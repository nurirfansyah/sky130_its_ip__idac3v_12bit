magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 6540 -3232 6550 -3219
rect 6474 -3274 6550 -3232
rect 6674 -3574 6774 -3450
rect 6674 -3628 6676 -3574
rect 6359 -4371 6503 -4324
rect 6540 -4371 6557 -4270
rect 6359 -4382 6475 -4371
rect 6445 -4407 6475 -4382
rect 6457 -4906 6475 -4407
rect 7639 -4848 7686 -4483
rect 7693 -4848 7740 -4537
rect 7608 -4943 7811 -4848
rect 7608 -5067 8313 -4943
rect 7608 -6152 8366 -5067
rect 7219 -6170 8366 -6152
rect 7657 -6181 8366 -6170
rect 7657 -6217 8331 -6181
rect 7840 -6235 8331 -6217
<< error_s >>
rect 3344 -2965 3460 -2899
rect 3460 -3219 3846 -3153
rect 3196 -3232 3206 -3219
rect 3130 -3274 3206 -3232
rect 3258 -3274 3846 -3219
rect 3130 -3277 3846 -3274
rect 3130 -3514 3274 -3277
rect 3460 -3299 3846 -3277
rect 3384 -3385 3846 -3299
rect 3388 -3393 3588 -3385
rect 3404 -3397 3572 -3393
rect 3130 -3600 3304 -3514
rect 3330 -3574 3430 -3450
rect 3330 -3628 3332 -3574
rect 3015 -4371 3159 -4324
rect 3196 -4371 3213 -4270
rect 3015 -4382 3787 -4371
rect 3101 -4407 3787 -4382
rect 3113 -4436 3787 -4407
rect 3113 -4848 3846 -4436
rect 4295 -4848 4342 -4483
rect 4349 -4848 4396 -4537
rect 3113 -4906 4467 -4848
rect 2540 -4943 4467 -4906
rect 2540 -5067 4969 -4943
rect 2540 -6022 5022 -5067
rect 5884 -6022 6348 -4906
rect 3131 -6087 5022 -6022
rect 3722 -6147 5022 -6087
rect 3751 -6152 5022 -6147
rect 3875 -6170 5022 -6152
rect 4313 -6181 5022 -6170
rect 4313 -6217 4987 -6181
rect 4496 -6235 4987 -6217
<< error_ps >>
rect 6474 -3514 6618 -3274
rect 6474 -3600 6648 -3514
rect 6475 -4436 7131 -4371
rect 6475 -4848 7190 -4436
rect 6475 -4906 7608 -4848
rect 6348 -6022 7608 -4906
rect 6475 -6087 7608 -6022
rect 7066 -6147 7608 -6087
rect 7095 -6152 7608 -6147
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use icell1scs  x1
timestamp 1717439242
transform 1 0 66 0 1 258
box -66 -6595 5022 200
use icell1scs  x2
timestamp 1717439242
transform 1 0 3410 0 1 258
box -66 -6595 5022 200
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
