magic
tech sky130A
magscale 1 2
timestamp 1717444414
<< nwell >>
rect 1168 -1780 1202 -1632
rect 2972 -1922 3030 -1866
rect 2366 -1992 2424 -1942
<< pwell >>
rect 1168 -2512 4842 -2182
<< locali >>
rect 2378 -2102 2412 -1982
rect 2984 -2104 3018 -1912
<< viali >>
rect 2984 -1912 3018 -1878
rect 2378 -1982 2412 -1948
rect 1288 -2144 1322 -2110
rect 2154 -2136 2188 -2102
rect 2258 -2136 2292 -2102
rect 2378 -2136 2412 -2102
rect 2496 -2136 2530 -2102
rect 2864 -2148 2898 -2114
rect 2984 -2138 3018 -2104
rect 3114 -2138 3148 -2104
rect 3288 -2136 3322 -2102
rect 3542 -2136 3576 -2102
rect 3900 -2146 3934 -2112
rect 4128 -2146 4162 -2112
rect 4328 -2164 4362 -2130
rect 3284 -2246 3318 -2212
rect 1480 -2300 1514 -2266
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 1212 -1632 4774 -1630
rect 1168 -1780 4774 -1632
rect 0 -2000 200 -1800
rect 2972 -1872 3030 -1866
rect 1283 -1878 3030 -1872
rect 1283 -1912 2984 -1878
rect 3018 -1880 3030 -1878
rect 3018 -1912 4366 -1880
rect 1283 -1914 4366 -1912
rect 1283 -2104 1325 -1914
rect 2972 -1922 4366 -1914
rect 2366 -1948 2424 -1942
rect 2366 -1982 2378 -1948
rect 2412 -1950 2424 -1948
rect 2412 -1982 4166 -1950
rect 2366 -1992 4166 -1982
rect 2150 -2062 3938 -2020
rect 2150 -2090 2192 -2062
rect 2142 -2102 2200 -2090
rect 1276 -2110 1334 -2104
rect 1276 -2144 1288 -2110
rect 1322 -2144 1334 -2110
rect 1276 -2156 1334 -2144
rect 2142 -2136 2154 -2102
rect 2188 -2136 2200 -2102
rect 2142 -2148 2200 -2136
rect 2246 -2098 2298 -2090
rect 2372 -2098 2418 -2096
rect 2490 -2098 2542 -2090
rect 2246 -2102 2542 -2098
rect 2246 -2136 2258 -2102
rect 2292 -2136 2378 -2102
rect 2412 -2136 2496 -2102
rect 2530 -2136 2542 -2102
rect 2246 -2140 2542 -2136
rect 2246 -2148 2298 -2140
rect 2372 -2142 2418 -2140
rect 2490 -2148 2542 -2140
rect 2854 -2114 2906 -2100
rect 2854 -2148 2864 -2114
rect 2898 -2148 2906 -2114
rect 0 -2400 200 -2200
rect 1472 -2266 1526 -2254
rect 1472 -2300 1480 -2266
rect 1514 -2274 1526 -2266
rect 2150 -2274 2192 -2148
rect 2854 -2158 2906 -2148
rect 2954 -2104 3170 -2090
rect 2954 -2138 2984 -2104
rect 3018 -2138 3114 -2104
rect 3148 -2138 3170 -2104
rect 2954 -2150 3170 -2138
rect 3278 -2098 3330 -2090
rect 3536 -2098 3588 -2090
rect 3278 -2102 3588 -2098
rect 3896 -2100 3938 -2062
rect 3278 -2136 3288 -2102
rect 3322 -2136 3542 -2102
rect 3576 -2136 3588 -2102
rect 3278 -2140 3588 -2136
rect 3278 -2148 3330 -2140
rect 3536 -2148 3588 -2140
rect 3890 -2112 3942 -2100
rect 4124 -2106 4166 -1992
rect 3890 -2146 3900 -2112
rect 3934 -2146 3942 -2112
rect 3890 -2158 3942 -2146
rect 4116 -2112 4174 -2106
rect 4116 -2146 4128 -2112
rect 4162 -2146 4174 -2112
rect 4324 -2124 4366 -1922
rect 4116 -2158 4174 -2146
rect 4316 -2130 4374 -2124
rect 2858 -2208 2900 -2158
rect 4316 -2164 4328 -2130
rect 4362 -2164 4374 -2130
rect 4316 -2176 4374 -2164
rect 3278 -2208 3330 -2200
rect 2858 -2212 3330 -2208
rect 2858 -2246 3284 -2212
rect 3318 -2246 3330 -2212
rect 2858 -2250 3330 -2246
rect 3278 -2258 3330 -2250
rect 1514 -2300 2192 -2274
rect 1472 -2316 2192 -2300
rect 1168 -2492 4774 -2344
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use pcell1scs  x1
timestamp 1717434410
transform -1 0 4548 0 -1 1272
box 710 -1488 3380 2844
use ncell1scs  x2
timestamp 1717414943
transform -1 0 3682 0 -1 -6068
box 149 -3548 2514 -422
use sky130_fd_sc_hvl__nand2_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 3490 0 1 -2469
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 3070 0 1 -2469
box -66 -43 354 897
use sky130_fd_sc_hvl__and2_1  x5 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 1234 0 1 -2469
box -66 -43 738 897
use sky130_fd_sc_hvl__inv_1  x6
timestamp 1710522493
transform 1 0 2038 0 1 -2469
box -66 -43 354 897
use sky130_fd_sc_hvl__nand2_1  x7
timestamp 1710522493
transform 1 0 2458 0 1 -2469
box -66 -43 546 897
use sky130_fd_sc_hvl__and2_1  x8
timestamp 1710522493
transform 1 0 4102 0 1 -2469
box -66 -43 738 897
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
