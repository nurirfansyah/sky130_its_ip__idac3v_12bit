magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 3344 -2965 3460 -2899
rect 6688 -2965 6804 -2899
rect 10032 -2965 10148 -2899
rect 13376 -2965 13492 -2899
rect 16720 -2965 16836 -2899
rect 20064 -2965 20180 -2899
rect 23408 -2965 23524 -2899
rect 26752 -2965 26868 -2899
rect 30096 -2965 30212 -2899
rect 33440 -2965 33556 -2899
rect 36784 -2965 36900 -2899
rect 40128 -2965 40244 -2899
rect 43472 -2965 43588 -2899
rect 46816 -2965 46932 -2899
rect 50160 -2965 50276 -2899
rect 53504 -2965 53620 -2899
rect 56848 -2965 56964 -2899
rect 60192 -2965 60308 -2899
rect 63536 -2965 63652 -2899
rect 66880 -2965 66996 -2899
rect 70224 -2965 70340 -2899
rect 73568 -2965 73684 -2899
rect 76912 -2965 77028 -2899
rect 80256 -2965 80372 -2899
rect 83600 -2965 83716 -2899
rect 86944 -2965 87060 -2899
rect 90288 -2965 90404 -2899
rect 93632 -2965 93748 -2899
rect 96976 -2965 97092 -2899
rect 100320 -2965 100436 -2899
rect 103664 -2965 103780 -2899
rect 110352 -2965 110468 -2899
rect 113696 -2965 113812 -2899
rect 117040 -2965 117156 -2899
rect 120384 -2965 120500 -2899
rect 123728 -2965 123844 -2899
rect 127072 -2965 127188 -2899
rect 130416 -2965 130532 -2899
rect 133760 -2965 133876 -2899
rect 137104 -2965 137220 -2899
rect 140448 -2965 140564 -2899
rect 143792 -2965 143908 -2899
rect 147136 -2965 147252 -2899
rect 150480 -2965 150596 -2899
rect 153824 -2965 153940 -2899
rect 157168 -2965 157284 -2899
rect 160512 -2965 160628 -2899
rect 163856 -2965 163972 -2899
rect 167200 -2965 167316 -2899
rect 170544 -2965 170660 -2899
rect 173888 -2965 174004 -2899
rect 177232 -2965 177348 -2899
rect 180576 -2965 180692 -2899
rect 183920 -2965 184036 -2899
rect 187264 -2965 187380 -2899
rect 190608 -2965 190724 -2899
rect 193952 -2965 194068 -2899
rect 197296 -2965 197412 -2899
rect 200640 -2965 200756 -2899
rect 203984 -2965 204100 -2899
rect 207328 -2965 207444 -2899
rect 210672 -2965 210788 -2899
rect 3460 -3219 3846 -3153
rect 6804 -3219 7190 -3153
rect 10148 -3219 10534 -3153
rect 13492 -3219 13878 -3153
rect 16836 -3219 17222 -3153
rect 20180 -3219 20566 -3153
rect 23524 -3219 23910 -3153
rect 26868 -3219 27254 -3153
rect 30212 -3219 30598 -3153
rect 33556 -3219 33942 -3153
rect 36900 -3219 37286 -3153
rect 40244 -3219 40630 -3153
rect 43588 -3219 43974 -3153
rect 46932 -3219 47318 -3153
rect 50276 -3219 50662 -3153
rect 53620 -3219 54006 -3153
rect 56964 -3219 57350 -3153
rect 60308 -3219 60694 -3153
rect 63652 -3219 64038 -3153
rect 66996 -3219 67382 -3153
rect 70340 -3219 70726 -3153
rect 73684 -3219 74070 -3153
rect 77028 -3219 77414 -3153
rect 80372 -3219 80758 -3153
rect 83716 -3219 84102 -3153
rect 87060 -3219 87446 -3153
rect 90404 -3219 90790 -3153
rect 93748 -3219 94134 -3153
rect 97092 -3219 97478 -3153
rect 100436 -3219 100822 -3153
rect 103780 -3219 104166 -3153
rect 3196 -3232 3206 -3219
rect 3130 -3274 3206 -3232
rect 3258 -3274 3846 -3219
rect 6540 -3232 6550 -3219
rect 3130 -3277 3846 -3274
rect 3130 -3514 3274 -3277
rect 3460 -3299 3846 -3277
rect 3384 -3385 3846 -3299
rect 6474 -3274 6550 -3232
rect 6602 -3274 7190 -3219
rect 9884 -3232 9894 -3219
rect 6474 -3277 7190 -3274
rect 3388 -3393 3588 -3385
rect 3404 -3397 3572 -3393
rect 3130 -3600 3304 -3514
rect 3330 -3574 3430 -3450
rect 6474 -3514 6618 -3277
rect 6804 -3299 7190 -3277
rect 6728 -3385 7190 -3299
rect 9818 -3274 9894 -3232
rect 9946 -3274 10534 -3219
rect 13228 -3232 13238 -3219
rect 9818 -3277 10534 -3274
rect 6732 -3393 6932 -3385
rect 6748 -3397 6916 -3393
rect 3330 -3628 3332 -3574
rect 6474 -3600 6648 -3514
rect 6674 -3574 6774 -3450
rect 9818 -3514 9962 -3277
rect 10148 -3299 10534 -3277
rect 10072 -3385 10534 -3299
rect 13162 -3274 13238 -3232
rect 13290 -3274 13878 -3219
rect 16572 -3232 16582 -3219
rect 13162 -3277 13878 -3274
rect 10076 -3393 10276 -3385
rect 10092 -3397 10260 -3393
rect 6674 -3628 6676 -3574
rect 9818 -3600 9992 -3514
rect 10018 -3574 10118 -3450
rect 13162 -3514 13306 -3277
rect 13492 -3299 13878 -3277
rect 13416 -3385 13878 -3299
rect 16506 -3274 16582 -3232
rect 16634 -3274 17222 -3219
rect 19916 -3232 19926 -3219
rect 16506 -3277 17222 -3274
rect 13420 -3393 13620 -3385
rect 13436 -3397 13604 -3393
rect 10018 -3628 10020 -3574
rect 13162 -3600 13336 -3514
rect 13362 -3574 13462 -3450
rect 16506 -3514 16650 -3277
rect 16836 -3299 17222 -3277
rect 16760 -3385 17222 -3299
rect 19850 -3274 19926 -3232
rect 19978 -3274 20566 -3219
rect 23260 -3232 23270 -3219
rect 19850 -3277 20566 -3274
rect 16764 -3393 16964 -3385
rect 16780 -3397 16948 -3393
rect 13362 -3628 13364 -3574
rect 16506 -3600 16680 -3514
rect 16706 -3574 16806 -3450
rect 19850 -3514 19994 -3277
rect 20180 -3299 20566 -3277
rect 20104 -3385 20566 -3299
rect 23194 -3274 23270 -3232
rect 23322 -3274 23910 -3219
rect 26604 -3232 26614 -3219
rect 23194 -3277 23910 -3274
rect 20108 -3393 20308 -3385
rect 20124 -3397 20292 -3393
rect 16706 -3628 16708 -3574
rect 19850 -3600 20024 -3514
rect 20050 -3574 20150 -3450
rect 23194 -3514 23338 -3277
rect 23524 -3299 23910 -3277
rect 23448 -3385 23910 -3299
rect 26538 -3274 26614 -3232
rect 26666 -3274 27254 -3219
rect 29948 -3232 29958 -3219
rect 26538 -3277 27254 -3274
rect 23452 -3393 23652 -3385
rect 23468 -3397 23636 -3393
rect 20050 -3628 20052 -3574
rect 23194 -3600 23368 -3514
rect 23394 -3574 23494 -3450
rect 26538 -3514 26682 -3277
rect 26868 -3299 27254 -3277
rect 26792 -3385 27254 -3299
rect 29882 -3274 29958 -3232
rect 30010 -3274 30598 -3219
rect 33292 -3232 33302 -3219
rect 29882 -3277 30598 -3274
rect 26796 -3393 26996 -3385
rect 26812 -3397 26980 -3393
rect 23394 -3628 23396 -3574
rect 26538 -3600 26712 -3514
rect 26738 -3574 26838 -3450
rect 29882 -3514 30026 -3277
rect 30212 -3299 30598 -3277
rect 30136 -3385 30598 -3299
rect 33226 -3274 33302 -3232
rect 33354 -3274 33942 -3219
rect 36636 -3232 36646 -3219
rect 33226 -3277 33942 -3274
rect 30140 -3393 30340 -3385
rect 30156 -3397 30324 -3393
rect 26738 -3628 26740 -3574
rect 29882 -3600 30056 -3514
rect 30082 -3574 30182 -3450
rect 33226 -3514 33370 -3277
rect 33556 -3299 33942 -3277
rect 33480 -3385 33942 -3299
rect 36570 -3274 36646 -3232
rect 36698 -3274 37286 -3219
rect 39980 -3232 39990 -3219
rect 36570 -3277 37286 -3274
rect 33484 -3393 33684 -3385
rect 33500 -3397 33668 -3393
rect 30082 -3628 30084 -3574
rect 33226 -3600 33400 -3514
rect 33426 -3574 33526 -3450
rect 36570 -3514 36714 -3277
rect 36900 -3299 37286 -3277
rect 36824 -3385 37286 -3299
rect 39914 -3274 39990 -3232
rect 40042 -3274 40630 -3219
rect 43324 -3232 43334 -3219
rect 39914 -3277 40630 -3274
rect 36828 -3393 37028 -3385
rect 36844 -3397 37012 -3393
rect 33426 -3628 33428 -3574
rect 36570 -3600 36744 -3514
rect 36770 -3574 36870 -3450
rect 39914 -3514 40058 -3277
rect 40244 -3299 40630 -3277
rect 40168 -3385 40630 -3299
rect 43258 -3274 43334 -3232
rect 43386 -3274 43974 -3219
rect 46668 -3232 46678 -3219
rect 43258 -3277 43974 -3274
rect 40172 -3393 40372 -3385
rect 40188 -3397 40356 -3393
rect 36770 -3628 36772 -3574
rect 39914 -3600 40088 -3514
rect 40114 -3574 40214 -3450
rect 43258 -3514 43402 -3277
rect 43588 -3299 43974 -3277
rect 43512 -3385 43974 -3299
rect 46602 -3274 46678 -3232
rect 46730 -3274 47318 -3219
rect 50012 -3232 50022 -3219
rect 46602 -3277 47318 -3274
rect 43516 -3393 43716 -3385
rect 43532 -3397 43700 -3393
rect 40114 -3628 40116 -3574
rect 43258 -3600 43432 -3514
rect 43458 -3574 43558 -3450
rect 46602 -3514 46746 -3277
rect 46932 -3299 47318 -3277
rect 46856 -3385 47318 -3299
rect 49946 -3274 50022 -3232
rect 50074 -3274 50662 -3219
rect 53356 -3232 53366 -3219
rect 49946 -3277 50662 -3274
rect 46860 -3393 47060 -3385
rect 46876 -3397 47044 -3393
rect 43458 -3628 43460 -3574
rect 46602 -3600 46776 -3514
rect 46802 -3574 46902 -3450
rect 49946 -3514 50090 -3277
rect 50276 -3299 50662 -3277
rect 50200 -3385 50662 -3299
rect 53290 -3274 53366 -3232
rect 53418 -3274 54006 -3219
rect 56700 -3232 56710 -3219
rect 53290 -3277 54006 -3274
rect 50204 -3393 50404 -3385
rect 50220 -3397 50388 -3393
rect 46802 -3628 46804 -3574
rect 49946 -3600 50120 -3514
rect 50146 -3574 50246 -3450
rect 53290 -3514 53434 -3277
rect 53620 -3299 54006 -3277
rect 53544 -3385 54006 -3299
rect 56634 -3274 56710 -3232
rect 56762 -3274 57350 -3219
rect 60044 -3232 60054 -3219
rect 56634 -3277 57350 -3274
rect 53548 -3393 53748 -3385
rect 53564 -3397 53732 -3393
rect 50146 -3628 50148 -3574
rect 53290 -3600 53464 -3514
rect 53490 -3574 53590 -3450
rect 56634 -3514 56778 -3277
rect 56964 -3299 57350 -3277
rect 56888 -3385 57350 -3299
rect 59978 -3274 60054 -3232
rect 60106 -3274 60694 -3219
rect 63388 -3232 63398 -3219
rect 59978 -3277 60694 -3274
rect 56892 -3393 57092 -3385
rect 56908 -3397 57076 -3393
rect 53490 -3628 53492 -3574
rect 56634 -3600 56808 -3514
rect 56834 -3574 56934 -3450
rect 59978 -3514 60122 -3277
rect 60308 -3299 60694 -3277
rect 60232 -3385 60694 -3299
rect 63322 -3274 63398 -3232
rect 63450 -3274 64038 -3219
rect 66732 -3232 66742 -3219
rect 63322 -3277 64038 -3274
rect 60236 -3393 60436 -3385
rect 60252 -3397 60420 -3393
rect 56834 -3628 56836 -3574
rect 59978 -3600 60152 -3514
rect 60178 -3574 60278 -3450
rect 63322 -3514 63466 -3277
rect 63652 -3299 64038 -3277
rect 63576 -3385 64038 -3299
rect 66666 -3274 66742 -3232
rect 66794 -3274 67382 -3219
rect 70076 -3232 70086 -3219
rect 66666 -3277 67382 -3274
rect 63580 -3393 63780 -3385
rect 63596 -3397 63764 -3393
rect 60178 -3628 60180 -3574
rect 63322 -3600 63496 -3514
rect 63522 -3574 63622 -3450
rect 66666 -3514 66810 -3277
rect 66996 -3299 67382 -3277
rect 66920 -3385 67382 -3299
rect 70010 -3274 70086 -3232
rect 70138 -3274 70726 -3219
rect 73420 -3232 73430 -3219
rect 70010 -3277 70726 -3274
rect 66924 -3393 67124 -3385
rect 66940 -3397 67108 -3393
rect 63522 -3628 63524 -3574
rect 66666 -3600 66840 -3514
rect 66866 -3574 66966 -3450
rect 70010 -3514 70154 -3277
rect 70340 -3299 70726 -3277
rect 70264 -3385 70726 -3299
rect 73354 -3274 73430 -3232
rect 73482 -3274 74070 -3219
rect 76764 -3232 76774 -3219
rect 73354 -3277 74070 -3274
rect 70268 -3393 70468 -3385
rect 70284 -3397 70452 -3393
rect 66866 -3628 66868 -3574
rect 70010 -3600 70184 -3514
rect 70210 -3574 70310 -3450
rect 73354 -3514 73498 -3277
rect 73684 -3299 74070 -3277
rect 73608 -3385 74070 -3299
rect 76698 -3274 76774 -3232
rect 76826 -3274 77414 -3219
rect 80108 -3232 80118 -3219
rect 76698 -3277 77414 -3274
rect 73612 -3393 73812 -3385
rect 73628 -3397 73796 -3393
rect 70210 -3628 70212 -3574
rect 73354 -3600 73528 -3514
rect 73554 -3574 73654 -3450
rect 76698 -3514 76842 -3277
rect 77028 -3299 77414 -3277
rect 76952 -3385 77414 -3299
rect 80042 -3274 80118 -3232
rect 80170 -3274 80758 -3219
rect 83452 -3232 83462 -3219
rect 80042 -3277 80758 -3274
rect 76956 -3393 77156 -3385
rect 76972 -3397 77140 -3393
rect 73554 -3628 73556 -3574
rect 76698 -3600 76872 -3514
rect 76898 -3574 76998 -3450
rect 80042 -3514 80186 -3277
rect 80372 -3299 80758 -3277
rect 80296 -3385 80758 -3299
rect 83386 -3274 83462 -3232
rect 83514 -3274 84102 -3219
rect 86796 -3232 86806 -3219
rect 83386 -3277 84102 -3274
rect 80300 -3393 80500 -3385
rect 80316 -3397 80484 -3393
rect 76898 -3628 76900 -3574
rect 80042 -3600 80216 -3514
rect 80242 -3574 80342 -3450
rect 83386 -3514 83530 -3277
rect 83716 -3299 84102 -3277
rect 83640 -3385 84102 -3299
rect 86730 -3274 86806 -3232
rect 86858 -3274 87446 -3219
rect 90140 -3232 90150 -3219
rect 86730 -3277 87446 -3274
rect 83644 -3393 83844 -3385
rect 83660 -3397 83828 -3393
rect 80242 -3628 80244 -3574
rect 83386 -3600 83560 -3514
rect 83586 -3574 83686 -3450
rect 86730 -3514 86874 -3277
rect 87060 -3299 87446 -3277
rect 86984 -3385 87446 -3299
rect 90074 -3274 90150 -3232
rect 90202 -3274 90790 -3219
rect 93484 -3232 93494 -3219
rect 90074 -3277 90790 -3274
rect 86988 -3393 87188 -3385
rect 87004 -3397 87172 -3393
rect 83586 -3628 83588 -3574
rect 86730 -3600 86904 -3514
rect 86930 -3574 87030 -3450
rect 90074 -3514 90218 -3277
rect 90404 -3299 90790 -3277
rect 90328 -3385 90790 -3299
rect 93418 -3274 93494 -3232
rect 93546 -3274 94134 -3219
rect 96828 -3232 96838 -3219
rect 93418 -3277 94134 -3274
rect 90332 -3393 90532 -3385
rect 90348 -3397 90516 -3393
rect 86930 -3628 86932 -3574
rect 90074 -3600 90248 -3514
rect 90274 -3574 90374 -3450
rect 93418 -3514 93562 -3277
rect 93748 -3299 94134 -3277
rect 93672 -3385 94134 -3299
rect 96762 -3274 96838 -3232
rect 96890 -3274 97478 -3219
rect 100172 -3232 100182 -3219
rect 96762 -3277 97478 -3274
rect 93676 -3393 93876 -3385
rect 93692 -3397 93860 -3393
rect 90274 -3628 90276 -3574
rect 93418 -3600 93592 -3514
rect 93618 -3574 93718 -3450
rect 96762 -3514 96906 -3277
rect 97092 -3299 97478 -3277
rect 97016 -3385 97478 -3299
rect 100106 -3274 100182 -3232
rect 100234 -3274 100822 -3219
rect 103516 -3232 103526 -3219
rect 100106 -3277 100822 -3274
rect 97020 -3393 97220 -3385
rect 97036 -3397 97204 -3393
rect 93618 -3628 93620 -3574
rect 96762 -3600 96936 -3514
rect 96962 -3574 97062 -3450
rect 100106 -3514 100250 -3277
rect 100436 -3299 100822 -3277
rect 100360 -3385 100822 -3299
rect 103450 -3274 103526 -3232
rect 103578 -3274 104166 -3219
rect 103450 -3277 104166 -3274
rect 100364 -3393 100564 -3385
rect 100380 -3397 100548 -3393
rect 96962 -3628 96964 -3574
rect 100106 -3600 100280 -3514
rect 100306 -3574 100406 -3450
rect 103450 -3514 103594 -3277
rect 103780 -3299 104166 -3277
rect 103704 -3385 104166 -3299
rect 110204 -3232 110214 -3219
rect 103708 -3393 103908 -3385
rect 103724 -3397 103892 -3393
rect 100306 -3628 100308 -3574
rect 103450 -3600 103624 -3514
rect 103650 -3574 103750 -3450
rect 110138 -3274 110214 -3232
rect 110266 -3274 110468 -3219
rect 103650 -3628 103652 -3574
rect 110282 -3277 110468 -3274
rect 113812 -3219 114198 -3153
rect 117156 -3219 117542 -3153
rect 120500 -3219 120886 -3153
rect 123844 -3219 124230 -3153
rect 127188 -3219 127574 -3153
rect 130532 -3219 130918 -3153
rect 133876 -3219 134262 -3153
rect 137220 -3219 137606 -3153
rect 140564 -3219 140950 -3153
rect 143908 -3219 144294 -3153
rect 147252 -3219 147638 -3153
rect 150596 -3219 150982 -3153
rect 153940 -3219 154326 -3153
rect 157284 -3219 157670 -3153
rect 160628 -3219 161014 -3153
rect 163972 -3219 164358 -3153
rect 167316 -3219 167702 -3153
rect 170660 -3219 171046 -3153
rect 174004 -3219 174390 -3153
rect 177348 -3219 177734 -3153
rect 180692 -3219 181078 -3153
rect 184036 -3219 184422 -3153
rect 187380 -3219 187766 -3153
rect 190724 -3219 191110 -3153
rect 194068 -3219 194454 -3153
rect 197412 -3219 197798 -3153
rect 200756 -3219 201142 -3153
rect 204100 -3219 204486 -3153
rect 207444 -3219 207830 -3153
rect 210788 -3219 211174 -3153
rect 113548 -3232 113558 -3219
rect 113482 -3274 113558 -3232
rect 113610 -3274 114198 -3219
rect 116892 -3232 116902 -3219
rect 113482 -3277 114198 -3274
rect 110396 -3393 110596 -3385
rect 110412 -3397 110580 -3393
rect 110338 -3574 110438 -3450
rect 113482 -3514 113626 -3277
rect 113812 -3299 114198 -3277
rect 113736 -3385 114198 -3299
rect 116826 -3274 116902 -3232
rect 116954 -3274 117542 -3219
rect 120236 -3232 120246 -3219
rect 116826 -3277 117542 -3274
rect 113740 -3393 113940 -3385
rect 113756 -3397 113924 -3393
rect 110338 -3628 110340 -3574
rect 113482 -3600 113656 -3514
rect 113682 -3574 113782 -3450
rect 116826 -3514 116970 -3277
rect 117156 -3299 117542 -3277
rect 117080 -3385 117542 -3299
rect 120170 -3274 120246 -3232
rect 120298 -3274 120886 -3219
rect 123580 -3232 123590 -3219
rect 120170 -3277 120886 -3274
rect 117084 -3393 117284 -3385
rect 117100 -3397 117268 -3393
rect 113682 -3628 113684 -3574
rect 116826 -3600 117000 -3514
rect 117026 -3574 117126 -3450
rect 120170 -3514 120314 -3277
rect 120500 -3299 120886 -3277
rect 120424 -3385 120886 -3299
rect 123514 -3274 123590 -3232
rect 123642 -3274 124230 -3219
rect 126924 -3232 126934 -3219
rect 123514 -3277 124230 -3274
rect 120428 -3393 120628 -3385
rect 120444 -3397 120612 -3393
rect 117026 -3628 117028 -3574
rect 120170 -3600 120344 -3514
rect 120370 -3574 120470 -3450
rect 123514 -3514 123658 -3277
rect 123844 -3299 124230 -3277
rect 123768 -3385 124230 -3299
rect 126858 -3274 126934 -3232
rect 126986 -3274 127574 -3219
rect 130268 -3232 130278 -3219
rect 126858 -3277 127574 -3274
rect 123772 -3393 123972 -3385
rect 123788 -3397 123956 -3393
rect 120370 -3628 120372 -3574
rect 123514 -3600 123688 -3514
rect 123714 -3574 123814 -3450
rect 126858 -3514 127002 -3277
rect 127188 -3299 127574 -3277
rect 127112 -3385 127574 -3299
rect 130202 -3274 130278 -3232
rect 130330 -3274 130918 -3219
rect 133612 -3232 133622 -3219
rect 130202 -3277 130918 -3274
rect 127116 -3393 127316 -3385
rect 127132 -3397 127300 -3393
rect 123714 -3628 123716 -3574
rect 126858 -3600 127032 -3514
rect 127058 -3574 127158 -3450
rect 130202 -3514 130346 -3277
rect 130532 -3299 130918 -3277
rect 130456 -3385 130918 -3299
rect 133546 -3274 133622 -3232
rect 133674 -3274 134262 -3219
rect 136956 -3232 136966 -3219
rect 133546 -3277 134262 -3274
rect 130460 -3393 130660 -3385
rect 130476 -3397 130644 -3393
rect 127058 -3628 127060 -3574
rect 130202 -3600 130376 -3514
rect 130402 -3574 130502 -3450
rect 133546 -3514 133690 -3277
rect 133876 -3299 134262 -3277
rect 133800 -3385 134262 -3299
rect 136890 -3274 136966 -3232
rect 137018 -3274 137606 -3219
rect 140300 -3232 140310 -3219
rect 136890 -3277 137606 -3274
rect 133804 -3393 134004 -3385
rect 133820 -3397 133988 -3393
rect 130402 -3628 130404 -3574
rect 133546 -3600 133720 -3514
rect 133746 -3574 133846 -3450
rect 136890 -3514 137034 -3277
rect 137220 -3299 137606 -3277
rect 137144 -3385 137606 -3299
rect 140234 -3274 140310 -3232
rect 140362 -3274 140950 -3219
rect 143644 -3232 143654 -3219
rect 140234 -3277 140950 -3274
rect 137148 -3393 137348 -3385
rect 137164 -3397 137332 -3393
rect 133746 -3628 133748 -3574
rect 136890 -3600 137064 -3514
rect 137090 -3574 137190 -3450
rect 140234 -3514 140378 -3277
rect 140564 -3299 140950 -3277
rect 140488 -3385 140950 -3299
rect 143578 -3274 143654 -3232
rect 143706 -3274 144294 -3219
rect 146988 -3232 146998 -3219
rect 143578 -3277 144294 -3274
rect 140492 -3393 140692 -3385
rect 140508 -3397 140676 -3393
rect 137090 -3628 137092 -3574
rect 140234 -3600 140408 -3514
rect 140434 -3574 140534 -3450
rect 143578 -3514 143722 -3277
rect 143908 -3299 144294 -3277
rect 143832 -3385 144294 -3299
rect 146922 -3274 146998 -3232
rect 147050 -3274 147638 -3219
rect 150332 -3232 150342 -3219
rect 146922 -3277 147638 -3274
rect 143836 -3393 144036 -3385
rect 143852 -3397 144020 -3393
rect 140434 -3628 140436 -3574
rect 143578 -3600 143752 -3514
rect 143778 -3574 143878 -3450
rect 146922 -3514 147066 -3277
rect 147252 -3299 147638 -3277
rect 147176 -3385 147638 -3299
rect 150266 -3274 150342 -3232
rect 150394 -3274 150982 -3219
rect 153676 -3232 153686 -3219
rect 150266 -3277 150982 -3274
rect 147180 -3393 147380 -3385
rect 147196 -3397 147364 -3393
rect 143778 -3628 143780 -3574
rect 146922 -3600 147096 -3514
rect 147122 -3574 147222 -3450
rect 150266 -3514 150410 -3277
rect 150596 -3299 150982 -3277
rect 150520 -3385 150982 -3299
rect 153610 -3274 153686 -3232
rect 153738 -3274 154326 -3219
rect 157020 -3232 157030 -3219
rect 153610 -3277 154326 -3274
rect 150524 -3393 150724 -3385
rect 150540 -3397 150708 -3393
rect 147122 -3628 147124 -3574
rect 150266 -3600 150440 -3514
rect 150466 -3574 150566 -3450
rect 153610 -3514 153754 -3277
rect 153940 -3299 154326 -3277
rect 153864 -3385 154326 -3299
rect 156954 -3274 157030 -3232
rect 157082 -3274 157670 -3219
rect 160364 -3232 160374 -3219
rect 156954 -3277 157670 -3274
rect 153868 -3393 154068 -3385
rect 153884 -3397 154052 -3393
rect 150466 -3628 150468 -3574
rect 153610 -3600 153784 -3514
rect 153810 -3574 153910 -3450
rect 156954 -3514 157098 -3277
rect 157284 -3299 157670 -3277
rect 157208 -3385 157670 -3299
rect 160298 -3274 160374 -3232
rect 160426 -3274 161014 -3219
rect 163708 -3232 163718 -3219
rect 160298 -3277 161014 -3274
rect 157212 -3393 157412 -3385
rect 157228 -3397 157396 -3393
rect 153810 -3628 153812 -3574
rect 156954 -3600 157128 -3514
rect 157154 -3574 157254 -3450
rect 160298 -3514 160442 -3277
rect 160628 -3299 161014 -3277
rect 160552 -3385 161014 -3299
rect 163642 -3274 163718 -3232
rect 163770 -3274 164358 -3219
rect 167052 -3232 167062 -3219
rect 163642 -3277 164358 -3274
rect 160556 -3393 160756 -3385
rect 160572 -3397 160740 -3393
rect 157154 -3628 157156 -3574
rect 160298 -3600 160472 -3514
rect 160498 -3574 160598 -3450
rect 163642 -3514 163786 -3277
rect 163972 -3299 164358 -3277
rect 163896 -3385 164358 -3299
rect 166986 -3274 167062 -3232
rect 167114 -3274 167702 -3219
rect 170396 -3232 170406 -3219
rect 166986 -3277 167702 -3274
rect 163900 -3393 164100 -3385
rect 163916 -3397 164084 -3393
rect 160498 -3628 160500 -3574
rect 163642 -3600 163816 -3514
rect 163842 -3574 163942 -3450
rect 166986 -3514 167130 -3277
rect 167316 -3299 167702 -3277
rect 167240 -3385 167702 -3299
rect 170330 -3274 170406 -3232
rect 170458 -3274 171046 -3219
rect 173740 -3232 173750 -3219
rect 170330 -3277 171046 -3274
rect 167244 -3393 167444 -3385
rect 167260 -3397 167428 -3393
rect 163842 -3628 163844 -3574
rect 166986 -3600 167160 -3514
rect 167186 -3574 167286 -3450
rect 170330 -3514 170474 -3277
rect 170660 -3299 171046 -3277
rect 170584 -3385 171046 -3299
rect 173674 -3274 173750 -3232
rect 173802 -3274 174390 -3219
rect 177084 -3232 177094 -3219
rect 173674 -3277 174390 -3274
rect 170588 -3393 170788 -3385
rect 170604 -3397 170772 -3393
rect 167186 -3628 167188 -3574
rect 170330 -3600 170504 -3514
rect 170530 -3574 170630 -3450
rect 173674 -3514 173818 -3277
rect 174004 -3299 174390 -3277
rect 173928 -3385 174390 -3299
rect 177018 -3274 177094 -3232
rect 177146 -3274 177734 -3219
rect 180428 -3232 180438 -3219
rect 177018 -3277 177734 -3274
rect 173932 -3393 174132 -3385
rect 173948 -3397 174116 -3393
rect 170530 -3628 170532 -3574
rect 173674 -3600 173848 -3514
rect 173874 -3574 173974 -3450
rect 177018 -3514 177162 -3277
rect 177348 -3299 177734 -3277
rect 177272 -3385 177734 -3299
rect 180362 -3274 180438 -3232
rect 180490 -3274 181078 -3219
rect 183772 -3232 183782 -3219
rect 180362 -3277 181078 -3274
rect 177276 -3393 177476 -3385
rect 177292 -3397 177460 -3393
rect 173874 -3628 173876 -3574
rect 177018 -3600 177192 -3514
rect 177218 -3574 177318 -3450
rect 180362 -3514 180506 -3277
rect 180692 -3299 181078 -3277
rect 180616 -3385 181078 -3299
rect 183706 -3274 183782 -3232
rect 183834 -3274 184422 -3219
rect 187116 -3232 187126 -3219
rect 183706 -3277 184422 -3274
rect 180620 -3393 180820 -3385
rect 180636 -3397 180804 -3393
rect 177218 -3628 177220 -3574
rect 180362 -3600 180536 -3514
rect 180562 -3574 180662 -3450
rect 183706 -3514 183850 -3277
rect 184036 -3299 184422 -3277
rect 183960 -3385 184422 -3299
rect 187050 -3274 187126 -3232
rect 187178 -3274 187766 -3219
rect 190460 -3232 190470 -3219
rect 187050 -3277 187766 -3274
rect 183964 -3393 184164 -3385
rect 183980 -3397 184148 -3393
rect 180562 -3628 180564 -3574
rect 183706 -3600 183880 -3514
rect 183906 -3574 184006 -3450
rect 187050 -3514 187194 -3277
rect 187380 -3299 187766 -3277
rect 187304 -3385 187766 -3299
rect 190394 -3274 190470 -3232
rect 190522 -3274 191110 -3219
rect 193804 -3232 193814 -3219
rect 190394 -3277 191110 -3274
rect 187308 -3393 187508 -3385
rect 187324 -3397 187492 -3393
rect 183906 -3628 183908 -3574
rect 187050 -3600 187224 -3514
rect 187250 -3574 187350 -3450
rect 190394 -3514 190538 -3277
rect 190724 -3299 191110 -3277
rect 190648 -3385 191110 -3299
rect 193738 -3274 193814 -3232
rect 193866 -3274 194454 -3219
rect 197148 -3232 197158 -3219
rect 193738 -3277 194454 -3274
rect 190652 -3393 190852 -3385
rect 190668 -3397 190836 -3393
rect 187250 -3628 187252 -3574
rect 190394 -3600 190568 -3514
rect 190594 -3574 190694 -3450
rect 193738 -3514 193882 -3277
rect 194068 -3299 194454 -3277
rect 193992 -3385 194454 -3299
rect 197082 -3274 197158 -3232
rect 197210 -3274 197798 -3219
rect 200492 -3232 200502 -3219
rect 197082 -3277 197798 -3274
rect 193996 -3393 194196 -3385
rect 194012 -3397 194180 -3393
rect 190594 -3628 190596 -3574
rect 193738 -3600 193912 -3514
rect 193938 -3574 194038 -3450
rect 197082 -3514 197226 -3277
rect 197412 -3299 197798 -3277
rect 197336 -3385 197798 -3299
rect 200426 -3274 200502 -3232
rect 200554 -3274 201142 -3219
rect 203836 -3232 203846 -3219
rect 200426 -3277 201142 -3274
rect 197340 -3393 197540 -3385
rect 197356 -3397 197524 -3393
rect 193938 -3628 193940 -3574
rect 197082 -3600 197256 -3514
rect 197282 -3574 197382 -3450
rect 200426 -3514 200570 -3277
rect 200756 -3299 201142 -3277
rect 200680 -3385 201142 -3299
rect 203770 -3274 203846 -3232
rect 203898 -3274 204486 -3219
rect 207180 -3232 207190 -3219
rect 203770 -3277 204486 -3274
rect 200684 -3393 200884 -3385
rect 200700 -3397 200868 -3393
rect 197282 -3628 197284 -3574
rect 200426 -3600 200600 -3514
rect 200626 -3574 200726 -3450
rect 203770 -3514 203914 -3277
rect 204100 -3299 204486 -3277
rect 204024 -3385 204486 -3299
rect 207114 -3274 207190 -3232
rect 207242 -3274 207830 -3219
rect 210524 -3232 210534 -3219
rect 207114 -3277 207830 -3274
rect 204028 -3393 204228 -3385
rect 204044 -3397 204212 -3393
rect 200626 -3628 200628 -3574
rect 203770 -3600 203944 -3514
rect 203970 -3574 204070 -3450
rect 207114 -3514 207258 -3277
rect 207444 -3299 207830 -3277
rect 207368 -3385 207830 -3299
rect 210458 -3274 210534 -3232
rect 210586 -3274 211174 -3219
rect 213868 -3232 213878 -3219
rect 210458 -3277 211174 -3274
rect 207372 -3393 207572 -3385
rect 207388 -3397 207556 -3393
rect 203970 -3628 203972 -3574
rect 207114 -3600 207288 -3514
rect 207314 -3574 207414 -3450
rect 210458 -3514 210602 -3277
rect 210788 -3299 211174 -3277
rect 210712 -3385 211174 -3299
rect 213802 -3274 213878 -3232
rect 210716 -3393 210916 -3385
rect 210732 -3397 210900 -3393
rect 207314 -3628 207316 -3574
rect 210458 -3600 210632 -3514
rect 210658 -3574 210758 -3450
rect 213802 -3514 213946 -3274
rect 210658 -3628 210660 -3574
rect 213802 -3600 213976 -3514
rect 214002 -3574 214102 -3450
rect 214002 -3628 214004 -3574
rect 3015 -4371 3159 -4324
rect 3196 -4371 3213 -4270
rect 6359 -4371 6503 -4324
rect 6540 -4371 6557 -4270
rect 9703 -4371 9847 -4324
rect 9884 -4371 9901 -4270
rect 13047 -4371 13191 -4324
rect 13228 -4371 13245 -4270
rect 16391 -4371 16535 -4324
rect 16572 -4371 16589 -4270
rect 19735 -4371 19879 -4324
rect 19916 -4371 19933 -4270
rect 23079 -4371 23223 -4324
rect 23260 -4371 23277 -4270
rect 26423 -4371 26567 -4324
rect 26604 -4371 26621 -4270
rect 29767 -4371 29911 -4324
rect 29948 -4371 29965 -4270
rect 33111 -4371 33255 -4324
rect 33292 -4371 33309 -4270
rect 36455 -4371 36599 -4324
rect 36636 -4371 36653 -4270
rect 39799 -4371 39943 -4324
rect 39980 -4371 39997 -4270
rect 43143 -4371 43287 -4324
rect 43324 -4371 43341 -4270
rect 46487 -4371 46631 -4324
rect 46668 -4371 46685 -4270
rect 49831 -4371 49975 -4324
rect 50012 -4371 50029 -4270
rect 53175 -4371 53319 -4324
rect 53356 -4371 53373 -4270
rect 56519 -4371 56663 -4324
rect 56700 -4371 56717 -4270
rect 59863 -4371 60007 -4324
rect 60044 -4371 60061 -4270
rect 63207 -4371 63351 -4324
rect 63388 -4371 63405 -4270
rect 66551 -4371 66695 -4324
rect 66732 -4371 66749 -4270
rect 69895 -4371 70039 -4324
rect 70076 -4371 70093 -4270
rect 73239 -4371 73383 -4324
rect 73420 -4371 73437 -4270
rect 76583 -4371 76727 -4324
rect 76764 -4371 76781 -4270
rect 79927 -4371 80071 -4324
rect 80108 -4371 80125 -4270
rect 83271 -4371 83415 -4324
rect 83452 -4371 83469 -4270
rect 86615 -4371 86759 -4324
rect 86796 -4371 86813 -4270
rect 89959 -4371 90103 -4324
rect 90140 -4371 90157 -4270
rect 93303 -4371 93447 -4324
rect 93484 -4371 93501 -4270
rect 96647 -4371 96791 -4324
rect 96828 -4371 96845 -4270
rect 99991 -4371 100135 -4324
rect 100172 -4371 100189 -4270
rect 103335 -4371 103479 -4324
rect 103516 -4371 103533 -4270
rect 110023 -4371 110167 -4324
rect 110204 -4371 110221 -4270
rect 113367 -4371 113511 -4324
rect 113548 -4371 113565 -4270
rect 116711 -4371 116855 -4324
rect 116892 -4371 116909 -4270
rect 120055 -4371 120199 -4324
rect 120236 -4371 120253 -4270
rect 123399 -4371 123543 -4324
rect 123580 -4371 123597 -4270
rect 126743 -4371 126887 -4324
rect 126924 -4371 126941 -4270
rect 130087 -4371 130231 -4324
rect 130268 -4371 130285 -4270
rect 133431 -4371 133575 -4324
rect 133612 -4371 133629 -4270
rect 136775 -4371 136919 -4324
rect 136956 -4371 136973 -4270
rect 140119 -4371 140263 -4324
rect 140300 -4371 140317 -4270
rect 143463 -4371 143607 -4324
rect 143644 -4371 143661 -4270
rect 146807 -4371 146951 -4324
rect 146988 -4371 147005 -4270
rect 150151 -4371 150295 -4324
rect 150332 -4371 150349 -4270
rect 153495 -4371 153639 -4324
rect 153676 -4371 153693 -4270
rect 156839 -4371 156983 -4324
rect 157020 -4371 157037 -4270
rect 160183 -4371 160327 -4324
rect 160364 -4371 160381 -4270
rect 163527 -4371 163671 -4324
rect 163708 -4371 163725 -4270
rect 166871 -4371 167015 -4324
rect 167052 -4371 167069 -4270
rect 170215 -4371 170359 -4324
rect 170396 -4371 170413 -4270
rect 173559 -4371 173703 -4324
rect 173740 -4371 173757 -4270
rect 176903 -4371 177047 -4324
rect 177084 -4371 177101 -4270
rect 180247 -4371 180391 -4324
rect 180428 -4371 180445 -4270
rect 183591 -4371 183735 -4324
rect 183772 -4371 183789 -4270
rect 186935 -4371 187079 -4324
rect 187116 -4371 187133 -4270
rect 190279 -4371 190423 -4324
rect 190460 -4371 190477 -4270
rect 193623 -4371 193767 -4324
rect 193804 -4371 193821 -4270
rect 196967 -4371 197111 -4324
rect 197148 -4371 197165 -4270
rect 200311 -4371 200455 -4324
rect 200492 -4371 200509 -4270
rect 203655 -4371 203799 -4324
rect 203836 -4371 203853 -4270
rect 206999 -4371 207143 -4324
rect 207180 -4371 207197 -4270
rect 210343 -4371 210487 -4324
rect 210524 -4371 210541 -4270
rect 213687 -4371 213831 -4324
rect 213868 -4371 213885 -4270
rect 3015 -4382 3787 -4371
rect 6359 -4382 7131 -4371
rect 9703 -4382 10475 -4371
rect 13047 -4382 13819 -4371
rect 16391 -4382 17163 -4371
rect 19735 -4382 20507 -4371
rect 23079 -4382 23851 -4371
rect 26423 -4382 27195 -4371
rect 29767 -4382 30539 -4371
rect 33111 -4382 33883 -4371
rect 36455 -4382 37227 -4371
rect 39799 -4382 40571 -4371
rect 43143 -4382 43915 -4371
rect 46487 -4382 47259 -4371
rect 49831 -4382 50603 -4371
rect 53175 -4382 53947 -4371
rect 56519 -4382 57291 -4371
rect 59863 -4382 60635 -4371
rect 63207 -4382 63979 -4371
rect 66551 -4382 67323 -4371
rect 69895 -4382 70667 -4371
rect 73239 -4382 74011 -4371
rect 76583 -4382 77355 -4371
rect 79927 -4382 80699 -4371
rect 83271 -4382 84043 -4371
rect 86615 -4382 87387 -4371
rect 89959 -4382 90731 -4371
rect 93303 -4382 94075 -4371
rect 96647 -4382 97419 -4371
rect 99991 -4382 100763 -4371
rect 103335 -4382 104107 -4371
rect 110023 -4382 110139 -4371
rect 3101 -4407 3787 -4382
rect 6445 -4407 7131 -4382
rect 9789 -4407 10475 -4382
rect 13133 -4407 13819 -4382
rect 16477 -4407 17163 -4382
rect 19821 -4407 20507 -4382
rect 23165 -4407 23851 -4382
rect 26509 -4407 27195 -4382
rect 29853 -4407 30539 -4382
rect 33197 -4407 33883 -4382
rect 36541 -4407 37227 -4382
rect 39885 -4407 40571 -4382
rect 43229 -4407 43915 -4382
rect 46573 -4407 47259 -4382
rect 49917 -4407 50603 -4382
rect 53261 -4407 53947 -4382
rect 56605 -4407 57291 -4382
rect 59949 -4407 60635 -4382
rect 63293 -4407 63979 -4382
rect 66637 -4407 67323 -4382
rect 69981 -4407 70667 -4382
rect 73325 -4407 74011 -4382
rect 76669 -4407 77355 -4382
rect 80013 -4407 80699 -4382
rect 83357 -4407 84043 -4382
rect 86701 -4407 87387 -4382
rect 90045 -4407 90731 -4382
rect 93389 -4407 94075 -4382
rect 96733 -4407 97419 -4382
rect 100077 -4407 100763 -4382
rect 103421 -4407 104107 -4382
rect 110109 -4407 110139 -4382
rect 3113 -4436 3787 -4407
rect 6457 -4436 7131 -4407
rect 9801 -4436 10475 -4407
rect 13145 -4436 13819 -4407
rect 16489 -4436 17163 -4407
rect 19833 -4436 20507 -4407
rect 23177 -4436 23851 -4407
rect 26521 -4436 27195 -4407
rect 29865 -4436 30539 -4407
rect 33209 -4436 33883 -4407
rect 36553 -4436 37227 -4407
rect 39897 -4436 40571 -4407
rect 43241 -4436 43915 -4407
rect 46585 -4436 47259 -4407
rect 49929 -4436 50603 -4407
rect 53273 -4436 53947 -4407
rect 56617 -4436 57291 -4407
rect 59961 -4436 60635 -4407
rect 63305 -4436 63979 -4407
rect 66649 -4436 67323 -4407
rect 69993 -4436 70667 -4407
rect 73337 -4436 74011 -4407
rect 76681 -4436 77355 -4407
rect 80025 -4436 80699 -4407
rect 83369 -4436 84043 -4407
rect 86713 -4436 87387 -4407
rect 90057 -4436 90731 -4407
rect 93401 -4436 94075 -4407
rect 96745 -4436 97419 -4407
rect 100089 -4436 100763 -4407
rect 103433 -4436 104107 -4407
rect 3113 -4848 3846 -4436
rect 4295 -4848 4342 -4483
rect 4349 -4848 4396 -4537
rect 6457 -4848 7190 -4436
rect 7639 -4848 7686 -4483
rect 7693 -4848 7740 -4537
rect 9801 -4848 10534 -4436
rect 10983 -4848 11030 -4483
rect 11037 -4848 11084 -4537
rect 13145 -4848 13878 -4436
rect 14327 -4848 14374 -4483
rect 14381 -4848 14428 -4537
rect 16489 -4848 17222 -4436
rect 17671 -4848 17718 -4483
rect 17725 -4848 17772 -4537
rect 19833 -4848 20566 -4436
rect 21015 -4848 21062 -4483
rect 21069 -4848 21116 -4537
rect 23177 -4848 23910 -4436
rect 24359 -4848 24406 -4483
rect 24413 -4848 24460 -4537
rect 26521 -4848 27254 -4436
rect 27703 -4848 27750 -4483
rect 27757 -4848 27804 -4537
rect 29865 -4848 30598 -4436
rect 31047 -4848 31094 -4483
rect 31101 -4848 31148 -4537
rect 33209 -4848 33942 -4436
rect 34391 -4848 34438 -4483
rect 34445 -4848 34492 -4537
rect 36553 -4848 37286 -4436
rect 37735 -4848 37782 -4483
rect 37789 -4848 37836 -4537
rect 39897 -4848 40630 -4436
rect 41079 -4848 41126 -4483
rect 41133 -4848 41180 -4537
rect 43241 -4848 43974 -4436
rect 44423 -4848 44470 -4483
rect 44477 -4848 44524 -4537
rect 46585 -4848 47318 -4436
rect 47767 -4848 47814 -4483
rect 47821 -4848 47868 -4537
rect 49929 -4848 50662 -4436
rect 51111 -4848 51158 -4483
rect 51165 -4848 51212 -4537
rect 53273 -4848 54006 -4436
rect 54455 -4848 54502 -4483
rect 54509 -4848 54556 -4537
rect 56617 -4848 57350 -4436
rect 57799 -4848 57846 -4483
rect 57853 -4848 57900 -4537
rect 59961 -4848 60694 -4436
rect 61143 -4848 61190 -4483
rect 61197 -4848 61244 -4537
rect 63305 -4848 64038 -4436
rect 64487 -4848 64534 -4483
rect 64541 -4848 64588 -4537
rect 66649 -4848 67382 -4436
rect 67831 -4848 67878 -4483
rect 67885 -4848 67932 -4537
rect 69993 -4848 70726 -4436
rect 71175 -4848 71222 -4483
rect 71229 -4848 71276 -4537
rect 73337 -4848 74070 -4436
rect 74519 -4848 74566 -4483
rect 74573 -4848 74620 -4537
rect 76681 -4848 77414 -4436
rect 77863 -4848 77910 -4483
rect 77917 -4848 77964 -4537
rect 80025 -4848 80758 -4436
rect 81207 -4848 81254 -4483
rect 81261 -4848 81308 -4537
rect 83369 -4848 84102 -4436
rect 84551 -4848 84598 -4483
rect 84605 -4848 84652 -4537
rect 86713 -4848 87446 -4436
rect 87895 -4848 87942 -4483
rect 87949 -4848 87996 -4537
rect 90057 -4848 90790 -4436
rect 91239 -4848 91286 -4483
rect 91293 -4848 91340 -4537
rect 93401 -4848 94134 -4436
rect 94583 -4848 94630 -4483
rect 94637 -4848 94684 -4537
rect 96745 -4848 97478 -4436
rect 97927 -4848 97974 -4483
rect 97981 -4848 98028 -4537
rect 100089 -4848 100822 -4436
rect 101271 -4848 101318 -4483
rect 101325 -4848 101372 -4537
rect 103433 -4848 104166 -4436
rect 104615 -4848 104662 -4483
rect 104669 -4848 104716 -4537
rect 3113 -4906 4467 -4848
rect 6457 -4906 7811 -4848
rect 9801 -4906 11155 -4848
rect 13145 -4906 14499 -4848
rect 16489 -4906 17843 -4848
rect 19833 -4906 21187 -4848
rect 23177 -4906 24531 -4848
rect 26521 -4906 27875 -4848
rect 29865 -4906 31219 -4848
rect 33209 -4906 34563 -4848
rect 36553 -4906 37907 -4848
rect 39897 -4906 41251 -4848
rect 43241 -4906 44595 -4848
rect 46585 -4906 47939 -4848
rect 49929 -4906 51283 -4848
rect 53273 -4906 54627 -4848
rect 56617 -4906 57971 -4848
rect 59961 -4906 61315 -4848
rect 63305 -4906 64659 -4848
rect 66649 -4906 68003 -4848
rect 69993 -4906 71347 -4848
rect 73337 -4906 74691 -4848
rect 76681 -4906 78035 -4848
rect 80025 -4906 81379 -4848
rect 83369 -4906 84723 -4848
rect 86713 -4906 88067 -4848
rect 90057 -4906 91411 -4848
rect 93401 -4906 94755 -4848
rect 96745 -4906 98099 -4848
rect 100089 -4906 101443 -4848
rect 103433 -4906 104488 -4848
rect 2720 -4943 4467 -4906
rect 5884 -4943 7811 -4906
rect 9228 -4943 11155 -4906
rect 12572 -4943 14499 -4906
rect 15916 -4943 17843 -4906
rect 19260 -4943 21187 -4906
rect 22604 -4943 24531 -4906
rect 25948 -4943 27875 -4906
rect 29292 -4943 31219 -4906
rect 32636 -4943 34563 -4906
rect 35980 -4943 37907 -4906
rect 39324 -4943 41251 -4906
rect 42668 -4943 44595 -4906
rect 46012 -4943 47939 -4906
rect 49356 -4943 51283 -4906
rect 52700 -4943 54627 -4906
rect 56044 -4943 57971 -4906
rect 59388 -4943 61315 -4906
rect 62732 -4943 64659 -4906
rect 66076 -4943 68003 -4906
rect 69420 -4943 71347 -4906
rect 72764 -4943 74691 -4906
rect 76108 -4943 78035 -4906
rect 79452 -4943 81379 -4906
rect 82796 -4943 84723 -4906
rect 86140 -4943 88067 -4906
rect 89484 -4943 91411 -4906
rect 92828 -4943 94755 -4906
rect 96172 -4943 98099 -4906
rect 99516 -4943 101443 -4906
rect 2720 -5067 4969 -4943
rect 5884 -5067 8313 -4943
rect 9228 -5067 11657 -4943
rect 12572 -5067 15001 -4943
rect 15916 -5067 18345 -4943
rect 19260 -5067 21689 -4943
rect 22604 -5067 25033 -4943
rect 25948 -5067 28377 -4943
rect 29292 -5067 31721 -4943
rect 32636 -5067 35065 -4943
rect 35980 -5067 38409 -4943
rect 39324 -5067 41753 -4943
rect 42668 -5067 45097 -4943
rect 46012 -5067 48441 -4943
rect 49356 -5067 51785 -4943
rect 52700 -5067 55129 -4943
rect 56044 -5067 58473 -4943
rect 59388 -5067 61817 -4943
rect 62732 -5067 65161 -4943
rect 66076 -5067 68505 -4943
rect 69420 -5067 71849 -4943
rect 72764 -5067 75193 -4943
rect 76108 -5067 78537 -4943
rect 79452 -5067 81881 -4943
rect 82796 -5067 85225 -4943
rect 86140 -5067 88569 -4943
rect 89484 -5067 91913 -4943
rect 92828 -5067 95257 -4943
rect 96172 -5067 98601 -4943
rect 99516 -5067 101945 -4943
rect 2720 -6022 5022 -5067
rect 5884 -6022 8366 -5067
rect 9228 -6022 11710 -5067
rect 12572 -6022 15054 -5067
rect 15916 -6022 18398 -5067
rect 19260 -6022 21742 -5067
rect 22604 -6022 25086 -5067
rect 25948 -6022 28430 -5067
rect 29292 -6022 31774 -5067
rect 32636 -6022 35118 -5067
rect 35980 -6022 38462 -5067
rect 39324 -6022 41806 -5067
rect 42668 -6022 45150 -5067
rect 46012 -6022 48494 -5067
rect 49356 -6022 51838 -5067
rect 52700 -6022 55182 -5067
rect 56044 -6022 58526 -5067
rect 59388 -6022 61870 -5067
rect 62732 -6022 65214 -5067
rect 66076 -6022 68558 -5067
rect 69420 -6022 71902 -5067
rect 72764 -6022 75246 -5067
rect 76108 -6022 78590 -5067
rect 79452 -6022 81934 -5067
rect 82796 -6022 85278 -5067
rect 86140 -6022 88622 -5067
rect 89484 -6022 91966 -5067
rect 92828 -6022 95310 -5067
rect 96172 -6022 98654 -5067
rect 99516 -6022 101998 -5067
rect 102860 -6022 104488 -4906
rect 110121 -4906 110139 -4407
rect 113367 -4382 114139 -4371
rect 116711 -4382 117483 -4371
rect 120055 -4382 120827 -4371
rect 123399 -4382 124171 -4371
rect 126743 -4382 127515 -4371
rect 130087 -4382 130859 -4371
rect 133431 -4382 134203 -4371
rect 136775 -4382 137547 -4371
rect 140119 -4382 140891 -4371
rect 143463 -4382 144235 -4371
rect 146807 -4382 147579 -4371
rect 150151 -4382 150923 -4371
rect 153495 -4382 154267 -4371
rect 156839 -4382 157611 -4371
rect 160183 -4382 160955 -4371
rect 163527 -4382 164299 -4371
rect 166871 -4382 167643 -4371
rect 170215 -4382 170987 -4371
rect 173559 -4382 174331 -4371
rect 176903 -4382 177675 -4371
rect 180247 -4382 181019 -4371
rect 183591 -4382 184363 -4371
rect 186935 -4382 187707 -4371
rect 190279 -4382 191051 -4371
rect 193623 -4382 194395 -4371
rect 196967 -4382 197739 -4371
rect 200311 -4382 201083 -4371
rect 203655 -4382 204427 -4371
rect 206999 -4382 207771 -4371
rect 210343 -4382 211115 -4371
rect 213687 -4382 214459 -4371
rect 113453 -4407 114139 -4382
rect 116797 -4407 117483 -4382
rect 120141 -4407 120827 -4382
rect 123485 -4407 124171 -4382
rect 126829 -4407 127515 -4382
rect 130173 -4407 130859 -4382
rect 133517 -4407 134203 -4382
rect 136861 -4407 137547 -4382
rect 140205 -4407 140891 -4382
rect 143549 -4407 144235 -4382
rect 146893 -4407 147579 -4382
rect 150237 -4407 150923 -4382
rect 153581 -4407 154267 -4382
rect 156925 -4407 157611 -4382
rect 160269 -4407 160955 -4382
rect 163613 -4407 164299 -4382
rect 166957 -4407 167643 -4382
rect 170301 -4407 170987 -4382
rect 173645 -4407 174331 -4382
rect 176989 -4407 177675 -4382
rect 180333 -4407 181019 -4382
rect 183677 -4407 184363 -4382
rect 187021 -4407 187707 -4382
rect 190365 -4407 191051 -4382
rect 193709 -4407 194395 -4382
rect 197053 -4407 197739 -4382
rect 200397 -4407 201083 -4382
rect 203741 -4407 204427 -4382
rect 207085 -4407 207771 -4382
rect 210429 -4407 211115 -4382
rect 213773 -4407 214459 -4382
rect 113465 -4436 114139 -4407
rect 116809 -4436 117483 -4407
rect 120153 -4436 120827 -4407
rect 123497 -4436 124171 -4407
rect 126841 -4436 127515 -4407
rect 130185 -4436 130859 -4407
rect 133529 -4436 134203 -4407
rect 136873 -4436 137547 -4407
rect 140217 -4436 140891 -4407
rect 143561 -4436 144235 -4407
rect 146905 -4436 147579 -4407
rect 150249 -4436 150923 -4407
rect 153593 -4436 154267 -4407
rect 156937 -4436 157611 -4407
rect 160281 -4436 160955 -4407
rect 163625 -4436 164299 -4407
rect 166969 -4436 167643 -4407
rect 170313 -4436 170987 -4407
rect 173657 -4436 174331 -4407
rect 177001 -4436 177675 -4407
rect 180345 -4436 181019 -4407
rect 183689 -4436 184363 -4407
rect 187033 -4436 187707 -4407
rect 190377 -4436 191051 -4407
rect 193721 -4436 194395 -4407
rect 197065 -4436 197739 -4407
rect 200409 -4436 201083 -4407
rect 203753 -4436 204427 -4407
rect 207097 -4436 207771 -4407
rect 210441 -4436 211115 -4407
rect 213785 -4436 214459 -4407
rect 111303 -4848 111350 -4483
rect 111357 -4848 111404 -4537
rect 113465 -4848 114198 -4436
rect 114647 -4848 114694 -4483
rect 114701 -4848 114748 -4537
rect 116809 -4848 117542 -4436
rect 117991 -4848 118038 -4483
rect 118045 -4848 118092 -4537
rect 120153 -4848 120886 -4436
rect 121335 -4848 121382 -4483
rect 121389 -4848 121436 -4537
rect 123497 -4848 124230 -4436
rect 124679 -4848 124726 -4483
rect 124733 -4848 124780 -4537
rect 126841 -4848 127574 -4436
rect 128023 -4848 128070 -4483
rect 128077 -4848 128124 -4537
rect 130185 -4848 130918 -4436
rect 131367 -4848 131414 -4483
rect 131421 -4848 131468 -4537
rect 133529 -4848 134262 -4436
rect 134711 -4848 134758 -4483
rect 134765 -4848 134812 -4537
rect 136873 -4848 137606 -4436
rect 138055 -4848 138102 -4483
rect 138109 -4848 138156 -4537
rect 140217 -4848 140950 -4436
rect 141399 -4848 141446 -4483
rect 141453 -4848 141500 -4537
rect 143561 -4848 144294 -4436
rect 144743 -4848 144790 -4483
rect 144797 -4848 144844 -4537
rect 146905 -4848 147638 -4436
rect 148087 -4848 148134 -4483
rect 148141 -4848 148188 -4537
rect 150249 -4848 150982 -4436
rect 151431 -4848 151478 -4483
rect 151485 -4848 151532 -4537
rect 153593 -4848 154326 -4436
rect 154775 -4848 154822 -4483
rect 154829 -4848 154876 -4537
rect 156937 -4848 157670 -4436
rect 158119 -4848 158166 -4483
rect 158173 -4848 158220 -4537
rect 160281 -4848 161014 -4436
rect 161463 -4848 161510 -4483
rect 161517 -4848 161564 -4537
rect 163625 -4848 164358 -4436
rect 164807 -4848 164854 -4483
rect 164861 -4848 164908 -4537
rect 166969 -4848 167702 -4436
rect 168151 -4848 168198 -4483
rect 168205 -4848 168252 -4537
rect 170313 -4848 171046 -4436
rect 171495 -4848 171542 -4483
rect 171549 -4848 171596 -4537
rect 173657 -4848 174390 -4436
rect 174839 -4848 174886 -4483
rect 174893 -4848 174940 -4537
rect 177001 -4848 177734 -4436
rect 178183 -4848 178230 -4483
rect 178237 -4848 178284 -4537
rect 180345 -4848 181078 -4436
rect 181527 -4848 181574 -4483
rect 181581 -4848 181628 -4537
rect 183689 -4848 184422 -4436
rect 184871 -4848 184918 -4483
rect 184925 -4848 184972 -4537
rect 187033 -4848 187766 -4436
rect 188215 -4848 188262 -4483
rect 188269 -4848 188316 -4537
rect 190377 -4848 191110 -4436
rect 191559 -4848 191606 -4483
rect 191613 -4848 191660 -4537
rect 193721 -4848 194454 -4436
rect 194903 -4848 194950 -4483
rect 194957 -4848 195004 -4537
rect 197065 -4848 197798 -4436
rect 198247 -4848 198294 -4483
rect 198301 -4848 198348 -4537
rect 200409 -4848 201142 -4436
rect 201591 -4848 201638 -4483
rect 201645 -4848 201692 -4537
rect 203753 -4848 204486 -4436
rect 204935 -4848 204982 -4483
rect 204989 -4848 205036 -4537
rect 207097 -4848 207830 -4436
rect 208279 -4848 208326 -4483
rect 208333 -4848 208380 -4537
rect 210441 -4848 211174 -4436
rect 211623 -4848 211670 -4483
rect 211677 -4848 211724 -4537
rect 213785 -4848 214518 -4436
rect 214967 -4848 215014 -4483
rect 215021 -4848 215068 -4537
rect 3131 -6087 5022 -6022
rect 6475 -6087 8366 -6022
rect 9819 -6087 11710 -6022
rect 13163 -6087 15054 -6022
rect 16507 -6087 18398 -6022
rect 19851 -6087 21742 -6022
rect 23195 -6087 25086 -6022
rect 26539 -6087 28430 -6022
rect 29883 -6087 31774 -6022
rect 33227 -6087 35118 -6022
rect 36571 -6087 38462 -6022
rect 39915 -6087 41806 -6022
rect 43259 -6087 45150 -6022
rect 46603 -6087 48494 -6022
rect 49947 -6087 51838 -6022
rect 53291 -6087 55182 -6022
rect 56635 -6087 58526 -6022
rect 59979 -6087 61870 -6022
rect 63323 -6087 65214 -6022
rect 66667 -6087 68558 -6022
rect 70011 -6087 71902 -6022
rect 73355 -6087 75246 -6022
rect 76699 -6087 78590 -6022
rect 80043 -6087 81934 -6022
rect 83387 -6087 85278 -6022
rect 86731 -6087 88622 -6022
rect 90075 -6087 91966 -6022
rect 93419 -6087 95310 -6022
rect 96763 -6087 98654 -6022
rect 100107 -6087 101998 -6022
rect 103451 -6087 104488 -6022
rect 3722 -6147 5022 -6087
rect 7066 -6147 8366 -6087
rect 10410 -6147 11710 -6087
rect 13754 -6147 15054 -6087
rect 17098 -6147 18398 -6087
rect 20442 -6147 21742 -6087
rect 23786 -6147 25086 -6087
rect 27130 -6147 28430 -6087
rect 30474 -6147 31774 -6087
rect 33818 -6147 35118 -6087
rect 37162 -6147 38462 -6087
rect 40506 -6147 41806 -6087
rect 43850 -6147 45150 -6087
rect 47194 -6147 48494 -6087
rect 50538 -6147 51838 -6087
rect 53882 -6147 55182 -6087
rect 57226 -6147 58526 -6087
rect 60570 -6147 61870 -6087
rect 63914 -6147 65214 -6087
rect 67258 -6147 68558 -6087
rect 70602 -6147 71902 -6087
rect 73946 -6147 75246 -6087
rect 77290 -6147 78590 -6087
rect 80634 -6147 81934 -6087
rect 83978 -6147 85278 -6087
rect 87322 -6147 88622 -6087
rect 90666 -6147 91966 -6087
rect 94010 -6147 95310 -6087
rect 97354 -6147 98654 -6087
rect 100698 -6147 101998 -6087
rect 104042 -6147 104488 -6087
rect 3751 -6152 5022 -6147
rect 7095 -6152 8366 -6147
rect 10439 -6152 11710 -6147
rect 13783 -6152 15054 -6147
rect 17127 -6152 18398 -6147
rect 20471 -6152 21742 -6147
rect 23815 -6152 25086 -6147
rect 27159 -6152 28430 -6147
rect 30503 -6152 31774 -6147
rect 33847 -6152 35118 -6147
rect 37191 -6152 38462 -6147
rect 40535 -6152 41806 -6147
rect 43879 -6152 45150 -6147
rect 47223 -6152 48494 -6147
rect 50567 -6152 51838 -6147
rect 53911 -6152 55182 -6147
rect 57255 -6152 58526 -6147
rect 60599 -6152 61870 -6147
rect 63943 -6152 65214 -6147
rect 67287 -6152 68558 -6147
rect 70631 -6152 71902 -6147
rect 73975 -6152 75246 -6147
rect 77319 -6152 78590 -6147
rect 80663 -6152 81934 -6147
rect 84007 -6152 85278 -6147
rect 87351 -6152 88622 -6147
rect 90695 -6152 91966 -6147
rect 94039 -6152 95310 -6147
rect 97383 -6152 98654 -6147
rect 100727 -6152 101998 -6147
rect 104071 -6152 104488 -6147
rect 3875 -6170 5022 -6152
rect 7219 -6170 8366 -6152
rect 10563 -6170 11710 -6152
rect 13907 -6170 15054 -6152
rect 17251 -6170 18398 -6152
rect 20595 -6170 21742 -6152
rect 23939 -6170 25086 -6152
rect 27283 -6170 28430 -6152
rect 30627 -6170 31774 -6152
rect 33971 -6170 35118 -6152
rect 37315 -6170 38462 -6152
rect 40659 -6170 41806 -6152
rect 44003 -6170 45150 -6152
rect 47347 -6170 48494 -6152
rect 50691 -6170 51838 -6152
rect 54035 -6170 55182 -6152
rect 57379 -6170 58526 -6152
rect 60723 -6170 61870 -6152
rect 64067 -6170 65214 -6152
rect 67411 -6170 68558 -6152
rect 70755 -6170 71902 -6152
rect 74099 -6170 75246 -6152
rect 77443 -6170 78590 -6152
rect 80787 -6170 81934 -6152
rect 84131 -6170 85278 -6152
rect 87475 -6170 88622 -6152
rect 90819 -6170 91966 -6152
rect 94163 -6170 95310 -6152
rect 97507 -6170 98654 -6152
rect 100851 -6170 101998 -6152
rect 104195 -6170 104633 -6152
rect 4313 -6181 5022 -6170
rect 7657 -6181 8366 -6170
rect 11001 -6181 11710 -6170
rect 14345 -6181 15054 -6170
rect 17689 -6181 18398 -6170
rect 21033 -6181 21742 -6170
rect 24377 -6181 25086 -6170
rect 27721 -6181 28430 -6170
rect 31065 -6181 31774 -6170
rect 34409 -6181 35118 -6170
rect 37753 -6181 38462 -6170
rect 41097 -6181 41806 -6170
rect 44441 -6181 45150 -6170
rect 47785 -6181 48494 -6170
rect 51129 -6181 51838 -6170
rect 54473 -6181 55182 -6170
rect 57817 -6181 58526 -6170
rect 61161 -6181 61870 -6170
rect 64505 -6181 65214 -6170
rect 67849 -6181 68558 -6170
rect 71193 -6181 71902 -6170
rect 74537 -6181 75246 -6170
rect 77881 -6181 78590 -6170
rect 81225 -6181 81934 -6170
rect 84569 -6181 85278 -6170
rect 87913 -6181 88622 -6170
rect 91257 -6181 91966 -6170
rect 94601 -6181 95310 -6170
rect 97945 -6181 98654 -6170
rect 101289 -6181 101998 -6170
rect 4313 -6217 4987 -6181
rect 7657 -6217 8331 -6181
rect 11001 -6217 11675 -6181
rect 14345 -6217 15019 -6181
rect 17689 -6217 18363 -6181
rect 21033 -6217 21707 -6181
rect 24377 -6217 25051 -6181
rect 27721 -6217 28395 -6181
rect 31065 -6217 31739 -6181
rect 34409 -6217 35083 -6181
rect 37753 -6217 38427 -6181
rect 41097 -6217 41771 -6181
rect 44441 -6217 45115 -6181
rect 47785 -6217 48459 -6181
rect 51129 -6217 51803 -6181
rect 54473 -6217 55147 -6181
rect 57817 -6217 58491 -6181
rect 61161 -6217 61835 -6181
rect 64505 -6217 65179 -6181
rect 67849 -6217 68523 -6181
rect 71193 -6217 71867 -6181
rect 74537 -6217 75211 -6181
rect 77881 -6217 78555 -6181
rect 81225 -6217 81899 -6181
rect 84569 -6217 85243 -6181
rect 87913 -6217 88587 -6181
rect 91257 -6217 91931 -6181
rect 94601 -6217 95275 -6181
rect 97945 -6217 98619 -6181
rect 101289 -6217 101963 -6181
rect 105289 -6181 105342 -5067
rect 111272 -4943 111475 -4848
rect 113465 -4906 114819 -4848
rect 116809 -4906 118163 -4848
rect 120153 -4906 121507 -4848
rect 123497 -4906 124851 -4848
rect 126841 -4906 128195 -4848
rect 130185 -4906 131539 -4848
rect 133529 -4906 134883 -4848
rect 136873 -4906 138227 -4848
rect 140217 -4906 141571 -4848
rect 143561 -4906 144915 -4848
rect 146905 -4906 148259 -4848
rect 150249 -4906 151603 -4848
rect 153593 -4906 154947 -4848
rect 156937 -4906 158291 -4848
rect 160281 -4906 161635 -4848
rect 163625 -4906 164979 -4848
rect 166969 -4906 168323 -4848
rect 170313 -4906 171667 -4848
rect 173657 -4906 175011 -4848
rect 177001 -4906 178355 -4848
rect 180345 -4906 181699 -4848
rect 183689 -4906 185043 -4848
rect 187033 -4906 188387 -4848
rect 190377 -4906 191731 -4848
rect 193721 -4906 195075 -4848
rect 197065 -4906 198419 -4848
rect 200409 -4906 201763 -4848
rect 203753 -4906 205107 -4848
rect 207097 -4906 208451 -4848
rect 210441 -4906 211795 -4848
rect 213785 -4906 215139 -4848
rect 112892 -4943 114819 -4906
rect 116236 -4943 118163 -4906
rect 119580 -4943 121507 -4906
rect 122924 -4943 124851 -4906
rect 126268 -4943 128195 -4906
rect 129612 -4943 131539 -4906
rect 132956 -4943 134883 -4906
rect 136300 -4943 138227 -4906
rect 139644 -4943 141571 -4906
rect 142988 -4943 144915 -4906
rect 146332 -4943 148259 -4906
rect 149676 -4943 151603 -4906
rect 153020 -4943 154947 -4906
rect 156364 -4943 158291 -4906
rect 159708 -4943 161635 -4906
rect 163052 -4943 164979 -4906
rect 166396 -4943 168323 -4906
rect 169740 -4943 171667 -4906
rect 173084 -4943 175011 -4906
rect 176428 -4943 178355 -4906
rect 179772 -4943 181699 -4906
rect 183116 -4943 185043 -4906
rect 186460 -4943 188387 -4906
rect 189804 -4943 191731 -4906
rect 193148 -4943 195075 -4906
rect 196492 -4943 198419 -4906
rect 199836 -4943 201763 -4906
rect 203180 -4943 205107 -4906
rect 206524 -4943 208451 -4906
rect 209868 -4943 211795 -4906
rect 213212 -4943 215139 -4906
rect 111272 -5067 111977 -4943
rect 112892 -5067 115321 -4943
rect 116236 -5067 118665 -4943
rect 119580 -5067 122009 -4943
rect 122924 -5067 125353 -4943
rect 126268 -5067 128697 -4943
rect 129612 -5067 132041 -4943
rect 132956 -5067 135385 -4943
rect 136300 -5067 138729 -4943
rect 139644 -5067 142073 -4943
rect 142988 -5067 145417 -4943
rect 146332 -5067 148761 -4943
rect 149676 -5067 152105 -4943
rect 153020 -5067 155449 -4943
rect 156364 -5067 158793 -4943
rect 159708 -5067 162137 -4943
rect 163052 -5067 165481 -4943
rect 166396 -5067 168825 -4943
rect 169740 -5067 172169 -4943
rect 173084 -5067 175513 -4943
rect 176428 -5067 178857 -4943
rect 179772 -5067 182201 -4943
rect 183116 -5067 185545 -4943
rect 186460 -5067 188889 -4943
rect 189804 -5067 192233 -4943
rect 193148 -5067 195577 -4943
rect 196492 -5067 198921 -4943
rect 199836 -5067 202265 -4943
rect 203180 -5067 205609 -4943
rect 206524 -5067 208953 -4943
rect 209868 -5067 212297 -4943
rect 213212 -5067 215641 -4943
rect 111272 -6152 112030 -5067
rect 112892 -6022 115374 -5067
rect 116236 -6022 118718 -5067
rect 119580 -6022 122062 -5067
rect 122924 -6022 125406 -5067
rect 126268 -6022 128750 -5067
rect 129612 -6022 132094 -5067
rect 132956 -6022 135438 -5067
rect 136300 -6022 138782 -5067
rect 139644 -6022 142126 -5067
rect 142988 -6022 145470 -5067
rect 146332 -6022 148814 -5067
rect 149676 -6022 152158 -5067
rect 153020 -6022 155502 -5067
rect 156364 -6022 158846 -5067
rect 159708 -6022 162190 -5067
rect 163052 -6022 165534 -5067
rect 166396 -6022 168878 -5067
rect 169740 -6022 172222 -5067
rect 173084 -6022 175566 -5067
rect 176428 -6022 178910 -5067
rect 179772 -6022 182254 -5067
rect 183116 -6022 185598 -5067
rect 186460 -6022 188942 -5067
rect 189804 -6022 192286 -5067
rect 193148 -6022 195630 -5067
rect 196492 -6022 198974 -5067
rect 199836 -6022 202318 -5067
rect 203180 -6022 205662 -5067
rect 206524 -6022 209006 -5067
rect 209868 -6022 212350 -5067
rect 213212 -6022 215694 -5067
rect 113483 -6087 115374 -6022
rect 116827 -6087 118718 -6022
rect 120171 -6087 122062 -6022
rect 123515 -6087 125406 -6022
rect 126859 -6087 128750 -6022
rect 130203 -6087 132094 -6022
rect 133547 -6087 135438 -6022
rect 136891 -6087 138782 -6022
rect 140235 -6087 142126 -6022
rect 143579 -6087 145470 -6022
rect 146923 -6087 148814 -6022
rect 150267 -6087 152158 -6022
rect 153611 -6087 155502 -6022
rect 156955 -6087 158846 -6022
rect 160299 -6087 162190 -6022
rect 163643 -6087 165534 -6022
rect 166987 -6087 168878 -6022
rect 170331 -6087 172222 -6022
rect 173675 -6087 175566 -6022
rect 177019 -6087 178910 -6022
rect 180363 -6087 182254 -6022
rect 183707 -6087 185598 -6022
rect 187051 -6087 188942 -6022
rect 190395 -6087 192286 -6022
rect 193739 -6087 195630 -6022
rect 197083 -6087 198974 -6022
rect 200427 -6087 202318 -6022
rect 203771 -6087 205662 -6022
rect 207115 -6087 209006 -6022
rect 210459 -6087 212350 -6022
rect 213803 -6087 215694 -6022
rect 114074 -6147 115374 -6087
rect 117418 -6147 118718 -6087
rect 120762 -6147 122062 -6087
rect 124106 -6147 125406 -6087
rect 127450 -6147 128750 -6087
rect 130794 -6147 132094 -6087
rect 134138 -6147 135438 -6087
rect 137482 -6147 138782 -6087
rect 140826 -6147 142126 -6087
rect 144170 -6147 145470 -6087
rect 147514 -6147 148814 -6087
rect 150858 -6147 152158 -6087
rect 154202 -6147 155502 -6087
rect 157546 -6147 158846 -6087
rect 160890 -6147 162190 -6087
rect 164234 -6147 165534 -6087
rect 167578 -6147 168878 -6087
rect 170922 -6147 172222 -6087
rect 174266 -6147 175566 -6087
rect 177610 -6147 178910 -6087
rect 180954 -6147 182254 -6087
rect 184298 -6147 185598 -6087
rect 187642 -6147 188942 -6087
rect 190986 -6147 192286 -6087
rect 194330 -6147 195630 -6087
rect 197674 -6147 198974 -6087
rect 201018 -6147 202318 -6087
rect 204362 -6147 205662 -6087
rect 207706 -6147 209006 -6087
rect 211050 -6147 212350 -6087
rect 214394 -6147 215694 -6087
rect 114103 -6152 115374 -6147
rect 117447 -6152 118718 -6147
rect 120791 -6152 122062 -6147
rect 124135 -6152 125406 -6147
rect 127479 -6152 128750 -6147
rect 130823 -6152 132094 -6147
rect 134167 -6152 135438 -6147
rect 137511 -6152 138782 -6147
rect 140855 -6152 142126 -6147
rect 144199 -6152 145470 -6147
rect 147543 -6152 148814 -6147
rect 150887 -6152 152158 -6147
rect 154231 -6152 155502 -6147
rect 157575 -6152 158846 -6147
rect 160919 -6152 162190 -6147
rect 164263 -6152 165534 -6147
rect 167607 -6152 168878 -6147
rect 170951 -6152 172222 -6147
rect 174295 -6152 175566 -6147
rect 177639 -6152 178910 -6147
rect 180983 -6152 182254 -6147
rect 184327 -6152 185598 -6147
rect 187671 -6152 188942 -6147
rect 191015 -6152 192286 -6147
rect 194359 -6152 195630 -6147
rect 197703 -6152 198974 -6147
rect 201047 -6152 202318 -6147
rect 204391 -6152 205662 -6147
rect 207735 -6152 209006 -6147
rect 211079 -6152 212350 -6147
rect 214423 -6152 215694 -6147
rect 110883 -6170 112030 -6152
rect 114227 -6170 115374 -6152
rect 117571 -6170 118718 -6152
rect 120915 -6170 122062 -6152
rect 124259 -6170 125406 -6152
rect 127603 -6170 128750 -6152
rect 130947 -6170 132094 -6152
rect 134291 -6170 135438 -6152
rect 137635 -6170 138782 -6152
rect 140979 -6170 142126 -6152
rect 144323 -6170 145470 -6152
rect 147667 -6170 148814 -6152
rect 151011 -6170 152158 -6152
rect 154355 -6170 155502 -6152
rect 157699 -6170 158846 -6152
rect 161043 -6170 162190 -6152
rect 164387 -6170 165534 -6152
rect 167731 -6170 168878 -6152
rect 171075 -6170 172222 -6152
rect 174419 -6170 175566 -6152
rect 177763 -6170 178910 -6152
rect 181107 -6170 182254 -6152
rect 184451 -6170 185598 -6152
rect 187795 -6170 188942 -6152
rect 191139 -6170 192286 -6152
rect 194483 -6170 195630 -6152
rect 197827 -6170 198974 -6152
rect 201171 -6170 202318 -6152
rect 204515 -6170 205662 -6152
rect 207859 -6170 209006 -6152
rect 211203 -6170 212350 -6152
rect 214547 -6170 215694 -6152
rect 111321 -6181 112030 -6170
rect 114665 -6181 115374 -6170
rect 118009 -6181 118718 -6170
rect 121353 -6181 122062 -6170
rect 124697 -6181 125406 -6170
rect 128041 -6181 128750 -6170
rect 131385 -6181 132094 -6170
rect 134729 -6181 135438 -6170
rect 138073 -6181 138782 -6170
rect 141417 -6181 142126 -6170
rect 144761 -6181 145470 -6170
rect 148105 -6181 148814 -6170
rect 151449 -6181 152158 -6170
rect 154793 -6181 155502 -6170
rect 158137 -6181 158846 -6170
rect 161481 -6181 162190 -6170
rect 164825 -6181 165534 -6170
rect 168169 -6181 168878 -6170
rect 171513 -6181 172222 -6170
rect 174857 -6181 175566 -6170
rect 178201 -6181 178910 -6170
rect 181545 -6181 182254 -6170
rect 184889 -6181 185598 -6170
rect 188233 -6181 188942 -6170
rect 191577 -6181 192286 -6170
rect 194921 -6181 195630 -6170
rect 198265 -6181 198974 -6170
rect 201609 -6181 202318 -6170
rect 204953 -6181 205662 -6170
rect 208297 -6181 209006 -6170
rect 211641 -6181 212350 -6170
rect 214985 -6181 215694 -6170
rect 105289 -6217 105307 -6181
rect 111321 -6217 111995 -6181
rect 114665 -6217 115339 -6181
rect 118009 -6217 118683 -6181
rect 121353 -6217 122027 -6181
rect 124697 -6217 125371 -6181
rect 128041 -6217 128715 -6181
rect 131385 -6217 132059 -6181
rect 134729 -6217 135403 -6181
rect 138073 -6217 138747 -6181
rect 141417 -6217 142091 -6181
rect 144761 -6217 145435 -6181
rect 148105 -6217 148779 -6181
rect 151449 -6217 152123 -6181
rect 154793 -6217 155467 -6181
rect 158137 -6217 158811 -6181
rect 161481 -6217 162155 -6181
rect 164825 -6217 165499 -6181
rect 168169 -6217 168843 -6181
rect 171513 -6217 172187 -6181
rect 174857 -6217 175531 -6181
rect 178201 -6217 178875 -6181
rect 181545 -6217 182219 -6181
rect 184889 -6217 185563 -6181
rect 188233 -6217 188907 -6181
rect 191577 -6217 192251 -6181
rect 194921 -6217 195595 -6181
rect 198265 -6217 198939 -6181
rect 201609 -6217 202283 -6181
rect 204953 -6217 205627 -6181
rect 208297 -6217 208971 -6181
rect 211641 -6217 212315 -6181
rect 214985 -6217 215659 -6181
rect 4496 -6235 4987 -6217
rect 7840 -6235 8331 -6217
rect 11184 -6235 11675 -6217
rect 14528 -6235 15019 -6217
rect 17872 -6235 18363 -6217
rect 21216 -6235 21707 -6217
rect 24560 -6235 25051 -6217
rect 27904 -6235 28395 -6217
rect 31248 -6235 31739 -6217
rect 34592 -6235 35083 -6217
rect 37936 -6235 38427 -6217
rect 41280 -6235 41771 -6217
rect 44624 -6235 45115 -6217
rect 47968 -6235 48459 -6217
rect 51312 -6235 51803 -6217
rect 54656 -6235 55147 -6217
rect 58000 -6235 58491 -6217
rect 61344 -6235 61835 -6217
rect 64688 -6235 65179 -6217
rect 68032 -6235 68523 -6217
rect 71376 -6235 71867 -6217
rect 74720 -6235 75211 -6217
rect 78064 -6235 78555 -6217
rect 81408 -6235 81899 -6217
rect 84752 -6235 85243 -6217
rect 88096 -6235 88587 -6217
rect 91440 -6235 91931 -6217
rect 94784 -6235 95275 -6217
rect 98128 -6235 98619 -6217
rect 101472 -6235 101963 -6217
rect 104816 -6235 105307 -6217
rect 111504 -6235 111995 -6217
rect 114848 -6235 115339 -6217
rect 118192 -6235 118683 -6217
rect 121536 -6235 122027 -6217
rect 124880 -6235 125371 -6217
rect 128224 -6235 128715 -6217
rect 131568 -6235 132059 -6217
rect 134912 -6235 135403 -6217
rect 138256 -6235 138747 -6217
rect 141600 -6235 142091 -6217
rect 144944 -6235 145435 -6217
rect 148288 -6235 148779 -6217
rect 151632 -6235 152123 -6217
rect 154976 -6235 155467 -6217
rect 158320 -6235 158811 -6217
rect 161664 -6235 162155 -6217
rect 165008 -6235 165499 -6217
rect 168352 -6235 168843 -6217
rect 171696 -6235 172187 -6217
rect 175040 -6235 175531 -6217
rect 178384 -6235 178875 -6217
rect 181728 -6235 182219 -6217
rect 185072 -6235 185563 -6217
rect 188416 -6235 188907 -6217
rect 191760 -6235 192251 -6217
rect 195104 -6235 195595 -6217
rect 198448 -6235 198939 -6217
rect 201792 -6235 202283 -6217
rect 205136 -6235 205627 -6217
rect 208480 -6235 208971 -6217
rect 211824 -6235 212315 -6217
rect 215168 -6235 215659 -6217
<< error_s >>
rect 107008 -2965 107124 -2899
rect 107124 -3219 107510 -3153
rect 106860 -3232 106870 -3219
rect 106794 -3274 106870 -3232
rect 106922 -3274 107510 -3219
rect 106794 -3277 107510 -3274
rect 106794 -3514 106938 -3277
rect 107124 -3299 107510 -3277
rect 107048 -3385 107510 -3299
rect 107052 -3393 107252 -3385
rect 107068 -3397 107236 -3393
rect 106794 -3600 106968 -3514
rect 106994 -3574 107094 -3450
rect 106994 -3628 106996 -3574
rect 106679 -4371 106823 -4324
rect 106860 -4371 106877 -4270
rect 106679 -4382 107451 -4371
rect 106765 -4407 107451 -4382
rect 106777 -4436 107451 -4407
rect 106777 -4848 107510 -4436
rect 107959 -4848 108006 -4483
rect 108013 -4848 108060 -4537
rect 106777 -4906 108131 -4848
rect 106204 -4943 108131 -4906
rect 106204 -5067 108633 -4943
rect 106204 -6022 108686 -5067
rect 109548 -6022 110012 -4906
rect 106795 -6087 108686 -6022
rect 107386 -6147 108686 -6087
rect 107415 -6152 108686 -6147
rect 107539 -6170 108686 -6152
rect 107977 -6181 108686 -6170
rect 107977 -6217 108651 -6181
rect 108160 -6235 108651 -6217
<< error_ps >>
rect 110138 -3514 110282 -3274
rect 110468 -3299 110854 -3153
rect 110392 -3385 110854 -3299
rect 110138 -3600 110312 -3514
rect 2540 -6022 2720 -4906
rect 104488 -4943 104787 -4848
rect 110139 -4436 110795 -4371
rect 110139 -4848 110854 -4436
rect 110139 -4906 111272 -4848
rect 104488 -6152 105289 -4943
rect 104633 -6217 105289 -6152
rect 110012 -6022 111272 -4906
rect 110139 -6087 111272 -6022
rect 110730 -6147 111272 -6087
rect 110759 -6152 111272 -6147
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use icell32scs  x1
timestamp 1717439242
transform 1 0 0 0 1 0
box 0 -6337 108752 458
use icell32scs  x2
timestamp 1717439242
transform 1 0 107008 0 1 0
box 0 -6337 108752 458
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
