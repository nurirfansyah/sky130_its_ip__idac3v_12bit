magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 3344 -2965 3460 -2899
rect 6688 -2965 6804 -2899
rect 10032 -2965 10148 -2899
rect 13376 -2965 13492 -2899
rect 16720 -2965 16836 -2899
rect 20064 -2965 20180 -2899
rect 23408 -2965 23524 -2899
rect 26752 -2965 26868 -2899
rect 30096 -2965 30212 -2899
rect 33440 -2965 33556 -2899
rect 36784 -2965 36900 -2899
rect 40128 -2965 40244 -2899
rect 43472 -2965 43588 -2899
rect 46816 -2965 46932 -2899
rect 50160 -2965 50276 -2899
rect 53504 -2965 53620 -2899
rect 56848 -2965 56964 -2899
rect 60192 -2965 60308 -2899
rect 63536 -2965 63652 -2899
rect 66880 -2965 66996 -2899
rect 70224 -2965 70340 -2899
rect 73568 -2965 73684 -2899
rect 76912 -2965 77028 -2899
rect 80256 -2965 80372 -2899
rect 83600 -2965 83716 -2899
rect 86944 -2965 87060 -2899
rect 90288 -2965 90404 -2899
rect 93632 -2965 93748 -2899
rect 96976 -2965 97092 -2899
rect 100320 -2965 100436 -2899
rect 103664 -2965 103780 -2899
rect 107008 -2965 107124 -2899
rect 110352 -2965 110468 -2899
rect 113696 -2965 113812 -2899
rect 117040 -2965 117156 -2899
rect 120384 -2965 120500 -2899
rect 123728 -2965 123844 -2899
rect 127072 -2965 127188 -2899
rect 130416 -2965 130532 -2899
rect 133760 -2965 133876 -2899
rect 137104 -2965 137220 -2899
rect 140448 -2965 140564 -2899
rect 143792 -2965 143908 -2899
rect 147136 -2965 147252 -2899
rect 150480 -2965 150596 -2899
rect 153824 -2965 153940 -2899
rect 157168 -2965 157284 -2899
rect 160512 -2965 160628 -2899
rect 163856 -2965 163972 -2899
rect 167200 -2965 167316 -2899
rect 170544 -2965 170660 -2899
rect 173888 -2965 174004 -2899
rect 177232 -2965 177348 -2899
rect 180576 -2965 180692 -2899
rect 183920 -2965 184036 -2899
rect 187264 -2965 187380 -2899
rect 190608 -2965 190724 -2899
rect 193952 -2965 194068 -2899
rect 197296 -2965 197412 -2899
rect 200640 -2965 200756 -2899
rect 203984 -2965 204100 -2899
rect 207328 -2965 207444 -2899
rect 210672 -2965 210788 -2899
rect 217360 -2965 217476 -2899
rect 220704 -2965 220820 -2899
rect 224048 -2965 224164 -2899
rect 227392 -2965 227508 -2899
rect 230736 -2965 230852 -2899
rect 234080 -2965 234196 -2899
rect 237424 -2965 237540 -2899
rect 240768 -2965 240884 -2899
rect 244112 -2965 244228 -2899
rect 247456 -2965 247572 -2899
rect 250800 -2965 250916 -2899
rect 254144 -2965 254260 -2899
rect 257488 -2965 257604 -2899
rect 260832 -2965 260948 -2899
rect 264176 -2965 264292 -2899
rect 267520 -2965 267636 -2899
rect 270864 -2965 270980 -2899
rect 274208 -2965 274324 -2899
rect 277552 -2965 277668 -2899
rect 280896 -2965 281012 -2899
rect 284240 -2965 284356 -2899
rect 287584 -2965 287700 -2899
rect 290928 -2965 291044 -2899
rect 294272 -2965 294388 -2899
rect 297616 -2965 297732 -2899
rect 300960 -2965 301076 -2899
rect 304304 -2965 304420 -2899
rect 307648 -2965 307764 -2899
rect 310992 -2965 311108 -2899
rect 314336 -2965 314452 -2899
rect 317680 -2965 317796 -2899
rect 321024 -2965 321140 -2899
rect 324368 -2965 324484 -2899
rect 327712 -2965 327828 -2899
rect 331056 -2965 331172 -2899
rect 334400 -2965 334516 -2899
rect 337744 -2965 337860 -2899
rect 341088 -2965 341204 -2899
rect 344432 -2965 344548 -2899
rect 347776 -2965 347892 -2899
rect 351120 -2965 351236 -2899
rect 354464 -2965 354580 -2899
rect 357808 -2965 357924 -2899
rect 361152 -2965 361268 -2899
rect 364496 -2965 364612 -2899
rect 367840 -2965 367956 -2899
rect 371184 -2965 371300 -2899
rect 374528 -2965 374644 -2899
rect 377872 -2965 377988 -2899
rect 381216 -2965 381332 -2899
rect 384560 -2965 384676 -2899
rect 387904 -2965 388020 -2899
rect 391248 -2965 391364 -2899
rect 394592 -2965 394708 -2899
rect 397936 -2965 398052 -2899
rect 401280 -2965 401396 -2899
rect 404624 -2965 404740 -2899
rect 407968 -2965 408084 -2899
rect 411312 -2965 411428 -2899
rect 414656 -2965 414772 -2899
rect 418000 -2965 418116 -2899
rect 421344 -2965 421460 -2899
rect 424688 -2965 424804 -2899
rect 3460 -3219 3846 -3153
rect 6804 -3219 7190 -3153
rect 10148 -3219 10534 -3153
rect 13492 -3219 13878 -3153
rect 16836 -3219 17222 -3153
rect 20180 -3219 20566 -3153
rect 23524 -3219 23910 -3153
rect 26868 -3219 27254 -3153
rect 30212 -3219 30598 -3153
rect 33556 -3219 33942 -3153
rect 36900 -3219 37286 -3153
rect 40244 -3219 40630 -3153
rect 43588 -3219 43974 -3153
rect 46932 -3219 47318 -3153
rect 50276 -3219 50662 -3153
rect 53620 -3219 54006 -3153
rect 56964 -3219 57350 -3153
rect 60308 -3219 60694 -3153
rect 63652 -3219 64038 -3153
rect 66996 -3219 67382 -3153
rect 70340 -3219 70726 -3153
rect 73684 -3219 74070 -3153
rect 77028 -3219 77414 -3153
rect 80372 -3219 80758 -3153
rect 83716 -3219 84102 -3153
rect 87060 -3219 87446 -3153
rect 90404 -3219 90790 -3153
rect 93748 -3219 94134 -3153
rect 97092 -3219 97478 -3153
rect 100436 -3219 100822 -3153
rect 103780 -3219 104166 -3153
rect 107124 -3219 107510 -3153
rect 110468 -3219 110854 -3153
rect 113812 -3219 114198 -3153
rect 117156 -3219 117542 -3153
rect 120500 -3219 120886 -3153
rect 123844 -3219 124230 -3153
rect 127188 -3219 127574 -3153
rect 130532 -3219 130918 -3153
rect 133876 -3219 134262 -3153
rect 137220 -3219 137606 -3153
rect 140564 -3219 140950 -3153
rect 143908 -3219 144294 -3153
rect 147252 -3219 147638 -3153
rect 150596 -3219 150982 -3153
rect 153940 -3219 154326 -3153
rect 157284 -3219 157670 -3153
rect 160628 -3219 161014 -3153
rect 163972 -3219 164358 -3153
rect 167316 -3219 167702 -3153
rect 170660 -3219 171046 -3153
rect 174004 -3219 174390 -3153
rect 177348 -3219 177734 -3153
rect 180692 -3219 181078 -3153
rect 184036 -3219 184422 -3153
rect 187380 -3219 187766 -3153
rect 190724 -3219 191110 -3153
rect 194068 -3219 194454 -3153
rect 197412 -3219 197798 -3153
rect 200756 -3219 201142 -3153
rect 204100 -3219 204486 -3153
rect 207444 -3219 207830 -3153
rect 210788 -3219 211174 -3153
rect 3196 -3232 3206 -3219
rect 3130 -3274 3206 -3232
rect 3258 -3274 3846 -3219
rect 6540 -3232 6550 -3219
rect 3130 -3277 3846 -3274
rect 3130 -3514 3274 -3277
rect 3460 -3299 3846 -3277
rect 3384 -3385 3846 -3299
rect 6474 -3274 6550 -3232
rect 6602 -3274 7190 -3219
rect 9884 -3232 9894 -3219
rect 6474 -3277 7190 -3274
rect 3388 -3393 3588 -3385
rect 3404 -3397 3572 -3393
rect 3130 -3600 3304 -3514
rect 3330 -3574 3430 -3450
rect 6474 -3514 6618 -3277
rect 6804 -3299 7190 -3277
rect 6728 -3385 7190 -3299
rect 9818 -3274 9894 -3232
rect 9946 -3274 10534 -3219
rect 13228 -3232 13238 -3219
rect 9818 -3277 10534 -3274
rect 6732 -3393 6932 -3385
rect 6748 -3397 6916 -3393
rect 3330 -3628 3332 -3574
rect 6474 -3600 6648 -3514
rect 6674 -3574 6774 -3450
rect 9818 -3514 9962 -3277
rect 10148 -3299 10534 -3277
rect 10072 -3385 10534 -3299
rect 13162 -3274 13238 -3232
rect 13290 -3274 13878 -3219
rect 16572 -3232 16582 -3219
rect 13162 -3277 13878 -3274
rect 10076 -3393 10276 -3385
rect 10092 -3397 10260 -3393
rect 6674 -3628 6676 -3574
rect 9818 -3600 9992 -3514
rect 10018 -3574 10118 -3450
rect 13162 -3514 13306 -3277
rect 13492 -3299 13878 -3277
rect 13416 -3385 13878 -3299
rect 16506 -3274 16582 -3232
rect 16634 -3274 17222 -3219
rect 19916 -3232 19926 -3219
rect 16506 -3277 17222 -3274
rect 13420 -3393 13620 -3385
rect 13436 -3397 13604 -3393
rect 10018 -3628 10020 -3574
rect 13162 -3600 13336 -3514
rect 13362 -3574 13462 -3450
rect 16506 -3514 16650 -3277
rect 16836 -3299 17222 -3277
rect 16760 -3385 17222 -3299
rect 19850 -3274 19926 -3232
rect 19978 -3274 20566 -3219
rect 23260 -3232 23270 -3219
rect 19850 -3277 20566 -3274
rect 16764 -3393 16964 -3385
rect 16780 -3397 16948 -3393
rect 13362 -3628 13364 -3574
rect 16506 -3600 16680 -3514
rect 16706 -3574 16806 -3450
rect 19850 -3514 19994 -3277
rect 20180 -3299 20566 -3277
rect 20104 -3385 20566 -3299
rect 23194 -3274 23270 -3232
rect 23322 -3274 23910 -3219
rect 26604 -3232 26614 -3219
rect 23194 -3277 23910 -3274
rect 20108 -3393 20308 -3385
rect 20124 -3397 20292 -3393
rect 16706 -3628 16708 -3574
rect 19850 -3600 20024 -3514
rect 20050 -3574 20150 -3450
rect 23194 -3514 23338 -3277
rect 23524 -3299 23910 -3277
rect 23448 -3385 23910 -3299
rect 26538 -3274 26614 -3232
rect 26666 -3274 27254 -3219
rect 29948 -3232 29958 -3219
rect 26538 -3277 27254 -3274
rect 23452 -3393 23652 -3385
rect 23468 -3397 23636 -3393
rect 20050 -3628 20052 -3574
rect 23194 -3600 23368 -3514
rect 23394 -3574 23494 -3450
rect 26538 -3514 26682 -3277
rect 26868 -3299 27254 -3277
rect 26792 -3385 27254 -3299
rect 29882 -3274 29958 -3232
rect 30010 -3274 30598 -3219
rect 33292 -3232 33302 -3219
rect 29882 -3277 30598 -3274
rect 26796 -3393 26996 -3385
rect 26812 -3397 26980 -3393
rect 23394 -3628 23396 -3574
rect 26538 -3600 26712 -3514
rect 26738 -3574 26838 -3450
rect 29882 -3514 30026 -3277
rect 30212 -3299 30598 -3277
rect 30136 -3385 30598 -3299
rect 33226 -3274 33302 -3232
rect 33354 -3274 33942 -3219
rect 36636 -3232 36646 -3219
rect 33226 -3277 33942 -3274
rect 30140 -3393 30340 -3385
rect 30156 -3397 30324 -3393
rect 26738 -3628 26740 -3574
rect 29882 -3600 30056 -3514
rect 30082 -3574 30182 -3450
rect 33226 -3514 33370 -3277
rect 33556 -3299 33942 -3277
rect 33480 -3385 33942 -3299
rect 36570 -3274 36646 -3232
rect 36698 -3274 37286 -3219
rect 39980 -3232 39990 -3219
rect 36570 -3277 37286 -3274
rect 33484 -3393 33684 -3385
rect 33500 -3397 33668 -3393
rect 30082 -3628 30084 -3574
rect 33226 -3600 33400 -3514
rect 33426 -3574 33526 -3450
rect 36570 -3514 36714 -3277
rect 36900 -3299 37286 -3277
rect 36824 -3385 37286 -3299
rect 39914 -3274 39990 -3232
rect 40042 -3274 40630 -3219
rect 43324 -3232 43334 -3219
rect 39914 -3277 40630 -3274
rect 36828 -3393 37028 -3385
rect 36844 -3397 37012 -3393
rect 33426 -3628 33428 -3574
rect 36570 -3600 36744 -3514
rect 36770 -3574 36870 -3450
rect 39914 -3514 40058 -3277
rect 40244 -3299 40630 -3277
rect 40168 -3385 40630 -3299
rect 43258 -3274 43334 -3232
rect 43386 -3274 43974 -3219
rect 46668 -3232 46678 -3219
rect 43258 -3277 43974 -3274
rect 40172 -3393 40372 -3385
rect 40188 -3397 40356 -3393
rect 36770 -3628 36772 -3574
rect 39914 -3600 40088 -3514
rect 40114 -3574 40214 -3450
rect 43258 -3514 43402 -3277
rect 43588 -3299 43974 -3277
rect 43512 -3385 43974 -3299
rect 46602 -3274 46678 -3232
rect 46730 -3274 47318 -3219
rect 50012 -3232 50022 -3219
rect 46602 -3277 47318 -3274
rect 43516 -3393 43716 -3385
rect 43532 -3397 43700 -3393
rect 40114 -3628 40116 -3574
rect 43258 -3600 43432 -3514
rect 43458 -3574 43558 -3450
rect 46602 -3514 46746 -3277
rect 46932 -3299 47318 -3277
rect 46856 -3385 47318 -3299
rect 49946 -3274 50022 -3232
rect 50074 -3274 50662 -3219
rect 53356 -3232 53366 -3219
rect 49946 -3277 50662 -3274
rect 46860 -3393 47060 -3385
rect 46876 -3397 47044 -3393
rect 43458 -3628 43460 -3574
rect 46602 -3600 46776 -3514
rect 46802 -3574 46902 -3450
rect 49946 -3514 50090 -3277
rect 50276 -3299 50662 -3277
rect 50200 -3385 50662 -3299
rect 53290 -3274 53366 -3232
rect 53418 -3274 54006 -3219
rect 56700 -3232 56710 -3219
rect 53290 -3277 54006 -3274
rect 50204 -3393 50404 -3385
rect 50220 -3397 50388 -3393
rect 46802 -3628 46804 -3574
rect 49946 -3600 50120 -3514
rect 50146 -3574 50246 -3450
rect 53290 -3514 53434 -3277
rect 53620 -3299 54006 -3277
rect 53544 -3385 54006 -3299
rect 56634 -3274 56710 -3232
rect 56762 -3274 57350 -3219
rect 60044 -3232 60054 -3219
rect 56634 -3277 57350 -3274
rect 53548 -3393 53748 -3385
rect 53564 -3397 53732 -3393
rect 50146 -3628 50148 -3574
rect 53290 -3600 53464 -3514
rect 53490 -3574 53590 -3450
rect 56634 -3514 56778 -3277
rect 56964 -3299 57350 -3277
rect 56888 -3385 57350 -3299
rect 59978 -3274 60054 -3232
rect 60106 -3274 60694 -3219
rect 63388 -3232 63398 -3219
rect 59978 -3277 60694 -3274
rect 56892 -3393 57092 -3385
rect 56908 -3397 57076 -3393
rect 53490 -3628 53492 -3574
rect 56634 -3600 56808 -3514
rect 56834 -3574 56934 -3450
rect 59978 -3514 60122 -3277
rect 60308 -3299 60694 -3277
rect 60232 -3385 60694 -3299
rect 63322 -3274 63398 -3232
rect 63450 -3274 64038 -3219
rect 66732 -3232 66742 -3219
rect 63322 -3277 64038 -3274
rect 60236 -3393 60436 -3385
rect 60252 -3397 60420 -3393
rect 56834 -3628 56836 -3574
rect 59978 -3600 60152 -3514
rect 60178 -3574 60278 -3450
rect 63322 -3514 63466 -3277
rect 63652 -3299 64038 -3277
rect 63576 -3385 64038 -3299
rect 66666 -3274 66742 -3232
rect 66794 -3274 67382 -3219
rect 70076 -3232 70086 -3219
rect 66666 -3277 67382 -3274
rect 63580 -3393 63780 -3385
rect 63596 -3397 63764 -3393
rect 60178 -3628 60180 -3574
rect 63322 -3600 63496 -3514
rect 63522 -3574 63622 -3450
rect 66666 -3514 66810 -3277
rect 66996 -3299 67382 -3277
rect 66920 -3385 67382 -3299
rect 70010 -3274 70086 -3232
rect 70138 -3274 70726 -3219
rect 73420 -3232 73430 -3219
rect 70010 -3277 70726 -3274
rect 66924 -3393 67124 -3385
rect 66940 -3397 67108 -3393
rect 63522 -3628 63524 -3574
rect 66666 -3600 66840 -3514
rect 66866 -3574 66966 -3450
rect 70010 -3514 70154 -3277
rect 70340 -3299 70726 -3277
rect 70264 -3385 70726 -3299
rect 73354 -3274 73430 -3232
rect 73482 -3274 74070 -3219
rect 76764 -3232 76774 -3219
rect 73354 -3277 74070 -3274
rect 70268 -3393 70468 -3385
rect 70284 -3397 70452 -3393
rect 66866 -3628 66868 -3574
rect 70010 -3600 70184 -3514
rect 70210 -3574 70310 -3450
rect 73354 -3514 73498 -3277
rect 73684 -3299 74070 -3277
rect 73608 -3385 74070 -3299
rect 76698 -3274 76774 -3232
rect 76826 -3274 77414 -3219
rect 80108 -3232 80118 -3219
rect 76698 -3277 77414 -3274
rect 73612 -3393 73812 -3385
rect 73628 -3397 73796 -3393
rect 70210 -3628 70212 -3574
rect 73354 -3600 73528 -3514
rect 73554 -3574 73654 -3450
rect 76698 -3514 76842 -3277
rect 77028 -3299 77414 -3277
rect 76952 -3385 77414 -3299
rect 80042 -3274 80118 -3232
rect 80170 -3274 80758 -3219
rect 83452 -3232 83462 -3219
rect 80042 -3277 80758 -3274
rect 76956 -3393 77156 -3385
rect 76972 -3397 77140 -3393
rect 73554 -3628 73556 -3574
rect 76698 -3600 76872 -3514
rect 76898 -3574 76998 -3450
rect 80042 -3514 80186 -3277
rect 80372 -3299 80758 -3277
rect 80296 -3385 80758 -3299
rect 83386 -3274 83462 -3232
rect 83514 -3274 84102 -3219
rect 86796 -3232 86806 -3219
rect 83386 -3277 84102 -3274
rect 80300 -3393 80500 -3385
rect 80316 -3397 80484 -3393
rect 76898 -3628 76900 -3574
rect 80042 -3600 80216 -3514
rect 80242 -3574 80342 -3450
rect 83386 -3514 83530 -3277
rect 83716 -3299 84102 -3277
rect 83640 -3385 84102 -3299
rect 86730 -3274 86806 -3232
rect 86858 -3274 87446 -3219
rect 90140 -3232 90150 -3219
rect 86730 -3277 87446 -3274
rect 83644 -3393 83844 -3385
rect 83660 -3397 83828 -3393
rect 80242 -3628 80244 -3574
rect 83386 -3600 83560 -3514
rect 83586 -3574 83686 -3450
rect 86730 -3514 86874 -3277
rect 87060 -3299 87446 -3277
rect 86984 -3385 87446 -3299
rect 90074 -3274 90150 -3232
rect 90202 -3274 90790 -3219
rect 93484 -3232 93494 -3219
rect 90074 -3277 90790 -3274
rect 86988 -3393 87188 -3385
rect 87004 -3397 87172 -3393
rect 83586 -3628 83588 -3574
rect 86730 -3600 86904 -3514
rect 86930 -3574 87030 -3450
rect 90074 -3514 90218 -3277
rect 90404 -3299 90790 -3277
rect 90328 -3385 90790 -3299
rect 93418 -3274 93494 -3232
rect 93546 -3274 94134 -3219
rect 96828 -3232 96838 -3219
rect 93418 -3277 94134 -3274
rect 90332 -3393 90532 -3385
rect 90348 -3397 90516 -3393
rect 86930 -3628 86932 -3574
rect 90074 -3600 90248 -3514
rect 90274 -3574 90374 -3450
rect 93418 -3514 93562 -3277
rect 93748 -3299 94134 -3277
rect 93672 -3385 94134 -3299
rect 96762 -3274 96838 -3232
rect 96890 -3274 97478 -3219
rect 100172 -3232 100182 -3219
rect 96762 -3277 97478 -3274
rect 93676 -3393 93876 -3385
rect 93692 -3397 93860 -3393
rect 90274 -3628 90276 -3574
rect 93418 -3600 93592 -3514
rect 93618 -3574 93718 -3450
rect 96762 -3514 96906 -3277
rect 97092 -3299 97478 -3277
rect 97016 -3385 97478 -3299
rect 100106 -3274 100182 -3232
rect 100234 -3274 100822 -3219
rect 103516 -3232 103526 -3219
rect 100106 -3277 100822 -3274
rect 97020 -3393 97220 -3385
rect 97036 -3397 97204 -3393
rect 93618 -3628 93620 -3574
rect 96762 -3600 96936 -3514
rect 96962 -3574 97062 -3450
rect 100106 -3514 100250 -3277
rect 100436 -3299 100822 -3277
rect 100360 -3385 100822 -3299
rect 103450 -3274 103526 -3232
rect 103578 -3274 104166 -3219
rect 106860 -3232 106870 -3219
rect 103450 -3277 104166 -3274
rect 100364 -3393 100564 -3385
rect 100380 -3397 100548 -3393
rect 96962 -3628 96964 -3574
rect 100106 -3600 100280 -3514
rect 100306 -3574 100406 -3450
rect 103450 -3514 103594 -3277
rect 103780 -3299 104166 -3277
rect 103704 -3385 104166 -3299
rect 106794 -3274 106870 -3232
rect 106922 -3274 107510 -3219
rect 110204 -3232 110214 -3219
rect 106794 -3277 107510 -3274
rect 103708 -3393 103908 -3385
rect 103724 -3397 103892 -3393
rect 100306 -3628 100308 -3574
rect 103450 -3600 103624 -3514
rect 103650 -3574 103750 -3450
rect 106794 -3514 106938 -3277
rect 107124 -3299 107510 -3277
rect 107048 -3385 107510 -3299
rect 110138 -3274 110214 -3232
rect 110266 -3274 110854 -3219
rect 113548 -3232 113558 -3219
rect 110138 -3277 110854 -3274
rect 107052 -3393 107252 -3385
rect 107068 -3397 107236 -3393
rect 103650 -3628 103652 -3574
rect 106794 -3600 106968 -3514
rect 106994 -3574 107094 -3450
rect 110138 -3514 110282 -3277
rect 110468 -3299 110854 -3277
rect 110392 -3385 110854 -3299
rect 113482 -3274 113558 -3232
rect 113610 -3274 114198 -3219
rect 116892 -3232 116902 -3219
rect 113482 -3277 114198 -3274
rect 110396 -3393 110596 -3385
rect 110412 -3397 110580 -3393
rect 106994 -3628 106996 -3574
rect 110138 -3600 110312 -3514
rect 110338 -3574 110438 -3450
rect 113482 -3514 113626 -3277
rect 113812 -3299 114198 -3277
rect 113736 -3385 114198 -3299
rect 116826 -3274 116902 -3232
rect 116954 -3274 117542 -3219
rect 120236 -3232 120246 -3219
rect 116826 -3277 117542 -3274
rect 113740 -3393 113940 -3385
rect 113756 -3397 113924 -3393
rect 110338 -3628 110340 -3574
rect 113482 -3600 113656 -3514
rect 113682 -3574 113782 -3450
rect 116826 -3514 116970 -3277
rect 117156 -3299 117542 -3277
rect 117080 -3385 117542 -3299
rect 120170 -3274 120246 -3232
rect 120298 -3274 120886 -3219
rect 123580 -3232 123590 -3219
rect 120170 -3277 120886 -3274
rect 117084 -3393 117284 -3385
rect 117100 -3397 117268 -3393
rect 113682 -3628 113684 -3574
rect 116826 -3600 117000 -3514
rect 117026 -3574 117126 -3450
rect 120170 -3514 120314 -3277
rect 120500 -3299 120886 -3277
rect 120424 -3385 120886 -3299
rect 123514 -3274 123590 -3232
rect 123642 -3274 124230 -3219
rect 126924 -3232 126934 -3219
rect 123514 -3277 124230 -3274
rect 120428 -3393 120628 -3385
rect 120444 -3397 120612 -3393
rect 117026 -3628 117028 -3574
rect 120170 -3600 120344 -3514
rect 120370 -3574 120470 -3450
rect 123514 -3514 123658 -3277
rect 123844 -3299 124230 -3277
rect 123768 -3385 124230 -3299
rect 126858 -3274 126934 -3232
rect 126986 -3274 127574 -3219
rect 130268 -3232 130278 -3219
rect 126858 -3277 127574 -3274
rect 123772 -3393 123972 -3385
rect 123788 -3397 123956 -3393
rect 120370 -3628 120372 -3574
rect 123514 -3600 123688 -3514
rect 123714 -3574 123814 -3450
rect 126858 -3514 127002 -3277
rect 127188 -3299 127574 -3277
rect 127112 -3385 127574 -3299
rect 130202 -3274 130278 -3232
rect 130330 -3274 130918 -3219
rect 133612 -3232 133622 -3219
rect 130202 -3277 130918 -3274
rect 127116 -3393 127316 -3385
rect 127132 -3397 127300 -3393
rect 123714 -3628 123716 -3574
rect 126858 -3600 127032 -3514
rect 127058 -3574 127158 -3450
rect 130202 -3514 130346 -3277
rect 130532 -3299 130918 -3277
rect 130456 -3385 130918 -3299
rect 133546 -3274 133622 -3232
rect 133674 -3274 134262 -3219
rect 136956 -3232 136966 -3219
rect 133546 -3277 134262 -3274
rect 130460 -3393 130660 -3385
rect 130476 -3397 130644 -3393
rect 127058 -3628 127060 -3574
rect 130202 -3600 130376 -3514
rect 130402 -3574 130502 -3450
rect 133546 -3514 133690 -3277
rect 133876 -3299 134262 -3277
rect 133800 -3385 134262 -3299
rect 136890 -3274 136966 -3232
rect 137018 -3274 137606 -3219
rect 140300 -3232 140310 -3219
rect 136890 -3277 137606 -3274
rect 133804 -3393 134004 -3385
rect 133820 -3397 133988 -3393
rect 130402 -3628 130404 -3574
rect 133546 -3600 133720 -3514
rect 133746 -3574 133846 -3450
rect 136890 -3514 137034 -3277
rect 137220 -3299 137606 -3277
rect 137144 -3385 137606 -3299
rect 140234 -3274 140310 -3232
rect 140362 -3274 140950 -3219
rect 143644 -3232 143654 -3219
rect 140234 -3277 140950 -3274
rect 137148 -3393 137348 -3385
rect 137164 -3397 137332 -3393
rect 133746 -3628 133748 -3574
rect 136890 -3600 137064 -3514
rect 137090 -3574 137190 -3450
rect 140234 -3514 140378 -3277
rect 140564 -3299 140950 -3277
rect 140488 -3385 140950 -3299
rect 143578 -3274 143654 -3232
rect 143706 -3274 144294 -3219
rect 146988 -3232 146998 -3219
rect 143578 -3277 144294 -3274
rect 140492 -3393 140692 -3385
rect 140508 -3397 140676 -3393
rect 137090 -3628 137092 -3574
rect 140234 -3600 140408 -3514
rect 140434 -3574 140534 -3450
rect 143578 -3514 143722 -3277
rect 143908 -3299 144294 -3277
rect 143832 -3385 144294 -3299
rect 146922 -3274 146998 -3232
rect 147050 -3274 147638 -3219
rect 150332 -3232 150342 -3219
rect 146922 -3277 147638 -3274
rect 143836 -3393 144036 -3385
rect 143852 -3397 144020 -3393
rect 140434 -3628 140436 -3574
rect 143578 -3600 143752 -3514
rect 143778 -3574 143878 -3450
rect 146922 -3514 147066 -3277
rect 147252 -3299 147638 -3277
rect 147176 -3385 147638 -3299
rect 150266 -3274 150342 -3232
rect 150394 -3274 150982 -3219
rect 153676 -3232 153686 -3219
rect 150266 -3277 150982 -3274
rect 147180 -3393 147380 -3385
rect 147196 -3397 147364 -3393
rect 143778 -3628 143780 -3574
rect 146922 -3600 147096 -3514
rect 147122 -3574 147222 -3450
rect 150266 -3514 150410 -3277
rect 150596 -3299 150982 -3277
rect 150520 -3385 150982 -3299
rect 153610 -3274 153686 -3232
rect 153738 -3274 154326 -3219
rect 157020 -3232 157030 -3219
rect 153610 -3277 154326 -3274
rect 150524 -3393 150724 -3385
rect 150540 -3397 150708 -3393
rect 147122 -3628 147124 -3574
rect 150266 -3600 150440 -3514
rect 150466 -3574 150566 -3450
rect 153610 -3514 153754 -3277
rect 153940 -3299 154326 -3277
rect 153864 -3385 154326 -3299
rect 156954 -3274 157030 -3232
rect 157082 -3274 157670 -3219
rect 160364 -3232 160374 -3219
rect 156954 -3277 157670 -3274
rect 153868 -3393 154068 -3385
rect 153884 -3397 154052 -3393
rect 150466 -3628 150468 -3574
rect 153610 -3600 153784 -3514
rect 153810 -3574 153910 -3450
rect 156954 -3514 157098 -3277
rect 157284 -3299 157670 -3277
rect 157208 -3385 157670 -3299
rect 160298 -3274 160374 -3232
rect 160426 -3274 161014 -3219
rect 163708 -3232 163718 -3219
rect 160298 -3277 161014 -3274
rect 157212 -3393 157412 -3385
rect 157228 -3397 157396 -3393
rect 153810 -3628 153812 -3574
rect 156954 -3600 157128 -3514
rect 157154 -3574 157254 -3450
rect 160298 -3514 160442 -3277
rect 160628 -3299 161014 -3277
rect 160552 -3385 161014 -3299
rect 163642 -3274 163718 -3232
rect 163770 -3274 164358 -3219
rect 167052 -3232 167062 -3219
rect 163642 -3277 164358 -3274
rect 160556 -3393 160756 -3385
rect 160572 -3397 160740 -3393
rect 157154 -3628 157156 -3574
rect 160298 -3600 160472 -3514
rect 160498 -3574 160598 -3450
rect 163642 -3514 163786 -3277
rect 163972 -3299 164358 -3277
rect 163896 -3385 164358 -3299
rect 166986 -3274 167062 -3232
rect 167114 -3274 167702 -3219
rect 170396 -3232 170406 -3219
rect 166986 -3277 167702 -3274
rect 163900 -3393 164100 -3385
rect 163916 -3397 164084 -3393
rect 160498 -3628 160500 -3574
rect 163642 -3600 163816 -3514
rect 163842 -3574 163942 -3450
rect 166986 -3514 167130 -3277
rect 167316 -3299 167702 -3277
rect 167240 -3385 167702 -3299
rect 170330 -3274 170406 -3232
rect 170458 -3274 171046 -3219
rect 173740 -3232 173750 -3219
rect 170330 -3277 171046 -3274
rect 167244 -3393 167444 -3385
rect 167260 -3397 167428 -3393
rect 163842 -3628 163844 -3574
rect 166986 -3600 167160 -3514
rect 167186 -3574 167286 -3450
rect 170330 -3514 170474 -3277
rect 170660 -3299 171046 -3277
rect 170584 -3385 171046 -3299
rect 173674 -3274 173750 -3232
rect 173802 -3274 174390 -3219
rect 177084 -3232 177094 -3219
rect 173674 -3277 174390 -3274
rect 170588 -3393 170788 -3385
rect 170604 -3397 170772 -3393
rect 167186 -3628 167188 -3574
rect 170330 -3600 170504 -3514
rect 170530 -3574 170630 -3450
rect 173674 -3514 173818 -3277
rect 174004 -3299 174390 -3277
rect 173928 -3385 174390 -3299
rect 177018 -3274 177094 -3232
rect 177146 -3274 177734 -3219
rect 180428 -3232 180438 -3219
rect 177018 -3277 177734 -3274
rect 173932 -3393 174132 -3385
rect 173948 -3397 174116 -3393
rect 170530 -3628 170532 -3574
rect 173674 -3600 173848 -3514
rect 173874 -3574 173974 -3450
rect 177018 -3514 177162 -3277
rect 177348 -3299 177734 -3277
rect 177272 -3385 177734 -3299
rect 180362 -3274 180438 -3232
rect 180490 -3274 181078 -3219
rect 183772 -3232 183782 -3219
rect 180362 -3277 181078 -3274
rect 177276 -3393 177476 -3385
rect 177292 -3397 177460 -3393
rect 173874 -3628 173876 -3574
rect 177018 -3600 177192 -3514
rect 177218 -3574 177318 -3450
rect 180362 -3514 180506 -3277
rect 180692 -3299 181078 -3277
rect 180616 -3385 181078 -3299
rect 183706 -3274 183782 -3232
rect 183834 -3274 184422 -3219
rect 187116 -3232 187126 -3219
rect 183706 -3277 184422 -3274
rect 180620 -3393 180820 -3385
rect 180636 -3397 180804 -3393
rect 177218 -3628 177220 -3574
rect 180362 -3600 180536 -3514
rect 180562 -3574 180662 -3450
rect 183706 -3514 183850 -3277
rect 184036 -3299 184422 -3277
rect 183960 -3385 184422 -3299
rect 187050 -3274 187126 -3232
rect 187178 -3274 187766 -3219
rect 190460 -3232 190470 -3219
rect 187050 -3277 187766 -3274
rect 183964 -3393 184164 -3385
rect 183980 -3397 184148 -3393
rect 180562 -3628 180564 -3574
rect 183706 -3600 183880 -3514
rect 183906 -3574 184006 -3450
rect 187050 -3514 187194 -3277
rect 187380 -3299 187766 -3277
rect 187304 -3385 187766 -3299
rect 190394 -3274 190470 -3232
rect 190522 -3274 191110 -3219
rect 193804 -3232 193814 -3219
rect 190394 -3277 191110 -3274
rect 187308 -3393 187508 -3385
rect 187324 -3397 187492 -3393
rect 183906 -3628 183908 -3574
rect 187050 -3600 187224 -3514
rect 187250 -3574 187350 -3450
rect 190394 -3514 190538 -3277
rect 190724 -3299 191110 -3277
rect 190648 -3385 191110 -3299
rect 193738 -3274 193814 -3232
rect 193866 -3274 194454 -3219
rect 197148 -3232 197158 -3219
rect 193738 -3277 194454 -3274
rect 190652 -3393 190852 -3385
rect 190668 -3397 190836 -3393
rect 187250 -3628 187252 -3574
rect 190394 -3600 190568 -3514
rect 190594 -3574 190694 -3450
rect 193738 -3514 193882 -3277
rect 194068 -3299 194454 -3277
rect 193992 -3385 194454 -3299
rect 197082 -3274 197158 -3232
rect 197210 -3274 197798 -3219
rect 200492 -3232 200502 -3219
rect 197082 -3277 197798 -3274
rect 193996 -3393 194196 -3385
rect 194012 -3397 194180 -3393
rect 190594 -3628 190596 -3574
rect 193738 -3600 193912 -3514
rect 193938 -3574 194038 -3450
rect 197082 -3514 197226 -3277
rect 197412 -3299 197798 -3277
rect 197336 -3385 197798 -3299
rect 200426 -3274 200502 -3232
rect 200554 -3274 201142 -3219
rect 203836 -3232 203846 -3219
rect 200426 -3277 201142 -3274
rect 197340 -3393 197540 -3385
rect 197356 -3397 197524 -3393
rect 193938 -3628 193940 -3574
rect 197082 -3600 197256 -3514
rect 197282 -3574 197382 -3450
rect 200426 -3514 200570 -3277
rect 200756 -3299 201142 -3277
rect 200680 -3385 201142 -3299
rect 203770 -3274 203846 -3232
rect 203898 -3274 204486 -3219
rect 207180 -3232 207190 -3219
rect 203770 -3277 204486 -3274
rect 200684 -3393 200884 -3385
rect 200700 -3397 200868 -3393
rect 197282 -3628 197284 -3574
rect 200426 -3600 200600 -3514
rect 200626 -3574 200726 -3450
rect 203770 -3514 203914 -3277
rect 204100 -3299 204486 -3277
rect 204024 -3385 204486 -3299
rect 207114 -3274 207190 -3232
rect 207242 -3274 207830 -3219
rect 210524 -3232 210534 -3219
rect 207114 -3277 207830 -3274
rect 204028 -3393 204228 -3385
rect 204044 -3397 204212 -3393
rect 200626 -3628 200628 -3574
rect 203770 -3600 203944 -3514
rect 203970 -3574 204070 -3450
rect 207114 -3514 207258 -3277
rect 207444 -3299 207830 -3277
rect 207368 -3385 207830 -3299
rect 210458 -3274 210534 -3232
rect 210586 -3274 211174 -3219
rect 210458 -3277 211174 -3274
rect 207372 -3393 207572 -3385
rect 207388 -3397 207556 -3393
rect 203970 -3628 203972 -3574
rect 207114 -3600 207288 -3514
rect 207314 -3574 207414 -3450
rect 210458 -3514 210602 -3277
rect 210788 -3299 211174 -3277
rect 210712 -3385 211174 -3299
rect 217212 -3232 217222 -3219
rect 210716 -3393 210916 -3385
rect 210732 -3397 210900 -3393
rect 207314 -3628 207316 -3574
rect 210458 -3600 210632 -3514
rect 210658 -3574 210758 -3450
rect 217146 -3274 217222 -3232
rect 217274 -3274 217476 -3219
rect 210658 -3628 210660 -3574
rect 217290 -3277 217476 -3274
rect 220820 -3219 221206 -3153
rect 224164 -3219 224550 -3153
rect 227508 -3219 227894 -3153
rect 230852 -3219 231238 -3153
rect 234196 -3219 234582 -3153
rect 237540 -3219 237926 -3153
rect 240884 -3219 241270 -3153
rect 244228 -3219 244614 -3153
rect 247572 -3219 247958 -3153
rect 250916 -3219 251302 -3153
rect 254260 -3219 254646 -3153
rect 257604 -3219 257990 -3153
rect 260948 -3219 261334 -3153
rect 264292 -3219 264678 -3153
rect 267636 -3219 268022 -3153
rect 270980 -3219 271366 -3153
rect 274324 -3219 274710 -3153
rect 277668 -3219 278054 -3153
rect 281012 -3219 281398 -3153
rect 284356 -3219 284742 -3153
rect 287700 -3219 288086 -3153
rect 291044 -3219 291430 -3153
rect 294388 -3219 294774 -3153
rect 297732 -3219 298118 -3153
rect 301076 -3219 301462 -3153
rect 304420 -3219 304806 -3153
rect 307764 -3219 308150 -3153
rect 311108 -3219 311494 -3153
rect 314452 -3219 314838 -3153
rect 317796 -3219 318182 -3153
rect 321140 -3219 321526 -3153
rect 324484 -3219 324870 -3153
rect 327828 -3219 328214 -3153
rect 331172 -3219 331558 -3153
rect 334516 -3219 334902 -3153
rect 337860 -3219 338246 -3153
rect 341204 -3219 341590 -3153
rect 344548 -3219 344934 -3153
rect 347892 -3219 348278 -3153
rect 351236 -3219 351622 -3153
rect 354580 -3219 354966 -3153
rect 357924 -3219 358310 -3153
rect 361268 -3219 361654 -3153
rect 364612 -3219 364998 -3153
rect 367956 -3219 368342 -3153
rect 371300 -3219 371686 -3153
rect 374644 -3219 375030 -3153
rect 377988 -3219 378374 -3153
rect 381332 -3219 381718 -3153
rect 384676 -3219 385062 -3153
rect 388020 -3219 388406 -3153
rect 391364 -3219 391750 -3153
rect 394708 -3219 395094 -3153
rect 398052 -3219 398438 -3153
rect 401396 -3219 401782 -3153
rect 404740 -3219 405126 -3153
rect 408084 -3219 408470 -3153
rect 411428 -3219 411814 -3153
rect 414772 -3219 415158 -3153
rect 418116 -3219 418502 -3153
rect 421460 -3219 421846 -3153
rect 424804 -3219 425190 -3153
rect 220556 -3232 220566 -3219
rect 220490 -3274 220566 -3232
rect 220618 -3274 221206 -3219
rect 223900 -3232 223910 -3219
rect 220490 -3277 221206 -3274
rect 217404 -3393 217604 -3385
rect 217420 -3397 217588 -3393
rect 217346 -3574 217446 -3450
rect 220490 -3514 220634 -3277
rect 220820 -3299 221206 -3277
rect 220744 -3385 221206 -3299
rect 223834 -3274 223910 -3232
rect 223962 -3274 224550 -3219
rect 227244 -3232 227254 -3219
rect 223834 -3277 224550 -3274
rect 220748 -3393 220948 -3385
rect 220764 -3397 220932 -3393
rect 217346 -3628 217348 -3574
rect 220490 -3600 220664 -3514
rect 220690 -3574 220790 -3450
rect 223834 -3514 223978 -3277
rect 224164 -3299 224550 -3277
rect 224088 -3385 224550 -3299
rect 227178 -3274 227254 -3232
rect 227306 -3274 227894 -3219
rect 230588 -3232 230598 -3219
rect 227178 -3277 227894 -3274
rect 224092 -3393 224292 -3385
rect 224108 -3397 224276 -3393
rect 220690 -3628 220692 -3574
rect 223834 -3600 224008 -3514
rect 224034 -3574 224134 -3450
rect 227178 -3514 227322 -3277
rect 227508 -3299 227894 -3277
rect 227432 -3385 227894 -3299
rect 230522 -3274 230598 -3232
rect 230650 -3274 231238 -3219
rect 233932 -3232 233942 -3219
rect 230522 -3277 231238 -3274
rect 227436 -3393 227636 -3385
rect 227452 -3397 227620 -3393
rect 224034 -3628 224036 -3574
rect 227178 -3600 227352 -3514
rect 227378 -3574 227478 -3450
rect 230522 -3514 230666 -3277
rect 230852 -3299 231238 -3277
rect 230776 -3385 231238 -3299
rect 233866 -3274 233942 -3232
rect 233994 -3274 234582 -3219
rect 237276 -3232 237286 -3219
rect 233866 -3277 234582 -3274
rect 230780 -3393 230980 -3385
rect 230796 -3397 230964 -3393
rect 227378 -3628 227380 -3574
rect 230522 -3600 230696 -3514
rect 230722 -3574 230822 -3450
rect 233866 -3514 234010 -3277
rect 234196 -3299 234582 -3277
rect 234120 -3385 234582 -3299
rect 237210 -3274 237286 -3232
rect 237338 -3274 237926 -3219
rect 240620 -3232 240630 -3219
rect 237210 -3277 237926 -3274
rect 234124 -3393 234324 -3385
rect 234140 -3397 234308 -3393
rect 230722 -3628 230724 -3574
rect 233866 -3600 234040 -3514
rect 234066 -3574 234166 -3450
rect 237210 -3514 237354 -3277
rect 237540 -3299 237926 -3277
rect 237464 -3385 237926 -3299
rect 240554 -3274 240630 -3232
rect 240682 -3274 241270 -3219
rect 243964 -3232 243974 -3219
rect 240554 -3277 241270 -3274
rect 237468 -3393 237668 -3385
rect 237484 -3397 237652 -3393
rect 234066 -3628 234068 -3574
rect 237210 -3600 237384 -3514
rect 237410 -3574 237510 -3450
rect 240554 -3514 240698 -3277
rect 240884 -3299 241270 -3277
rect 240808 -3385 241270 -3299
rect 243898 -3274 243974 -3232
rect 244026 -3274 244614 -3219
rect 247308 -3232 247318 -3219
rect 243898 -3277 244614 -3274
rect 240812 -3393 241012 -3385
rect 240828 -3397 240996 -3393
rect 237410 -3628 237412 -3574
rect 240554 -3600 240728 -3514
rect 240754 -3574 240854 -3450
rect 243898 -3514 244042 -3277
rect 244228 -3299 244614 -3277
rect 244152 -3385 244614 -3299
rect 247242 -3274 247318 -3232
rect 247370 -3274 247958 -3219
rect 250652 -3232 250662 -3219
rect 247242 -3277 247958 -3274
rect 244156 -3393 244356 -3385
rect 244172 -3397 244340 -3393
rect 240754 -3628 240756 -3574
rect 243898 -3600 244072 -3514
rect 244098 -3574 244198 -3450
rect 247242 -3514 247386 -3277
rect 247572 -3299 247958 -3277
rect 247496 -3385 247958 -3299
rect 250586 -3274 250662 -3232
rect 250714 -3274 251302 -3219
rect 253996 -3232 254006 -3219
rect 250586 -3277 251302 -3274
rect 247500 -3393 247700 -3385
rect 247516 -3397 247684 -3393
rect 244098 -3628 244100 -3574
rect 247242 -3600 247416 -3514
rect 247442 -3574 247542 -3450
rect 250586 -3514 250730 -3277
rect 250916 -3299 251302 -3277
rect 250840 -3385 251302 -3299
rect 253930 -3274 254006 -3232
rect 254058 -3274 254646 -3219
rect 257340 -3232 257350 -3219
rect 253930 -3277 254646 -3274
rect 250844 -3393 251044 -3385
rect 250860 -3397 251028 -3393
rect 247442 -3628 247444 -3574
rect 250586 -3600 250760 -3514
rect 250786 -3574 250886 -3450
rect 253930 -3514 254074 -3277
rect 254260 -3299 254646 -3277
rect 254184 -3385 254646 -3299
rect 257274 -3274 257350 -3232
rect 257402 -3274 257990 -3219
rect 260684 -3232 260694 -3219
rect 257274 -3277 257990 -3274
rect 254188 -3393 254388 -3385
rect 254204 -3397 254372 -3393
rect 250786 -3628 250788 -3574
rect 253930 -3600 254104 -3514
rect 254130 -3574 254230 -3450
rect 257274 -3514 257418 -3277
rect 257604 -3299 257990 -3277
rect 257528 -3385 257990 -3299
rect 260618 -3274 260694 -3232
rect 260746 -3274 261334 -3219
rect 264028 -3232 264038 -3219
rect 260618 -3277 261334 -3274
rect 257532 -3393 257732 -3385
rect 257548 -3397 257716 -3393
rect 254130 -3628 254132 -3574
rect 257274 -3600 257448 -3514
rect 257474 -3574 257574 -3450
rect 260618 -3514 260762 -3277
rect 260948 -3299 261334 -3277
rect 260872 -3385 261334 -3299
rect 263962 -3274 264038 -3232
rect 264090 -3274 264678 -3219
rect 267372 -3232 267382 -3219
rect 263962 -3277 264678 -3274
rect 260876 -3393 261076 -3385
rect 260892 -3397 261060 -3393
rect 257474 -3628 257476 -3574
rect 260618 -3600 260792 -3514
rect 260818 -3574 260918 -3450
rect 263962 -3514 264106 -3277
rect 264292 -3299 264678 -3277
rect 264216 -3385 264678 -3299
rect 267306 -3274 267382 -3232
rect 267434 -3274 268022 -3219
rect 270716 -3232 270726 -3219
rect 267306 -3277 268022 -3274
rect 264220 -3393 264420 -3385
rect 264236 -3397 264404 -3393
rect 260818 -3628 260820 -3574
rect 263962 -3600 264136 -3514
rect 264162 -3574 264262 -3450
rect 267306 -3514 267450 -3277
rect 267636 -3299 268022 -3277
rect 267560 -3385 268022 -3299
rect 270650 -3274 270726 -3232
rect 270778 -3274 271366 -3219
rect 274060 -3232 274070 -3219
rect 270650 -3277 271366 -3274
rect 267564 -3393 267764 -3385
rect 267580 -3397 267748 -3393
rect 264162 -3628 264164 -3574
rect 267306 -3600 267480 -3514
rect 267506 -3574 267606 -3450
rect 270650 -3514 270794 -3277
rect 270980 -3299 271366 -3277
rect 270904 -3385 271366 -3299
rect 273994 -3274 274070 -3232
rect 274122 -3274 274710 -3219
rect 277404 -3232 277414 -3219
rect 273994 -3277 274710 -3274
rect 270908 -3393 271108 -3385
rect 270924 -3397 271092 -3393
rect 267506 -3628 267508 -3574
rect 270650 -3600 270824 -3514
rect 270850 -3574 270950 -3450
rect 273994 -3514 274138 -3277
rect 274324 -3299 274710 -3277
rect 274248 -3385 274710 -3299
rect 277338 -3274 277414 -3232
rect 277466 -3274 278054 -3219
rect 280748 -3232 280758 -3219
rect 277338 -3277 278054 -3274
rect 274252 -3393 274452 -3385
rect 274268 -3397 274436 -3393
rect 270850 -3628 270852 -3574
rect 273994 -3600 274168 -3514
rect 274194 -3574 274294 -3450
rect 277338 -3514 277482 -3277
rect 277668 -3299 278054 -3277
rect 277592 -3385 278054 -3299
rect 280682 -3274 280758 -3232
rect 280810 -3274 281398 -3219
rect 284092 -3232 284102 -3219
rect 280682 -3277 281398 -3274
rect 277596 -3393 277796 -3385
rect 277612 -3397 277780 -3393
rect 274194 -3628 274196 -3574
rect 277338 -3600 277512 -3514
rect 277538 -3574 277638 -3450
rect 280682 -3514 280826 -3277
rect 281012 -3299 281398 -3277
rect 280936 -3385 281398 -3299
rect 284026 -3274 284102 -3232
rect 284154 -3274 284742 -3219
rect 287436 -3232 287446 -3219
rect 284026 -3277 284742 -3274
rect 280940 -3393 281140 -3385
rect 280956 -3397 281124 -3393
rect 277538 -3628 277540 -3574
rect 280682 -3600 280856 -3514
rect 280882 -3574 280982 -3450
rect 284026 -3514 284170 -3277
rect 284356 -3299 284742 -3277
rect 284280 -3385 284742 -3299
rect 287370 -3274 287446 -3232
rect 287498 -3274 288086 -3219
rect 290780 -3232 290790 -3219
rect 287370 -3277 288086 -3274
rect 284284 -3393 284484 -3385
rect 284300 -3397 284468 -3393
rect 280882 -3628 280884 -3574
rect 284026 -3600 284200 -3514
rect 284226 -3574 284326 -3450
rect 287370 -3514 287514 -3277
rect 287700 -3299 288086 -3277
rect 287624 -3385 288086 -3299
rect 290714 -3274 290790 -3232
rect 290842 -3274 291430 -3219
rect 294124 -3232 294134 -3219
rect 290714 -3277 291430 -3274
rect 287628 -3393 287828 -3385
rect 287644 -3397 287812 -3393
rect 284226 -3628 284228 -3574
rect 287370 -3600 287544 -3514
rect 287570 -3574 287670 -3450
rect 290714 -3514 290858 -3277
rect 291044 -3299 291430 -3277
rect 290968 -3385 291430 -3299
rect 294058 -3274 294134 -3232
rect 294186 -3274 294774 -3219
rect 297468 -3232 297478 -3219
rect 294058 -3277 294774 -3274
rect 290972 -3393 291172 -3385
rect 290988 -3397 291156 -3393
rect 287570 -3628 287572 -3574
rect 290714 -3600 290888 -3514
rect 290914 -3574 291014 -3450
rect 294058 -3514 294202 -3277
rect 294388 -3299 294774 -3277
rect 294312 -3385 294774 -3299
rect 297402 -3274 297478 -3232
rect 297530 -3274 298118 -3219
rect 300812 -3232 300822 -3219
rect 297402 -3277 298118 -3274
rect 294316 -3393 294516 -3385
rect 294332 -3397 294500 -3393
rect 290914 -3628 290916 -3574
rect 294058 -3600 294232 -3514
rect 294258 -3574 294358 -3450
rect 297402 -3514 297546 -3277
rect 297732 -3299 298118 -3277
rect 297656 -3385 298118 -3299
rect 300746 -3274 300822 -3232
rect 300874 -3274 301462 -3219
rect 304156 -3232 304166 -3219
rect 300746 -3277 301462 -3274
rect 297660 -3393 297860 -3385
rect 297676 -3397 297844 -3393
rect 294258 -3628 294260 -3574
rect 297402 -3600 297576 -3514
rect 297602 -3574 297702 -3450
rect 300746 -3514 300890 -3277
rect 301076 -3299 301462 -3277
rect 301000 -3385 301462 -3299
rect 304090 -3274 304166 -3232
rect 304218 -3274 304806 -3219
rect 307500 -3232 307510 -3219
rect 304090 -3277 304806 -3274
rect 301004 -3393 301204 -3385
rect 301020 -3397 301188 -3393
rect 297602 -3628 297604 -3574
rect 300746 -3600 300920 -3514
rect 300946 -3574 301046 -3450
rect 304090 -3514 304234 -3277
rect 304420 -3299 304806 -3277
rect 304344 -3385 304806 -3299
rect 307434 -3274 307510 -3232
rect 307562 -3274 308150 -3219
rect 310844 -3232 310854 -3219
rect 307434 -3277 308150 -3274
rect 304348 -3393 304548 -3385
rect 304364 -3397 304532 -3393
rect 300946 -3628 300948 -3574
rect 304090 -3600 304264 -3514
rect 304290 -3574 304390 -3450
rect 307434 -3514 307578 -3277
rect 307764 -3299 308150 -3277
rect 307688 -3385 308150 -3299
rect 310778 -3274 310854 -3232
rect 310906 -3274 311494 -3219
rect 314188 -3232 314198 -3219
rect 310778 -3277 311494 -3274
rect 307692 -3393 307892 -3385
rect 307708 -3397 307876 -3393
rect 304290 -3628 304292 -3574
rect 307434 -3600 307608 -3514
rect 307634 -3574 307734 -3450
rect 310778 -3514 310922 -3277
rect 311108 -3299 311494 -3277
rect 311032 -3385 311494 -3299
rect 314122 -3274 314198 -3232
rect 314250 -3274 314838 -3219
rect 317532 -3232 317542 -3219
rect 314122 -3277 314838 -3274
rect 311036 -3393 311236 -3385
rect 311052 -3397 311220 -3393
rect 307634 -3628 307636 -3574
rect 310778 -3600 310952 -3514
rect 310978 -3574 311078 -3450
rect 314122 -3514 314266 -3277
rect 314452 -3299 314838 -3277
rect 314376 -3385 314838 -3299
rect 317466 -3274 317542 -3232
rect 317594 -3274 318182 -3219
rect 320876 -3232 320886 -3219
rect 317466 -3277 318182 -3274
rect 314380 -3393 314580 -3385
rect 314396 -3397 314564 -3393
rect 310978 -3628 310980 -3574
rect 314122 -3600 314296 -3514
rect 314322 -3574 314422 -3450
rect 317466 -3514 317610 -3277
rect 317796 -3299 318182 -3277
rect 317720 -3385 318182 -3299
rect 320810 -3274 320886 -3232
rect 320938 -3274 321526 -3219
rect 324220 -3232 324230 -3219
rect 320810 -3277 321526 -3274
rect 317724 -3393 317924 -3385
rect 317740 -3397 317908 -3393
rect 314322 -3628 314324 -3574
rect 317466 -3600 317640 -3514
rect 317666 -3574 317766 -3450
rect 320810 -3514 320954 -3277
rect 321140 -3299 321526 -3277
rect 321064 -3385 321526 -3299
rect 324154 -3274 324230 -3232
rect 324282 -3274 324870 -3219
rect 327564 -3232 327574 -3219
rect 324154 -3277 324870 -3274
rect 321068 -3393 321268 -3385
rect 321084 -3397 321252 -3393
rect 317666 -3628 317668 -3574
rect 320810 -3600 320984 -3514
rect 321010 -3574 321110 -3450
rect 324154 -3514 324298 -3277
rect 324484 -3299 324870 -3277
rect 324408 -3385 324870 -3299
rect 327498 -3274 327574 -3232
rect 327626 -3274 328214 -3219
rect 330908 -3232 330918 -3219
rect 327498 -3277 328214 -3274
rect 324412 -3393 324612 -3385
rect 324428 -3397 324596 -3393
rect 321010 -3628 321012 -3574
rect 324154 -3600 324328 -3514
rect 324354 -3574 324454 -3450
rect 327498 -3514 327642 -3277
rect 327828 -3299 328214 -3277
rect 327752 -3385 328214 -3299
rect 330842 -3274 330918 -3232
rect 330970 -3274 331558 -3219
rect 334252 -3232 334262 -3219
rect 330842 -3277 331558 -3274
rect 327756 -3393 327956 -3385
rect 327772 -3397 327940 -3393
rect 324354 -3628 324356 -3574
rect 327498 -3600 327672 -3514
rect 327698 -3574 327798 -3450
rect 330842 -3514 330986 -3277
rect 331172 -3299 331558 -3277
rect 331096 -3385 331558 -3299
rect 334186 -3274 334262 -3232
rect 334314 -3274 334902 -3219
rect 337596 -3232 337606 -3219
rect 334186 -3277 334902 -3274
rect 331100 -3393 331300 -3385
rect 331116 -3397 331284 -3393
rect 327698 -3628 327700 -3574
rect 330842 -3600 331016 -3514
rect 331042 -3574 331142 -3450
rect 334186 -3514 334330 -3277
rect 334516 -3299 334902 -3277
rect 334440 -3385 334902 -3299
rect 337530 -3274 337606 -3232
rect 337658 -3274 338246 -3219
rect 340940 -3232 340950 -3219
rect 337530 -3277 338246 -3274
rect 334444 -3393 334644 -3385
rect 334460 -3397 334628 -3393
rect 331042 -3628 331044 -3574
rect 334186 -3600 334360 -3514
rect 334386 -3574 334486 -3450
rect 337530 -3514 337674 -3277
rect 337860 -3299 338246 -3277
rect 337784 -3385 338246 -3299
rect 340874 -3274 340950 -3232
rect 341002 -3274 341590 -3219
rect 344284 -3232 344294 -3219
rect 340874 -3277 341590 -3274
rect 337788 -3393 337988 -3385
rect 337804 -3397 337972 -3393
rect 334386 -3628 334388 -3574
rect 337530 -3600 337704 -3514
rect 337730 -3574 337830 -3450
rect 340874 -3514 341018 -3277
rect 341204 -3299 341590 -3277
rect 341128 -3385 341590 -3299
rect 344218 -3274 344294 -3232
rect 344346 -3274 344934 -3219
rect 347628 -3232 347638 -3219
rect 344218 -3277 344934 -3274
rect 341132 -3393 341332 -3385
rect 341148 -3397 341316 -3393
rect 337730 -3628 337732 -3574
rect 340874 -3600 341048 -3514
rect 341074 -3574 341174 -3450
rect 344218 -3514 344362 -3277
rect 344548 -3299 344934 -3277
rect 344472 -3385 344934 -3299
rect 347562 -3274 347638 -3232
rect 347690 -3274 348278 -3219
rect 350972 -3232 350982 -3219
rect 347562 -3277 348278 -3274
rect 344476 -3393 344676 -3385
rect 344492 -3397 344660 -3393
rect 341074 -3628 341076 -3574
rect 344218 -3600 344392 -3514
rect 344418 -3574 344518 -3450
rect 347562 -3514 347706 -3277
rect 347892 -3299 348278 -3277
rect 347816 -3385 348278 -3299
rect 350906 -3274 350982 -3232
rect 351034 -3274 351622 -3219
rect 354316 -3232 354326 -3219
rect 350906 -3277 351622 -3274
rect 347820 -3393 348020 -3385
rect 347836 -3397 348004 -3393
rect 344418 -3628 344420 -3574
rect 347562 -3600 347736 -3514
rect 347762 -3574 347862 -3450
rect 350906 -3514 351050 -3277
rect 351236 -3299 351622 -3277
rect 351160 -3385 351622 -3299
rect 354250 -3274 354326 -3232
rect 354378 -3274 354966 -3219
rect 357660 -3232 357670 -3219
rect 354250 -3277 354966 -3274
rect 351164 -3393 351364 -3385
rect 351180 -3397 351348 -3393
rect 347762 -3628 347764 -3574
rect 350906 -3600 351080 -3514
rect 351106 -3574 351206 -3450
rect 354250 -3514 354394 -3277
rect 354580 -3299 354966 -3277
rect 354504 -3385 354966 -3299
rect 357594 -3274 357670 -3232
rect 357722 -3274 358310 -3219
rect 361004 -3232 361014 -3219
rect 357594 -3277 358310 -3274
rect 354508 -3393 354708 -3385
rect 354524 -3397 354692 -3393
rect 351106 -3628 351108 -3574
rect 354250 -3600 354424 -3514
rect 354450 -3574 354550 -3450
rect 357594 -3514 357738 -3277
rect 357924 -3299 358310 -3277
rect 357848 -3385 358310 -3299
rect 360938 -3274 361014 -3232
rect 361066 -3274 361654 -3219
rect 364348 -3232 364358 -3219
rect 360938 -3277 361654 -3274
rect 357852 -3393 358052 -3385
rect 357868 -3397 358036 -3393
rect 354450 -3628 354452 -3574
rect 357594 -3600 357768 -3514
rect 357794 -3574 357894 -3450
rect 360938 -3514 361082 -3277
rect 361268 -3299 361654 -3277
rect 361192 -3385 361654 -3299
rect 364282 -3274 364358 -3232
rect 364410 -3274 364998 -3219
rect 367692 -3232 367702 -3219
rect 364282 -3277 364998 -3274
rect 361196 -3393 361396 -3385
rect 361212 -3397 361380 -3393
rect 357794 -3628 357796 -3574
rect 360938 -3600 361112 -3514
rect 361138 -3574 361238 -3450
rect 364282 -3514 364426 -3277
rect 364612 -3299 364998 -3277
rect 364536 -3385 364998 -3299
rect 367626 -3274 367702 -3232
rect 367754 -3274 368342 -3219
rect 371036 -3232 371046 -3219
rect 367626 -3277 368342 -3274
rect 364540 -3393 364740 -3385
rect 364556 -3397 364724 -3393
rect 361138 -3628 361140 -3574
rect 364282 -3600 364456 -3514
rect 364482 -3574 364582 -3450
rect 367626 -3514 367770 -3277
rect 367956 -3299 368342 -3277
rect 367880 -3385 368342 -3299
rect 370970 -3274 371046 -3232
rect 371098 -3274 371686 -3219
rect 374380 -3232 374390 -3219
rect 370970 -3277 371686 -3274
rect 367884 -3393 368084 -3385
rect 367900 -3397 368068 -3393
rect 364482 -3628 364484 -3574
rect 367626 -3600 367800 -3514
rect 367826 -3574 367926 -3450
rect 370970 -3514 371114 -3277
rect 371300 -3299 371686 -3277
rect 371224 -3385 371686 -3299
rect 374314 -3274 374390 -3232
rect 374442 -3274 375030 -3219
rect 377724 -3232 377734 -3219
rect 374314 -3277 375030 -3274
rect 371228 -3393 371428 -3385
rect 371244 -3397 371412 -3393
rect 367826 -3628 367828 -3574
rect 370970 -3600 371144 -3514
rect 371170 -3574 371270 -3450
rect 374314 -3514 374458 -3277
rect 374644 -3299 375030 -3277
rect 374568 -3385 375030 -3299
rect 377658 -3274 377734 -3232
rect 377786 -3274 378374 -3219
rect 381068 -3232 381078 -3219
rect 377658 -3277 378374 -3274
rect 374572 -3393 374772 -3385
rect 374588 -3397 374756 -3393
rect 371170 -3628 371172 -3574
rect 374314 -3600 374488 -3514
rect 374514 -3574 374614 -3450
rect 377658 -3514 377802 -3277
rect 377988 -3299 378374 -3277
rect 377912 -3385 378374 -3299
rect 381002 -3274 381078 -3232
rect 381130 -3274 381718 -3219
rect 384412 -3232 384422 -3219
rect 381002 -3277 381718 -3274
rect 377916 -3393 378116 -3385
rect 377932 -3397 378100 -3393
rect 374514 -3628 374516 -3574
rect 377658 -3600 377832 -3514
rect 377858 -3574 377958 -3450
rect 381002 -3514 381146 -3277
rect 381332 -3299 381718 -3277
rect 381256 -3385 381718 -3299
rect 384346 -3274 384422 -3232
rect 384474 -3274 385062 -3219
rect 387756 -3232 387766 -3219
rect 384346 -3277 385062 -3274
rect 381260 -3393 381460 -3385
rect 381276 -3397 381444 -3393
rect 377858 -3628 377860 -3574
rect 381002 -3600 381176 -3514
rect 381202 -3574 381302 -3450
rect 384346 -3514 384490 -3277
rect 384676 -3299 385062 -3277
rect 384600 -3385 385062 -3299
rect 387690 -3274 387766 -3232
rect 387818 -3274 388406 -3219
rect 391100 -3232 391110 -3219
rect 387690 -3277 388406 -3274
rect 384604 -3393 384804 -3385
rect 384620 -3397 384788 -3393
rect 381202 -3628 381204 -3574
rect 384346 -3600 384520 -3514
rect 384546 -3574 384646 -3450
rect 387690 -3514 387834 -3277
rect 388020 -3299 388406 -3277
rect 387944 -3385 388406 -3299
rect 391034 -3274 391110 -3232
rect 391162 -3274 391750 -3219
rect 394444 -3232 394454 -3219
rect 391034 -3277 391750 -3274
rect 387948 -3393 388148 -3385
rect 387964 -3397 388132 -3393
rect 384546 -3628 384548 -3574
rect 387690 -3600 387864 -3514
rect 387890 -3574 387990 -3450
rect 391034 -3514 391178 -3277
rect 391364 -3299 391750 -3277
rect 391288 -3385 391750 -3299
rect 394378 -3274 394454 -3232
rect 394506 -3274 395094 -3219
rect 397788 -3232 397798 -3219
rect 394378 -3277 395094 -3274
rect 391292 -3393 391492 -3385
rect 391308 -3397 391476 -3393
rect 387890 -3628 387892 -3574
rect 391034 -3600 391208 -3514
rect 391234 -3574 391334 -3450
rect 394378 -3514 394522 -3277
rect 394708 -3299 395094 -3277
rect 394632 -3385 395094 -3299
rect 397722 -3274 397798 -3232
rect 397850 -3274 398438 -3219
rect 401132 -3232 401142 -3219
rect 397722 -3277 398438 -3274
rect 394636 -3393 394836 -3385
rect 394652 -3397 394820 -3393
rect 391234 -3628 391236 -3574
rect 394378 -3600 394552 -3514
rect 394578 -3574 394678 -3450
rect 397722 -3514 397866 -3277
rect 398052 -3299 398438 -3277
rect 397976 -3385 398438 -3299
rect 401066 -3274 401142 -3232
rect 401194 -3274 401782 -3219
rect 404476 -3232 404486 -3219
rect 401066 -3277 401782 -3274
rect 397980 -3393 398180 -3385
rect 397996 -3397 398164 -3393
rect 394578 -3628 394580 -3574
rect 397722 -3600 397896 -3514
rect 397922 -3574 398022 -3450
rect 401066 -3514 401210 -3277
rect 401396 -3299 401782 -3277
rect 401320 -3385 401782 -3299
rect 404410 -3274 404486 -3232
rect 404538 -3274 405126 -3219
rect 407820 -3232 407830 -3219
rect 404410 -3277 405126 -3274
rect 401324 -3393 401524 -3385
rect 401340 -3397 401508 -3393
rect 397922 -3628 397924 -3574
rect 401066 -3600 401240 -3514
rect 401266 -3574 401366 -3450
rect 404410 -3514 404554 -3277
rect 404740 -3299 405126 -3277
rect 404664 -3385 405126 -3299
rect 407754 -3274 407830 -3232
rect 407882 -3274 408470 -3219
rect 411164 -3232 411174 -3219
rect 407754 -3277 408470 -3274
rect 404668 -3393 404868 -3385
rect 404684 -3397 404852 -3393
rect 401266 -3628 401268 -3574
rect 404410 -3600 404584 -3514
rect 404610 -3574 404710 -3450
rect 407754 -3514 407898 -3277
rect 408084 -3299 408470 -3277
rect 408008 -3385 408470 -3299
rect 411098 -3274 411174 -3232
rect 411226 -3274 411814 -3219
rect 414508 -3232 414518 -3219
rect 411098 -3277 411814 -3274
rect 408012 -3393 408212 -3385
rect 408028 -3397 408196 -3393
rect 404610 -3628 404612 -3574
rect 407754 -3600 407928 -3514
rect 407954 -3574 408054 -3450
rect 411098 -3514 411242 -3277
rect 411428 -3299 411814 -3277
rect 411352 -3385 411814 -3299
rect 414442 -3274 414518 -3232
rect 414570 -3274 415158 -3219
rect 417852 -3232 417862 -3219
rect 414442 -3277 415158 -3274
rect 411356 -3393 411556 -3385
rect 411372 -3397 411540 -3393
rect 407954 -3628 407956 -3574
rect 411098 -3600 411272 -3514
rect 411298 -3574 411398 -3450
rect 414442 -3514 414586 -3277
rect 414772 -3299 415158 -3277
rect 414696 -3385 415158 -3299
rect 417786 -3274 417862 -3232
rect 417914 -3274 418502 -3219
rect 421196 -3232 421206 -3219
rect 417786 -3277 418502 -3274
rect 414700 -3393 414900 -3385
rect 414716 -3397 414884 -3393
rect 411298 -3628 411300 -3574
rect 414442 -3600 414616 -3514
rect 414642 -3574 414742 -3450
rect 417786 -3514 417930 -3277
rect 418116 -3299 418502 -3277
rect 418040 -3385 418502 -3299
rect 421130 -3274 421206 -3232
rect 421258 -3274 421846 -3219
rect 424540 -3232 424550 -3219
rect 421130 -3277 421846 -3274
rect 418044 -3393 418244 -3385
rect 418060 -3397 418228 -3393
rect 414642 -3628 414644 -3574
rect 417786 -3600 417960 -3514
rect 417986 -3574 418086 -3450
rect 421130 -3514 421274 -3277
rect 421460 -3299 421846 -3277
rect 421384 -3385 421846 -3299
rect 424474 -3274 424550 -3232
rect 424602 -3274 425190 -3219
rect 427884 -3232 427894 -3219
rect 424474 -3277 425190 -3274
rect 421388 -3393 421588 -3385
rect 421404 -3397 421572 -3393
rect 417986 -3628 417988 -3574
rect 421130 -3600 421304 -3514
rect 421330 -3574 421430 -3450
rect 424474 -3514 424618 -3277
rect 424804 -3299 425190 -3277
rect 424728 -3385 425190 -3299
rect 427818 -3274 427894 -3232
rect 424732 -3393 424932 -3385
rect 424748 -3397 424916 -3393
rect 421330 -3628 421332 -3574
rect 424474 -3600 424648 -3514
rect 424674 -3574 424774 -3450
rect 427818 -3514 427962 -3274
rect 424674 -3628 424676 -3574
rect 427818 -3600 427992 -3514
rect 428018 -3574 428118 -3450
rect 428018 -3628 428020 -3574
rect 3015 -4371 3159 -4324
rect 3196 -4371 3213 -4270
rect 6359 -4371 6503 -4324
rect 6540 -4371 6557 -4270
rect 9703 -4371 9847 -4324
rect 9884 -4371 9901 -4270
rect 13047 -4371 13191 -4324
rect 13228 -4371 13245 -4270
rect 16391 -4371 16535 -4324
rect 16572 -4371 16589 -4270
rect 19735 -4371 19879 -4324
rect 19916 -4371 19933 -4270
rect 23079 -4371 23223 -4324
rect 23260 -4371 23277 -4270
rect 26423 -4371 26567 -4324
rect 26604 -4371 26621 -4270
rect 29767 -4371 29911 -4324
rect 29948 -4371 29965 -4270
rect 33111 -4371 33255 -4324
rect 33292 -4371 33309 -4270
rect 36455 -4371 36599 -4324
rect 36636 -4371 36653 -4270
rect 39799 -4371 39943 -4324
rect 39980 -4371 39997 -4270
rect 43143 -4371 43287 -4324
rect 43324 -4371 43341 -4270
rect 46487 -4371 46631 -4324
rect 46668 -4371 46685 -4270
rect 49831 -4371 49975 -4324
rect 50012 -4371 50029 -4270
rect 53175 -4371 53319 -4324
rect 53356 -4371 53373 -4270
rect 56519 -4371 56663 -4324
rect 56700 -4371 56717 -4270
rect 59863 -4371 60007 -4324
rect 60044 -4371 60061 -4270
rect 63207 -4371 63351 -4324
rect 63388 -4371 63405 -4270
rect 66551 -4371 66695 -4324
rect 66732 -4371 66749 -4270
rect 69895 -4371 70039 -4324
rect 70076 -4371 70093 -4270
rect 73239 -4371 73383 -4324
rect 73420 -4371 73437 -4270
rect 76583 -4371 76727 -4324
rect 76764 -4371 76781 -4270
rect 79927 -4371 80071 -4324
rect 80108 -4371 80125 -4270
rect 83271 -4371 83415 -4324
rect 83452 -4371 83469 -4270
rect 86615 -4371 86759 -4324
rect 86796 -4371 86813 -4270
rect 89959 -4371 90103 -4324
rect 90140 -4371 90157 -4270
rect 93303 -4371 93447 -4324
rect 93484 -4371 93501 -4270
rect 96647 -4371 96791 -4324
rect 96828 -4371 96845 -4270
rect 99991 -4371 100135 -4324
rect 100172 -4371 100189 -4270
rect 103335 -4371 103479 -4324
rect 103516 -4371 103533 -4270
rect 106679 -4371 106823 -4324
rect 106860 -4371 106877 -4270
rect 110023 -4371 110167 -4324
rect 110204 -4371 110221 -4270
rect 113367 -4371 113511 -4324
rect 113548 -4371 113565 -4270
rect 116711 -4371 116855 -4324
rect 116892 -4371 116909 -4270
rect 120055 -4371 120199 -4324
rect 120236 -4371 120253 -4270
rect 123399 -4371 123543 -4324
rect 123580 -4371 123597 -4270
rect 126743 -4371 126887 -4324
rect 126924 -4371 126941 -4270
rect 130087 -4371 130231 -4324
rect 130268 -4371 130285 -4270
rect 133431 -4371 133575 -4324
rect 133612 -4371 133629 -4270
rect 136775 -4371 136919 -4324
rect 136956 -4371 136973 -4270
rect 140119 -4371 140263 -4324
rect 140300 -4371 140317 -4270
rect 143463 -4371 143607 -4324
rect 143644 -4371 143661 -4270
rect 146807 -4371 146951 -4324
rect 146988 -4371 147005 -4270
rect 150151 -4371 150295 -4324
rect 150332 -4371 150349 -4270
rect 153495 -4371 153639 -4324
rect 153676 -4371 153693 -4270
rect 156839 -4371 156983 -4324
rect 157020 -4371 157037 -4270
rect 160183 -4371 160327 -4324
rect 160364 -4371 160381 -4270
rect 163527 -4371 163671 -4324
rect 163708 -4371 163725 -4270
rect 166871 -4371 167015 -4324
rect 167052 -4371 167069 -4270
rect 170215 -4371 170359 -4324
rect 170396 -4371 170413 -4270
rect 173559 -4371 173703 -4324
rect 173740 -4371 173757 -4270
rect 176903 -4371 177047 -4324
rect 177084 -4371 177101 -4270
rect 180247 -4371 180391 -4324
rect 180428 -4371 180445 -4270
rect 183591 -4371 183735 -4324
rect 183772 -4371 183789 -4270
rect 186935 -4371 187079 -4324
rect 187116 -4371 187133 -4270
rect 190279 -4371 190423 -4324
rect 190460 -4371 190477 -4270
rect 193623 -4371 193767 -4324
rect 193804 -4371 193821 -4270
rect 196967 -4371 197111 -4324
rect 197148 -4371 197165 -4270
rect 200311 -4371 200455 -4324
rect 200492 -4371 200509 -4270
rect 203655 -4371 203799 -4324
rect 203836 -4371 203853 -4270
rect 206999 -4371 207143 -4324
rect 207180 -4371 207197 -4270
rect 210343 -4371 210487 -4324
rect 210524 -4371 210541 -4270
rect 217031 -4371 217175 -4324
rect 217212 -4371 217229 -4270
rect 220375 -4371 220519 -4324
rect 220556 -4371 220573 -4270
rect 223719 -4371 223863 -4324
rect 223900 -4371 223917 -4270
rect 227063 -4371 227207 -4324
rect 227244 -4371 227261 -4270
rect 230407 -4371 230551 -4324
rect 230588 -4371 230605 -4270
rect 233751 -4371 233895 -4324
rect 233932 -4371 233949 -4270
rect 237095 -4371 237239 -4324
rect 237276 -4371 237293 -4270
rect 240439 -4371 240583 -4324
rect 240620 -4371 240637 -4270
rect 243783 -4371 243927 -4324
rect 243964 -4371 243981 -4270
rect 247127 -4371 247271 -4324
rect 247308 -4371 247325 -4270
rect 250471 -4371 250615 -4324
rect 250652 -4371 250669 -4270
rect 253815 -4371 253959 -4324
rect 253996 -4371 254013 -4270
rect 257159 -4371 257303 -4324
rect 257340 -4371 257357 -4270
rect 260503 -4371 260647 -4324
rect 260684 -4371 260701 -4270
rect 263847 -4371 263991 -4324
rect 264028 -4371 264045 -4270
rect 267191 -4371 267335 -4324
rect 267372 -4371 267389 -4270
rect 270535 -4371 270679 -4324
rect 270716 -4371 270733 -4270
rect 273879 -4371 274023 -4324
rect 274060 -4371 274077 -4270
rect 277223 -4371 277367 -4324
rect 277404 -4371 277421 -4270
rect 280567 -4371 280711 -4324
rect 280748 -4371 280765 -4270
rect 283911 -4371 284055 -4324
rect 284092 -4371 284109 -4270
rect 287255 -4371 287399 -4324
rect 287436 -4371 287453 -4270
rect 290599 -4371 290743 -4324
rect 290780 -4371 290797 -4270
rect 293943 -4371 294087 -4324
rect 294124 -4371 294141 -4270
rect 297287 -4371 297431 -4324
rect 297468 -4371 297485 -4270
rect 300631 -4371 300775 -4324
rect 300812 -4371 300829 -4270
rect 303975 -4371 304119 -4324
rect 304156 -4371 304173 -4270
rect 307319 -4371 307463 -4324
rect 307500 -4371 307517 -4270
rect 310663 -4371 310807 -4324
rect 310844 -4371 310861 -4270
rect 314007 -4371 314151 -4324
rect 314188 -4371 314205 -4270
rect 317351 -4371 317495 -4324
rect 317532 -4371 317549 -4270
rect 320695 -4371 320839 -4324
rect 320876 -4371 320893 -4270
rect 324039 -4371 324183 -4324
rect 324220 -4371 324237 -4270
rect 327383 -4371 327527 -4324
rect 327564 -4371 327581 -4270
rect 330727 -4371 330871 -4324
rect 330908 -4371 330925 -4270
rect 334071 -4371 334215 -4324
rect 334252 -4371 334269 -4270
rect 337415 -4371 337559 -4324
rect 337596 -4371 337613 -4270
rect 340759 -4371 340903 -4324
rect 340940 -4371 340957 -4270
rect 344103 -4371 344247 -4324
rect 344284 -4371 344301 -4270
rect 347447 -4371 347591 -4324
rect 347628 -4371 347645 -4270
rect 350791 -4371 350935 -4324
rect 350972 -4371 350989 -4270
rect 354135 -4371 354279 -4324
rect 354316 -4371 354333 -4270
rect 357479 -4371 357623 -4324
rect 357660 -4371 357677 -4270
rect 360823 -4371 360967 -4324
rect 361004 -4371 361021 -4270
rect 364167 -4371 364311 -4324
rect 364348 -4371 364365 -4270
rect 367511 -4371 367655 -4324
rect 367692 -4371 367709 -4270
rect 370855 -4371 370999 -4324
rect 371036 -4371 371053 -4270
rect 374199 -4371 374343 -4324
rect 374380 -4371 374397 -4270
rect 377543 -4371 377687 -4324
rect 377724 -4371 377741 -4270
rect 380887 -4371 381031 -4324
rect 381068 -4371 381085 -4270
rect 384231 -4371 384375 -4324
rect 384412 -4371 384429 -4270
rect 387575 -4371 387719 -4324
rect 387756 -4371 387773 -4270
rect 390919 -4371 391063 -4324
rect 391100 -4371 391117 -4270
rect 394263 -4371 394407 -4324
rect 394444 -4371 394461 -4270
rect 397607 -4371 397751 -4324
rect 397788 -4371 397805 -4270
rect 400951 -4371 401095 -4324
rect 401132 -4371 401149 -4270
rect 404295 -4371 404439 -4324
rect 404476 -4371 404493 -4270
rect 407639 -4371 407783 -4324
rect 407820 -4371 407837 -4270
rect 410983 -4371 411127 -4324
rect 411164 -4371 411181 -4270
rect 414327 -4371 414471 -4324
rect 414508 -4371 414525 -4270
rect 417671 -4371 417815 -4324
rect 417852 -4371 417869 -4270
rect 421015 -4371 421159 -4324
rect 421196 -4371 421213 -4270
rect 424359 -4371 424503 -4324
rect 424540 -4371 424557 -4270
rect 427703 -4371 427847 -4324
rect 427884 -4371 427901 -4270
rect 3015 -4382 3787 -4371
rect 6359 -4382 7131 -4371
rect 9703 -4382 10475 -4371
rect 13047 -4382 13819 -4371
rect 16391 -4382 17163 -4371
rect 19735 -4382 20507 -4371
rect 23079 -4382 23851 -4371
rect 26423 -4382 27195 -4371
rect 29767 -4382 30539 -4371
rect 33111 -4382 33883 -4371
rect 36455 -4382 37227 -4371
rect 39799 -4382 40571 -4371
rect 43143 -4382 43915 -4371
rect 46487 -4382 47259 -4371
rect 49831 -4382 50603 -4371
rect 53175 -4382 53947 -4371
rect 56519 -4382 57291 -4371
rect 59863 -4382 60635 -4371
rect 63207 -4382 63979 -4371
rect 66551 -4382 67323 -4371
rect 69895 -4382 70667 -4371
rect 73239 -4382 74011 -4371
rect 76583 -4382 77355 -4371
rect 79927 -4382 80699 -4371
rect 83271 -4382 84043 -4371
rect 86615 -4382 87387 -4371
rect 89959 -4382 90731 -4371
rect 93303 -4382 94075 -4371
rect 96647 -4382 97419 -4371
rect 99991 -4382 100763 -4371
rect 103335 -4382 104107 -4371
rect 106679 -4382 107451 -4371
rect 110023 -4382 110795 -4371
rect 113367 -4382 114139 -4371
rect 116711 -4382 117483 -4371
rect 120055 -4382 120827 -4371
rect 123399 -4382 124171 -4371
rect 126743 -4382 127515 -4371
rect 130087 -4382 130859 -4371
rect 133431 -4382 134203 -4371
rect 136775 -4382 137547 -4371
rect 140119 -4382 140891 -4371
rect 143463 -4382 144235 -4371
rect 146807 -4382 147579 -4371
rect 150151 -4382 150923 -4371
rect 153495 -4382 154267 -4371
rect 156839 -4382 157611 -4371
rect 160183 -4382 160955 -4371
rect 163527 -4382 164299 -4371
rect 166871 -4382 167643 -4371
rect 170215 -4382 170987 -4371
rect 173559 -4382 174331 -4371
rect 176903 -4382 177675 -4371
rect 180247 -4382 181019 -4371
rect 183591 -4382 184363 -4371
rect 186935 -4382 187707 -4371
rect 190279 -4382 191051 -4371
rect 193623 -4382 194395 -4371
rect 196967 -4382 197739 -4371
rect 200311 -4382 201083 -4371
rect 203655 -4382 204427 -4371
rect 206999 -4382 207771 -4371
rect 210343 -4382 211115 -4371
rect 217031 -4382 217147 -4371
rect 3101 -4407 3787 -4382
rect 6445 -4407 7131 -4382
rect 9789 -4407 10475 -4382
rect 13133 -4407 13819 -4382
rect 16477 -4407 17163 -4382
rect 19821 -4407 20507 -4382
rect 23165 -4407 23851 -4382
rect 26509 -4407 27195 -4382
rect 29853 -4407 30539 -4382
rect 33197 -4407 33883 -4382
rect 36541 -4407 37227 -4382
rect 39885 -4407 40571 -4382
rect 43229 -4407 43915 -4382
rect 46573 -4407 47259 -4382
rect 49917 -4407 50603 -4382
rect 53261 -4407 53947 -4382
rect 56605 -4407 57291 -4382
rect 59949 -4407 60635 -4382
rect 63293 -4407 63979 -4382
rect 66637 -4407 67323 -4382
rect 69981 -4407 70667 -4382
rect 73325 -4407 74011 -4382
rect 76669 -4407 77355 -4382
rect 80013 -4407 80699 -4382
rect 83357 -4407 84043 -4382
rect 86701 -4407 87387 -4382
rect 90045 -4407 90731 -4382
rect 93389 -4407 94075 -4382
rect 96733 -4407 97419 -4382
rect 100077 -4407 100763 -4382
rect 103421 -4407 104107 -4382
rect 106765 -4407 107451 -4382
rect 110109 -4407 110795 -4382
rect 113453 -4407 114139 -4382
rect 116797 -4407 117483 -4382
rect 120141 -4407 120827 -4382
rect 123485 -4407 124171 -4382
rect 126829 -4407 127515 -4382
rect 130173 -4407 130859 -4382
rect 133517 -4407 134203 -4382
rect 136861 -4407 137547 -4382
rect 140205 -4407 140891 -4382
rect 143549 -4407 144235 -4382
rect 146893 -4407 147579 -4382
rect 150237 -4407 150923 -4382
rect 153581 -4407 154267 -4382
rect 156925 -4407 157611 -4382
rect 160269 -4407 160955 -4382
rect 163613 -4407 164299 -4382
rect 166957 -4407 167643 -4382
rect 170301 -4407 170987 -4382
rect 173645 -4407 174331 -4382
rect 176989 -4407 177675 -4382
rect 180333 -4407 181019 -4382
rect 183677 -4407 184363 -4382
rect 187021 -4407 187707 -4382
rect 190365 -4407 191051 -4382
rect 193709 -4407 194395 -4382
rect 197053 -4407 197739 -4382
rect 200397 -4407 201083 -4382
rect 203741 -4407 204427 -4382
rect 207085 -4407 207771 -4382
rect 210429 -4407 211115 -4382
rect 217117 -4407 217147 -4382
rect 3113 -4436 3787 -4407
rect 6457 -4436 7131 -4407
rect 9801 -4436 10475 -4407
rect 13145 -4436 13819 -4407
rect 16489 -4436 17163 -4407
rect 19833 -4436 20507 -4407
rect 23177 -4436 23851 -4407
rect 26521 -4436 27195 -4407
rect 29865 -4436 30539 -4407
rect 33209 -4436 33883 -4407
rect 36553 -4436 37227 -4407
rect 39897 -4436 40571 -4407
rect 43241 -4436 43915 -4407
rect 46585 -4436 47259 -4407
rect 49929 -4436 50603 -4407
rect 53273 -4436 53947 -4407
rect 56617 -4436 57291 -4407
rect 59961 -4436 60635 -4407
rect 63305 -4436 63979 -4407
rect 66649 -4436 67323 -4407
rect 69993 -4436 70667 -4407
rect 73337 -4436 74011 -4407
rect 76681 -4436 77355 -4407
rect 80025 -4436 80699 -4407
rect 83369 -4436 84043 -4407
rect 86713 -4436 87387 -4407
rect 90057 -4436 90731 -4407
rect 93401 -4436 94075 -4407
rect 96745 -4436 97419 -4407
rect 100089 -4436 100763 -4407
rect 103433 -4436 104107 -4407
rect 106777 -4436 107451 -4407
rect 110121 -4436 110795 -4407
rect 113465 -4436 114139 -4407
rect 116809 -4436 117483 -4407
rect 120153 -4436 120827 -4407
rect 123497 -4436 124171 -4407
rect 126841 -4436 127515 -4407
rect 130185 -4436 130859 -4407
rect 133529 -4436 134203 -4407
rect 136873 -4436 137547 -4407
rect 140217 -4436 140891 -4407
rect 143561 -4436 144235 -4407
rect 146905 -4436 147579 -4407
rect 150249 -4436 150923 -4407
rect 153593 -4436 154267 -4407
rect 156937 -4436 157611 -4407
rect 160281 -4436 160955 -4407
rect 163625 -4436 164299 -4407
rect 166969 -4436 167643 -4407
rect 170313 -4436 170987 -4407
rect 173657 -4436 174331 -4407
rect 177001 -4436 177675 -4407
rect 180345 -4436 181019 -4407
rect 183689 -4436 184363 -4407
rect 187033 -4436 187707 -4407
rect 190377 -4436 191051 -4407
rect 193721 -4436 194395 -4407
rect 197065 -4436 197739 -4407
rect 200409 -4436 201083 -4407
rect 203753 -4436 204427 -4407
rect 207097 -4436 207771 -4407
rect 210441 -4436 211115 -4407
rect 3113 -4848 3846 -4436
rect 4295 -4848 4342 -4483
rect 4349 -4848 4396 -4537
rect 6457 -4848 7190 -4436
rect 7639 -4848 7686 -4483
rect 7693 -4848 7740 -4537
rect 9801 -4848 10534 -4436
rect 10983 -4848 11030 -4483
rect 11037 -4848 11084 -4537
rect 13145 -4848 13878 -4436
rect 14327 -4848 14374 -4483
rect 14381 -4848 14428 -4537
rect 16489 -4848 17222 -4436
rect 17671 -4848 17718 -4483
rect 17725 -4848 17772 -4537
rect 19833 -4848 20566 -4436
rect 21015 -4848 21062 -4483
rect 21069 -4848 21116 -4537
rect 23177 -4848 23910 -4436
rect 24359 -4848 24406 -4483
rect 24413 -4848 24460 -4537
rect 26521 -4848 27254 -4436
rect 27703 -4848 27750 -4483
rect 27757 -4848 27804 -4537
rect 29865 -4848 30598 -4436
rect 31047 -4848 31094 -4483
rect 31101 -4848 31148 -4537
rect 33209 -4848 33942 -4436
rect 34391 -4848 34438 -4483
rect 34445 -4848 34492 -4537
rect 36553 -4848 37286 -4436
rect 37735 -4848 37782 -4483
rect 37789 -4848 37836 -4537
rect 39897 -4848 40630 -4436
rect 41079 -4848 41126 -4483
rect 41133 -4848 41180 -4537
rect 43241 -4848 43974 -4436
rect 44423 -4848 44470 -4483
rect 44477 -4848 44524 -4537
rect 46585 -4848 47318 -4436
rect 47767 -4848 47814 -4483
rect 47821 -4848 47868 -4537
rect 49929 -4848 50662 -4436
rect 51111 -4848 51158 -4483
rect 51165 -4848 51212 -4537
rect 53273 -4848 54006 -4436
rect 54455 -4848 54502 -4483
rect 54509 -4848 54556 -4537
rect 56617 -4848 57350 -4436
rect 57799 -4848 57846 -4483
rect 57853 -4848 57900 -4537
rect 59961 -4848 60694 -4436
rect 61143 -4848 61190 -4483
rect 61197 -4848 61244 -4537
rect 63305 -4848 64038 -4436
rect 64487 -4848 64534 -4483
rect 64541 -4848 64588 -4537
rect 66649 -4848 67382 -4436
rect 67831 -4848 67878 -4483
rect 67885 -4848 67932 -4537
rect 69993 -4848 70726 -4436
rect 71175 -4848 71222 -4483
rect 71229 -4848 71276 -4537
rect 73337 -4848 74070 -4436
rect 74519 -4848 74566 -4483
rect 74573 -4848 74620 -4537
rect 76681 -4848 77414 -4436
rect 77863 -4848 77910 -4483
rect 77917 -4848 77964 -4537
rect 80025 -4848 80758 -4436
rect 81207 -4848 81254 -4483
rect 81261 -4848 81308 -4537
rect 83369 -4848 84102 -4436
rect 84551 -4848 84598 -4483
rect 84605 -4848 84652 -4537
rect 86713 -4848 87446 -4436
rect 87895 -4848 87942 -4483
rect 87949 -4848 87996 -4537
rect 90057 -4848 90790 -4436
rect 91239 -4848 91286 -4483
rect 91293 -4848 91340 -4537
rect 93401 -4848 94134 -4436
rect 94583 -4848 94630 -4483
rect 94637 -4848 94684 -4537
rect 96745 -4848 97478 -4436
rect 97927 -4848 97974 -4483
rect 97981 -4848 98028 -4537
rect 100089 -4848 100822 -4436
rect 101271 -4848 101318 -4483
rect 101325 -4848 101372 -4537
rect 103433 -4848 104166 -4436
rect 104615 -4848 104662 -4483
rect 104669 -4848 104716 -4537
rect 106777 -4848 107510 -4436
rect 107959 -4848 108006 -4483
rect 108013 -4848 108060 -4537
rect 110121 -4848 110854 -4436
rect 111303 -4848 111350 -4483
rect 111357 -4848 111404 -4537
rect 113465 -4848 114198 -4436
rect 114647 -4848 114694 -4483
rect 114701 -4848 114748 -4537
rect 116809 -4848 117542 -4436
rect 117991 -4848 118038 -4483
rect 118045 -4848 118092 -4537
rect 120153 -4848 120886 -4436
rect 121335 -4848 121382 -4483
rect 121389 -4848 121436 -4537
rect 123497 -4848 124230 -4436
rect 124679 -4848 124726 -4483
rect 124733 -4848 124780 -4537
rect 126841 -4848 127574 -4436
rect 128023 -4848 128070 -4483
rect 128077 -4848 128124 -4537
rect 130185 -4848 130918 -4436
rect 131367 -4848 131414 -4483
rect 131421 -4848 131468 -4537
rect 133529 -4848 134262 -4436
rect 134711 -4848 134758 -4483
rect 134765 -4848 134812 -4537
rect 136873 -4848 137606 -4436
rect 138055 -4848 138102 -4483
rect 138109 -4848 138156 -4537
rect 140217 -4848 140950 -4436
rect 141399 -4848 141446 -4483
rect 141453 -4848 141500 -4537
rect 143561 -4848 144294 -4436
rect 144743 -4848 144790 -4483
rect 144797 -4848 144844 -4537
rect 146905 -4848 147638 -4436
rect 148087 -4848 148134 -4483
rect 148141 -4848 148188 -4537
rect 150249 -4848 150982 -4436
rect 151431 -4848 151478 -4483
rect 151485 -4848 151532 -4537
rect 153593 -4848 154326 -4436
rect 154775 -4848 154822 -4483
rect 154829 -4848 154876 -4537
rect 156937 -4848 157670 -4436
rect 158119 -4848 158166 -4483
rect 158173 -4848 158220 -4537
rect 160281 -4848 161014 -4436
rect 161463 -4848 161510 -4483
rect 161517 -4848 161564 -4537
rect 163625 -4848 164358 -4436
rect 164807 -4848 164854 -4483
rect 164861 -4848 164908 -4537
rect 166969 -4848 167702 -4436
rect 168151 -4848 168198 -4483
rect 168205 -4848 168252 -4537
rect 170313 -4848 171046 -4436
rect 171495 -4848 171542 -4483
rect 171549 -4848 171596 -4537
rect 173657 -4848 174390 -4436
rect 174839 -4848 174886 -4483
rect 174893 -4848 174940 -4537
rect 177001 -4848 177734 -4436
rect 178183 -4848 178230 -4483
rect 178237 -4848 178284 -4537
rect 180345 -4848 181078 -4436
rect 181527 -4848 181574 -4483
rect 181581 -4848 181628 -4537
rect 183689 -4848 184422 -4436
rect 184871 -4848 184918 -4483
rect 184925 -4848 184972 -4537
rect 187033 -4848 187766 -4436
rect 188215 -4848 188262 -4483
rect 188269 -4848 188316 -4537
rect 190377 -4848 191110 -4436
rect 191559 -4848 191606 -4483
rect 191613 -4848 191660 -4537
rect 193721 -4848 194454 -4436
rect 194903 -4848 194950 -4483
rect 194957 -4848 195004 -4537
rect 197065 -4848 197798 -4436
rect 198247 -4848 198294 -4483
rect 198301 -4848 198348 -4537
rect 200409 -4848 201142 -4436
rect 201591 -4848 201638 -4483
rect 201645 -4848 201692 -4537
rect 203753 -4848 204486 -4436
rect 204935 -4848 204982 -4483
rect 204989 -4848 205036 -4537
rect 207097 -4848 207830 -4436
rect 208279 -4848 208326 -4483
rect 208333 -4848 208380 -4537
rect 210441 -4848 211174 -4436
rect 211623 -4848 211670 -4483
rect 211677 -4848 211724 -4537
rect 3113 -4906 4467 -4848
rect 6457 -4906 7811 -4848
rect 9801 -4906 11155 -4848
rect 13145 -4906 14499 -4848
rect 16489 -4906 17843 -4848
rect 19833 -4906 21187 -4848
rect 23177 -4906 24531 -4848
rect 26521 -4906 27875 -4848
rect 29865 -4906 31219 -4848
rect 33209 -4906 34563 -4848
rect 36553 -4906 37907 -4848
rect 39897 -4906 41251 -4848
rect 43241 -4906 44595 -4848
rect 46585 -4906 47939 -4848
rect 49929 -4906 51283 -4848
rect 53273 -4906 54627 -4848
rect 56617 -4906 57971 -4848
rect 59961 -4906 61315 -4848
rect 63305 -4906 64659 -4848
rect 66649 -4906 68003 -4848
rect 69993 -4906 71347 -4848
rect 73337 -4906 74691 -4848
rect 76681 -4906 78035 -4848
rect 80025 -4906 81379 -4848
rect 83369 -4906 84723 -4848
rect 86713 -4906 88067 -4848
rect 90057 -4906 91411 -4848
rect 93401 -4906 94755 -4848
rect 96745 -4906 98099 -4848
rect 100089 -4906 101443 -4848
rect 103433 -4906 104787 -4848
rect 106777 -4906 108131 -4848
rect 110121 -4906 111475 -4848
rect 113465 -4906 114819 -4848
rect 116809 -4906 118163 -4848
rect 120153 -4906 121507 -4848
rect 123497 -4906 124851 -4848
rect 126841 -4906 128195 -4848
rect 130185 -4906 131539 -4848
rect 133529 -4906 134883 -4848
rect 136873 -4906 138227 -4848
rect 140217 -4906 141571 -4848
rect 143561 -4906 144915 -4848
rect 146905 -4906 148259 -4848
rect 150249 -4906 151603 -4848
rect 153593 -4906 154947 -4848
rect 156937 -4906 158291 -4848
rect 160281 -4906 161635 -4848
rect 163625 -4906 164979 -4848
rect 166969 -4906 168323 -4848
rect 170313 -4906 171667 -4848
rect 173657 -4906 175011 -4848
rect 177001 -4906 178355 -4848
rect 180345 -4906 181699 -4848
rect 183689 -4906 185043 -4848
rect 187033 -4906 188387 -4848
rect 190377 -4906 191731 -4848
rect 193721 -4906 195075 -4848
rect 197065 -4906 198419 -4848
rect 200409 -4906 201763 -4848
rect 203753 -4906 205107 -4848
rect 207097 -4906 208451 -4848
rect 210441 -4906 211496 -4848
rect 2720 -4943 4467 -4906
rect 5884 -4943 7811 -4906
rect 9228 -4943 11155 -4906
rect 12572 -4943 14499 -4906
rect 15916 -4943 17843 -4906
rect 19260 -4943 21187 -4906
rect 22604 -4943 24531 -4906
rect 25948 -4943 27875 -4906
rect 29292 -4943 31219 -4906
rect 32636 -4943 34563 -4906
rect 35980 -4943 37907 -4906
rect 39324 -4943 41251 -4906
rect 42668 -4943 44595 -4906
rect 46012 -4943 47939 -4906
rect 49356 -4943 51283 -4906
rect 52700 -4943 54627 -4906
rect 56044 -4943 57971 -4906
rect 59388 -4943 61315 -4906
rect 62732 -4943 64659 -4906
rect 66076 -4943 68003 -4906
rect 69420 -4943 71347 -4906
rect 72764 -4943 74691 -4906
rect 76108 -4943 78035 -4906
rect 79452 -4943 81379 -4906
rect 82796 -4943 84723 -4906
rect 86140 -4943 88067 -4906
rect 89484 -4943 91411 -4906
rect 92828 -4943 94755 -4906
rect 96172 -4943 98099 -4906
rect 99516 -4943 101443 -4906
rect 102860 -4943 104787 -4906
rect 106204 -4943 108131 -4906
rect 109548 -4943 111475 -4906
rect 112892 -4943 114819 -4906
rect 116236 -4943 118163 -4906
rect 119580 -4943 121507 -4906
rect 122924 -4943 124851 -4906
rect 126268 -4943 128195 -4906
rect 129612 -4943 131539 -4906
rect 132956 -4943 134883 -4906
rect 136300 -4943 138227 -4906
rect 139644 -4943 141571 -4906
rect 142988 -4943 144915 -4906
rect 146332 -4943 148259 -4906
rect 149676 -4943 151603 -4906
rect 153020 -4943 154947 -4906
rect 156364 -4943 158291 -4906
rect 159708 -4943 161635 -4906
rect 163052 -4943 164979 -4906
rect 166396 -4943 168323 -4906
rect 169740 -4943 171667 -4906
rect 173084 -4943 175011 -4906
rect 176428 -4943 178355 -4906
rect 179772 -4943 181699 -4906
rect 183116 -4943 185043 -4906
rect 186460 -4943 188387 -4906
rect 189804 -4943 191731 -4906
rect 193148 -4943 195075 -4906
rect 196492 -4943 198419 -4906
rect 199836 -4943 201763 -4906
rect 203180 -4943 205107 -4906
rect 206524 -4943 208451 -4906
rect 2720 -5067 4969 -4943
rect 5884 -5067 8313 -4943
rect 9228 -5067 11657 -4943
rect 12572 -5067 15001 -4943
rect 15916 -5067 18345 -4943
rect 19260 -5067 21689 -4943
rect 22604 -5067 25033 -4943
rect 25948 -5067 28377 -4943
rect 29292 -5067 31721 -4943
rect 32636 -5067 35065 -4943
rect 35980 -5067 38409 -4943
rect 39324 -5067 41753 -4943
rect 42668 -5067 45097 -4943
rect 46012 -5067 48441 -4943
rect 49356 -5067 51785 -4943
rect 52700 -5067 55129 -4943
rect 56044 -5067 58473 -4943
rect 59388 -5067 61817 -4943
rect 62732 -5067 65161 -4943
rect 66076 -5067 68505 -4943
rect 69420 -5067 71849 -4943
rect 72764 -5067 75193 -4943
rect 76108 -5067 78537 -4943
rect 79452 -5067 81881 -4943
rect 82796 -5067 85225 -4943
rect 86140 -5067 88569 -4943
rect 89484 -5067 91913 -4943
rect 92828 -5067 95257 -4943
rect 96172 -5067 98601 -4943
rect 99516 -5067 101945 -4943
rect 102860 -5067 105289 -4943
rect 106204 -5067 108633 -4943
rect 109548 -5067 111977 -4943
rect 112892 -5067 115321 -4943
rect 116236 -5067 118665 -4943
rect 119580 -5067 122009 -4943
rect 122924 -5067 125353 -4943
rect 126268 -5067 128697 -4943
rect 129612 -5067 132041 -4943
rect 132956 -5067 135385 -4943
rect 136300 -5067 138729 -4943
rect 139644 -5067 142073 -4943
rect 142988 -5067 145417 -4943
rect 146332 -5067 148761 -4943
rect 149676 -5067 152105 -4943
rect 153020 -5067 155449 -4943
rect 156364 -5067 158793 -4943
rect 159708 -5067 162137 -4943
rect 163052 -5067 165481 -4943
rect 166396 -5067 168825 -4943
rect 169740 -5067 172169 -4943
rect 173084 -5067 175513 -4943
rect 176428 -5067 178857 -4943
rect 179772 -5067 182201 -4943
rect 183116 -5067 185545 -4943
rect 186460 -5067 188889 -4943
rect 189804 -5067 192233 -4943
rect 193148 -5067 195577 -4943
rect 196492 -5067 198921 -4943
rect 199836 -5067 202265 -4943
rect 203180 -5067 205609 -4943
rect 206524 -5067 208953 -4943
rect 2720 -6022 5022 -5067
rect 5884 -6022 8366 -5067
rect 9228 -6022 11710 -5067
rect 12572 -6022 15054 -5067
rect 15916 -6022 18398 -5067
rect 19260 -6022 21742 -5067
rect 22604 -6022 25086 -5067
rect 25948 -6022 28430 -5067
rect 29292 -6022 31774 -5067
rect 32636 -6022 35118 -5067
rect 35980 -6022 38462 -5067
rect 39324 -6022 41806 -5067
rect 42668 -6022 45150 -5067
rect 46012 -6022 48494 -5067
rect 49356 -6022 51838 -5067
rect 52700 -6022 55182 -5067
rect 56044 -6022 58526 -5067
rect 59388 -6022 61870 -5067
rect 62732 -6022 65214 -5067
rect 66076 -6022 68558 -5067
rect 69420 -6022 71902 -5067
rect 72764 -6022 75246 -5067
rect 76108 -6022 78590 -5067
rect 79452 -6022 81934 -5067
rect 82796 -6022 85278 -5067
rect 86140 -6022 88622 -5067
rect 89484 -6022 91966 -5067
rect 92828 -6022 95310 -5067
rect 96172 -6022 98654 -5067
rect 99516 -6022 101998 -5067
rect 102860 -6022 105342 -5067
rect 106204 -6022 108686 -5067
rect 109548 -6022 112030 -5067
rect 112892 -6022 115374 -5067
rect 116236 -6022 118718 -5067
rect 119580 -6022 122062 -5067
rect 122924 -6022 125406 -5067
rect 126268 -6022 128750 -5067
rect 129612 -6022 132094 -5067
rect 132956 -6022 135438 -5067
rect 136300 -6022 138782 -5067
rect 139644 -6022 142126 -5067
rect 142988 -6022 145470 -5067
rect 146332 -6022 148814 -5067
rect 149676 -6022 152158 -5067
rect 153020 -6022 155502 -5067
rect 156364 -6022 158846 -5067
rect 159708 -6022 162190 -5067
rect 163052 -6022 165534 -5067
rect 166396 -6022 168878 -5067
rect 169740 -6022 172222 -5067
rect 173084 -6022 175566 -5067
rect 176428 -6022 178910 -5067
rect 179772 -6022 182254 -5067
rect 183116 -6022 185598 -5067
rect 186460 -6022 188942 -5067
rect 189804 -6022 192286 -5067
rect 193148 -6022 195630 -5067
rect 196492 -6022 198974 -5067
rect 199836 -6022 202318 -5067
rect 203180 -6022 205662 -5067
rect 206524 -6022 209006 -5067
rect 209868 -6022 211496 -4906
rect 217129 -4906 217147 -4407
rect 220375 -4382 221147 -4371
rect 223719 -4382 224491 -4371
rect 227063 -4382 227835 -4371
rect 230407 -4382 231179 -4371
rect 233751 -4382 234523 -4371
rect 237095 -4382 237867 -4371
rect 240439 -4382 241211 -4371
rect 243783 -4382 244555 -4371
rect 247127 -4382 247899 -4371
rect 250471 -4382 251243 -4371
rect 253815 -4382 254587 -4371
rect 257159 -4382 257931 -4371
rect 260503 -4382 261275 -4371
rect 263847 -4382 264619 -4371
rect 267191 -4382 267963 -4371
rect 270535 -4382 271307 -4371
rect 273879 -4382 274651 -4371
rect 277223 -4382 277995 -4371
rect 280567 -4382 281339 -4371
rect 283911 -4382 284683 -4371
rect 287255 -4382 288027 -4371
rect 290599 -4382 291371 -4371
rect 293943 -4382 294715 -4371
rect 297287 -4382 298059 -4371
rect 300631 -4382 301403 -4371
rect 303975 -4382 304747 -4371
rect 307319 -4382 308091 -4371
rect 310663 -4382 311435 -4371
rect 314007 -4382 314779 -4371
rect 317351 -4382 318123 -4371
rect 320695 -4382 321467 -4371
rect 324039 -4382 324811 -4371
rect 327383 -4382 328155 -4371
rect 330727 -4382 331499 -4371
rect 334071 -4382 334843 -4371
rect 337415 -4382 338187 -4371
rect 340759 -4382 341531 -4371
rect 344103 -4382 344875 -4371
rect 347447 -4382 348219 -4371
rect 350791 -4382 351563 -4371
rect 354135 -4382 354907 -4371
rect 357479 -4382 358251 -4371
rect 360823 -4382 361595 -4371
rect 364167 -4382 364939 -4371
rect 367511 -4382 368283 -4371
rect 370855 -4382 371627 -4371
rect 374199 -4382 374971 -4371
rect 377543 -4382 378315 -4371
rect 380887 -4382 381659 -4371
rect 384231 -4382 385003 -4371
rect 387575 -4382 388347 -4371
rect 390919 -4382 391691 -4371
rect 394263 -4382 395035 -4371
rect 397607 -4382 398379 -4371
rect 400951 -4382 401723 -4371
rect 404295 -4382 405067 -4371
rect 407639 -4382 408411 -4371
rect 410983 -4382 411755 -4371
rect 414327 -4382 415099 -4371
rect 417671 -4382 418443 -4371
rect 421015 -4382 421787 -4371
rect 424359 -4382 425131 -4371
rect 427703 -4382 428475 -4371
rect 220461 -4407 221147 -4382
rect 223805 -4407 224491 -4382
rect 227149 -4407 227835 -4382
rect 230493 -4407 231179 -4382
rect 233837 -4407 234523 -4382
rect 237181 -4407 237867 -4382
rect 240525 -4407 241211 -4382
rect 243869 -4407 244555 -4382
rect 247213 -4407 247899 -4382
rect 250557 -4407 251243 -4382
rect 253901 -4407 254587 -4382
rect 257245 -4407 257931 -4382
rect 260589 -4407 261275 -4382
rect 263933 -4407 264619 -4382
rect 267277 -4407 267963 -4382
rect 270621 -4407 271307 -4382
rect 273965 -4407 274651 -4382
rect 277309 -4407 277995 -4382
rect 280653 -4407 281339 -4382
rect 283997 -4407 284683 -4382
rect 287341 -4407 288027 -4382
rect 290685 -4407 291371 -4382
rect 294029 -4407 294715 -4382
rect 297373 -4407 298059 -4382
rect 300717 -4407 301403 -4382
rect 304061 -4407 304747 -4382
rect 307405 -4407 308091 -4382
rect 310749 -4407 311435 -4382
rect 314093 -4407 314779 -4382
rect 317437 -4407 318123 -4382
rect 320781 -4407 321467 -4382
rect 324125 -4407 324811 -4382
rect 327469 -4407 328155 -4382
rect 330813 -4407 331499 -4382
rect 334157 -4407 334843 -4382
rect 337501 -4407 338187 -4382
rect 340845 -4407 341531 -4382
rect 344189 -4407 344875 -4382
rect 347533 -4407 348219 -4382
rect 350877 -4407 351563 -4382
rect 354221 -4407 354907 -4382
rect 357565 -4407 358251 -4382
rect 360909 -4407 361595 -4382
rect 364253 -4407 364939 -4382
rect 367597 -4407 368283 -4382
rect 370941 -4407 371627 -4382
rect 374285 -4407 374971 -4382
rect 377629 -4407 378315 -4382
rect 380973 -4407 381659 -4382
rect 384317 -4407 385003 -4382
rect 387661 -4407 388347 -4382
rect 391005 -4407 391691 -4382
rect 394349 -4407 395035 -4382
rect 397693 -4407 398379 -4382
rect 401037 -4407 401723 -4382
rect 404381 -4407 405067 -4382
rect 407725 -4407 408411 -4382
rect 411069 -4407 411755 -4382
rect 414413 -4407 415099 -4382
rect 417757 -4407 418443 -4382
rect 421101 -4407 421787 -4382
rect 424445 -4407 425131 -4382
rect 427789 -4407 428475 -4382
rect 220473 -4436 221147 -4407
rect 223817 -4436 224491 -4407
rect 227161 -4436 227835 -4407
rect 230505 -4436 231179 -4407
rect 233849 -4436 234523 -4407
rect 237193 -4436 237867 -4407
rect 240537 -4436 241211 -4407
rect 243881 -4436 244555 -4407
rect 247225 -4436 247899 -4407
rect 250569 -4436 251243 -4407
rect 253913 -4436 254587 -4407
rect 257257 -4436 257931 -4407
rect 260601 -4436 261275 -4407
rect 263945 -4436 264619 -4407
rect 267289 -4436 267963 -4407
rect 270633 -4436 271307 -4407
rect 273977 -4436 274651 -4407
rect 277321 -4436 277995 -4407
rect 280665 -4436 281339 -4407
rect 284009 -4436 284683 -4407
rect 287353 -4436 288027 -4407
rect 290697 -4436 291371 -4407
rect 294041 -4436 294715 -4407
rect 297385 -4436 298059 -4407
rect 300729 -4436 301403 -4407
rect 304073 -4436 304747 -4407
rect 307417 -4436 308091 -4407
rect 310761 -4436 311435 -4407
rect 314105 -4436 314779 -4407
rect 317449 -4436 318123 -4407
rect 320793 -4436 321467 -4407
rect 324137 -4436 324811 -4407
rect 327481 -4436 328155 -4407
rect 330825 -4436 331499 -4407
rect 334169 -4436 334843 -4407
rect 337513 -4436 338187 -4407
rect 340857 -4436 341531 -4407
rect 344201 -4436 344875 -4407
rect 347545 -4436 348219 -4407
rect 350889 -4436 351563 -4407
rect 354233 -4436 354907 -4407
rect 357577 -4436 358251 -4407
rect 360921 -4436 361595 -4407
rect 364265 -4436 364939 -4407
rect 367609 -4436 368283 -4407
rect 370953 -4436 371627 -4407
rect 374297 -4436 374971 -4407
rect 377641 -4436 378315 -4407
rect 380985 -4436 381659 -4407
rect 384329 -4436 385003 -4407
rect 387673 -4436 388347 -4407
rect 391017 -4436 391691 -4407
rect 394361 -4436 395035 -4407
rect 397705 -4436 398379 -4407
rect 401049 -4436 401723 -4407
rect 404393 -4436 405067 -4407
rect 407737 -4436 408411 -4407
rect 411081 -4436 411755 -4407
rect 414425 -4436 415099 -4407
rect 417769 -4436 418443 -4407
rect 421113 -4436 421787 -4407
rect 424457 -4436 425131 -4407
rect 427801 -4436 428475 -4407
rect 218311 -4848 218358 -4483
rect 218365 -4848 218412 -4537
rect 220473 -4848 221206 -4436
rect 221655 -4848 221702 -4483
rect 221709 -4848 221756 -4537
rect 223817 -4848 224550 -4436
rect 224999 -4848 225046 -4483
rect 225053 -4848 225100 -4537
rect 227161 -4848 227894 -4436
rect 228343 -4848 228390 -4483
rect 228397 -4848 228444 -4537
rect 230505 -4848 231238 -4436
rect 231687 -4848 231734 -4483
rect 231741 -4848 231788 -4537
rect 233849 -4848 234582 -4436
rect 235031 -4848 235078 -4483
rect 235085 -4848 235132 -4537
rect 237193 -4848 237926 -4436
rect 238375 -4848 238422 -4483
rect 238429 -4848 238476 -4537
rect 240537 -4848 241270 -4436
rect 241719 -4848 241766 -4483
rect 241773 -4848 241820 -4537
rect 243881 -4848 244614 -4436
rect 245063 -4848 245110 -4483
rect 245117 -4848 245164 -4537
rect 247225 -4848 247958 -4436
rect 248407 -4848 248454 -4483
rect 248461 -4848 248508 -4537
rect 250569 -4848 251302 -4436
rect 251751 -4848 251798 -4483
rect 251805 -4848 251852 -4537
rect 253913 -4848 254646 -4436
rect 255095 -4848 255142 -4483
rect 255149 -4848 255196 -4537
rect 257257 -4848 257990 -4436
rect 258439 -4848 258486 -4483
rect 258493 -4848 258540 -4537
rect 260601 -4848 261334 -4436
rect 261783 -4848 261830 -4483
rect 261837 -4848 261884 -4537
rect 263945 -4848 264678 -4436
rect 265127 -4848 265174 -4483
rect 265181 -4848 265228 -4537
rect 267289 -4848 268022 -4436
rect 268471 -4848 268518 -4483
rect 268525 -4848 268572 -4537
rect 270633 -4848 271366 -4436
rect 271815 -4848 271862 -4483
rect 271869 -4848 271916 -4537
rect 273977 -4848 274710 -4436
rect 275159 -4848 275206 -4483
rect 275213 -4848 275260 -4537
rect 277321 -4848 278054 -4436
rect 278503 -4848 278550 -4483
rect 278557 -4848 278604 -4537
rect 280665 -4848 281398 -4436
rect 281847 -4848 281894 -4483
rect 281901 -4848 281948 -4537
rect 284009 -4848 284742 -4436
rect 285191 -4848 285238 -4483
rect 285245 -4848 285292 -4537
rect 287353 -4848 288086 -4436
rect 288535 -4848 288582 -4483
rect 288589 -4848 288636 -4537
rect 290697 -4848 291430 -4436
rect 291879 -4848 291926 -4483
rect 291933 -4848 291980 -4537
rect 294041 -4848 294774 -4436
rect 295223 -4848 295270 -4483
rect 295277 -4848 295324 -4537
rect 297385 -4848 298118 -4436
rect 298567 -4848 298614 -4483
rect 298621 -4848 298668 -4537
rect 300729 -4848 301462 -4436
rect 301911 -4848 301958 -4483
rect 301965 -4848 302012 -4537
rect 304073 -4848 304806 -4436
rect 305255 -4848 305302 -4483
rect 305309 -4848 305356 -4537
rect 307417 -4848 308150 -4436
rect 308599 -4848 308646 -4483
rect 308653 -4848 308700 -4537
rect 310761 -4848 311494 -4436
rect 311943 -4848 311990 -4483
rect 311997 -4848 312044 -4537
rect 314105 -4848 314838 -4436
rect 315287 -4848 315334 -4483
rect 315341 -4848 315388 -4537
rect 317449 -4848 318182 -4436
rect 318631 -4848 318678 -4483
rect 318685 -4848 318732 -4537
rect 320793 -4848 321526 -4436
rect 321975 -4848 322022 -4483
rect 322029 -4848 322076 -4537
rect 324137 -4848 324870 -4436
rect 325319 -4848 325366 -4483
rect 325373 -4848 325420 -4537
rect 327481 -4848 328214 -4436
rect 328663 -4848 328710 -4483
rect 328717 -4848 328764 -4537
rect 330825 -4848 331558 -4436
rect 332007 -4848 332054 -4483
rect 332061 -4848 332108 -4537
rect 334169 -4848 334902 -4436
rect 335351 -4848 335398 -4483
rect 335405 -4848 335452 -4537
rect 337513 -4848 338246 -4436
rect 338695 -4848 338742 -4483
rect 338749 -4848 338796 -4537
rect 340857 -4848 341590 -4436
rect 342039 -4848 342086 -4483
rect 342093 -4848 342140 -4537
rect 344201 -4848 344934 -4436
rect 345383 -4848 345430 -4483
rect 345437 -4848 345484 -4537
rect 347545 -4848 348278 -4436
rect 348727 -4848 348774 -4483
rect 348781 -4848 348828 -4537
rect 350889 -4848 351622 -4436
rect 352071 -4848 352118 -4483
rect 352125 -4848 352172 -4537
rect 354233 -4848 354966 -4436
rect 355415 -4848 355462 -4483
rect 355469 -4848 355516 -4537
rect 357577 -4848 358310 -4436
rect 358759 -4848 358806 -4483
rect 358813 -4848 358860 -4537
rect 360921 -4848 361654 -4436
rect 362103 -4848 362150 -4483
rect 362157 -4848 362204 -4537
rect 364265 -4848 364998 -4436
rect 365447 -4848 365494 -4483
rect 365501 -4848 365548 -4537
rect 367609 -4848 368342 -4436
rect 368791 -4848 368838 -4483
rect 368845 -4848 368892 -4537
rect 370953 -4848 371686 -4436
rect 372135 -4848 372182 -4483
rect 372189 -4848 372236 -4537
rect 374297 -4848 375030 -4436
rect 375479 -4848 375526 -4483
rect 375533 -4848 375580 -4537
rect 377641 -4848 378374 -4436
rect 378823 -4848 378870 -4483
rect 378877 -4848 378924 -4537
rect 380985 -4848 381718 -4436
rect 382167 -4848 382214 -4483
rect 382221 -4848 382268 -4537
rect 384329 -4848 385062 -4436
rect 385511 -4848 385558 -4483
rect 385565 -4848 385612 -4537
rect 387673 -4848 388406 -4436
rect 388855 -4848 388902 -4483
rect 388909 -4848 388956 -4537
rect 391017 -4848 391750 -4436
rect 392199 -4848 392246 -4483
rect 392253 -4848 392300 -4537
rect 394361 -4848 395094 -4436
rect 395543 -4848 395590 -4483
rect 395597 -4848 395644 -4537
rect 397705 -4848 398438 -4436
rect 398887 -4848 398934 -4483
rect 398941 -4848 398988 -4537
rect 401049 -4848 401782 -4436
rect 402231 -4848 402278 -4483
rect 402285 -4848 402332 -4537
rect 404393 -4848 405126 -4436
rect 405575 -4848 405622 -4483
rect 405629 -4848 405676 -4537
rect 407737 -4848 408470 -4436
rect 408919 -4848 408966 -4483
rect 408973 -4848 409020 -4537
rect 411081 -4848 411814 -4436
rect 412263 -4848 412310 -4483
rect 412317 -4848 412364 -4537
rect 414425 -4848 415158 -4436
rect 415607 -4848 415654 -4483
rect 415661 -4848 415708 -4537
rect 417769 -4848 418502 -4436
rect 418951 -4848 418998 -4483
rect 419005 -4848 419052 -4537
rect 421113 -4848 421846 -4436
rect 422295 -4848 422342 -4483
rect 422349 -4848 422396 -4537
rect 424457 -4848 425190 -4436
rect 425639 -4848 425686 -4483
rect 425693 -4848 425740 -4537
rect 427801 -4848 428534 -4436
rect 428983 -4848 429030 -4483
rect 429037 -4848 429084 -4537
rect 3131 -6087 5022 -6022
rect 6475 -6087 8366 -6022
rect 9819 -6087 11710 -6022
rect 13163 -6087 15054 -6022
rect 16507 -6087 18398 -6022
rect 19851 -6087 21742 -6022
rect 23195 -6087 25086 -6022
rect 26539 -6087 28430 -6022
rect 29883 -6087 31774 -6022
rect 33227 -6087 35118 -6022
rect 36571 -6087 38462 -6022
rect 39915 -6087 41806 -6022
rect 43259 -6087 45150 -6022
rect 46603 -6087 48494 -6022
rect 49947 -6087 51838 -6022
rect 53291 -6087 55182 -6022
rect 56635 -6087 58526 -6022
rect 59979 -6087 61870 -6022
rect 63323 -6087 65214 -6022
rect 66667 -6087 68558 -6022
rect 70011 -6087 71902 -6022
rect 73355 -6087 75246 -6022
rect 76699 -6087 78590 -6022
rect 80043 -6087 81934 -6022
rect 83387 -6087 85278 -6022
rect 86731 -6087 88622 -6022
rect 90075 -6087 91966 -6022
rect 93419 -6087 95310 -6022
rect 96763 -6087 98654 -6022
rect 100107 -6087 101998 -6022
rect 103451 -6087 105342 -6022
rect 106795 -6087 108686 -6022
rect 110139 -6087 112030 -6022
rect 113483 -6087 115374 -6022
rect 116827 -6087 118718 -6022
rect 120171 -6087 122062 -6022
rect 123515 -6087 125406 -6022
rect 126859 -6087 128750 -6022
rect 130203 -6087 132094 -6022
rect 133547 -6087 135438 -6022
rect 136891 -6087 138782 -6022
rect 140235 -6087 142126 -6022
rect 143579 -6087 145470 -6022
rect 146923 -6087 148814 -6022
rect 150267 -6087 152158 -6022
rect 153611 -6087 155502 -6022
rect 156955 -6087 158846 -6022
rect 160299 -6087 162190 -6022
rect 163643 -6087 165534 -6022
rect 166987 -6087 168878 -6022
rect 170331 -6087 172222 -6022
rect 173675 -6087 175566 -6022
rect 177019 -6087 178910 -6022
rect 180363 -6087 182254 -6022
rect 183707 -6087 185598 -6022
rect 187051 -6087 188942 -6022
rect 190395 -6087 192286 -6022
rect 193739 -6087 195630 -6022
rect 197083 -6087 198974 -6022
rect 200427 -6087 202318 -6022
rect 203771 -6087 205662 -6022
rect 207115 -6087 209006 -6022
rect 210459 -6087 211496 -6022
rect 3722 -6147 5022 -6087
rect 7066 -6147 8366 -6087
rect 10410 -6147 11710 -6087
rect 13754 -6147 15054 -6087
rect 17098 -6147 18398 -6087
rect 20442 -6147 21742 -6087
rect 23786 -6147 25086 -6087
rect 27130 -6147 28430 -6087
rect 30474 -6147 31774 -6087
rect 33818 -6147 35118 -6087
rect 37162 -6147 38462 -6087
rect 40506 -6147 41806 -6087
rect 43850 -6147 45150 -6087
rect 47194 -6147 48494 -6087
rect 50538 -6147 51838 -6087
rect 53882 -6147 55182 -6087
rect 57226 -6147 58526 -6087
rect 60570 -6147 61870 -6087
rect 63914 -6147 65214 -6087
rect 67258 -6147 68558 -6087
rect 70602 -6147 71902 -6087
rect 73946 -6147 75246 -6087
rect 77290 -6147 78590 -6087
rect 80634 -6147 81934 -6087
rect 83978 -6147 85278 -6087
rect 87322 -6147 88622 -6087
rect 90666 -6147 91966 -6087
rect 94010 -6147 95310 -6087
rect 97354 -6147 98654 -6087
rect 100698 -6147 101998 -6087
rect 104042 -6147 105342 -6087
rect 107386 -6147 108686 -6087
rect 110730 -6147 112030 -6087
rect 114074 -6147 115374 -6087
rect 117418 -6147 118718 -6087
rect 120762 -6147 122062 -6087
rect 124106 -6147 125406 -6087
rect 127450 -6147 128750 -6087
rect 130794 -6147 132094 -6087
rect 134138 -6147 135438 -6087
rect 137482 -6147 138782 -6087
rect 140826 -6147 142126 -6087
rect 144170 -6147 145470 -6087
rect 147514 -6147 148814 -6087
rect 150858 -6147 152158 -6087
rect 154202 -6147 155502 -6087
rect 157546 -6147 158846 -6087
rect 160890 -6147 162190 -6087
rect 164234 -6147 165534 -6087
rect 167578 -6147 168878 -6087
rect 170922 -6147 172222 -6087
rect 174266 -6147 175566 -6087
rect 177610 -6147 178910 -6087
rect 180954 -6147 182254 -6087
rect 184298 -6147 185598 -6087
rect 187642 -6147 188942 -6087
rect 190986 -6147 192286 -6087
rect 194330 -6147 195630 -6087
rect 197674 -6147 198974 -6087
rect 201018 -6147 202318 -6087
rect 204362 -6147 205662 -6087
rect 207706 -6147 209006 -6087
rect 211050 -6147 211496 -6087
rect 3751 -6152 5022 -6147
rect 7095 -6152 8366 -6147
rect 10439 -6152 11710 -6147
rect 13783 -6152 15054 -6147
rect 17127 -6152 18398 -6147
rect 20471 -6152 21742 -6147
rect 23815 -6152 25086 -6147
rect 27159 -6152 28430 -6147
rect 30503 -6152 31774 -6147
rect 33847 -6152 35118 -6147
rect 37191 -6152 38462 -6147
rect 40535 -6152 41806 -6147
rect 43879 -6152 45150 -6147
rect 47223 -6152 48494 -6147
rect 50567 -6152 51838 -6147
rect 53911 -6152 55182 -6147
rect 57255 -6152 58526 -6147
rect 60599 -6152 61870 -6147
rect 63943 -6152 65214 -6147
rect 67287 -6152 68558 -6147
rect 70631 -6152 71902 -6147
rect 73975 -6152 75246 -6147
rect 77319 -6152 78590 -6147
rect 80663 -6152 81934 -6147
rect 84007 -6152 85278 -6147
rect 87351 -6152 88622 -6147
rect 90695 -6152 91966 -6147
rect 94039 -6152 95310 -6147
rect 97383 -6152 98654 -6147
rect 100727 -6152 101998 -6147
rect 104071 -6152 105342 -6147
rect 107415 -6152 108686 -6147
rect 110759 -6152 112030 -6147
rect 114103 -6152 115374 -6147
rect 117447 -6152 118718 -6147
rect 120791 -6152 122062 -6147
rect 124135 -6152 125406 -6147
rect 127479 -6152 128750 -6147
rect 130823 -6152 132094 -6147
rect 134167 -6152 135438 -6147
rect 137511 -6152 138782 -6147
rect 140855 -6152 142126 -6147
rect 144199 -6152 145470 -6147
rect 147543 -6152 148814 -6147
rect 150887 -6152 152158 -6147
rect 154231 -6152 155502 -6147
rect 157575 -6152 158846 -6147
rect 160919 -6152 162190 -6147
rect 164263 -6152 165534 -6147
rect 167607 -6152 168878 -6147
rect 170951 -6152 172222 -6147
rect 174295 -6152 175566 -6147
rect 177639 -6152 178910 -6147
rect 180983 -6152 182254 -6147
rect 184327 -6152 185598 -6147
rect 187671 -6152 188942 -6147
rect 191015 -6152 192286 -6147
rect 194359 -6152 195630 -6147
rect 197703 -6152 198974 -6147
rect 201047 -6152 202318 -6147
rect 204391 -6152 205662 -6147
rect 207735 -6152 209006 -6147
rect 211079 -6152 211496 -6147
rect 3875 -6170 5022 -6152
rect 7219 -6170 8366 -6152
rect 10563 -6170 11710 -6152
rect 13907 -6170 15054 -6152
rect 17251 -6170 18398 -6152
rect 20595 -6170 21742 -6152
rect 23939 -6170 25086 -6152
rect 27283 -6170 28430 -6152
rect 30627 -6170 31774 -6152
rect 33971 -6170 35118 -6152
rect 37315 -6170 38462 -6152
rect 40659 -6170 41806 -6152
rect 44003 -6170 45150 -6152
rect 47347 -6170 48494 -6152
rect 50691 -6170 51838 -6152
rect 54035 -6170 55182 -6152
rect 57379 -6170 58526 -6152
rect 60723 -6170 61870 -6152
rect 64067 -6170 65214 -6152
rect 67411 -6170 68558 -6152
rect 70755 -6170 71902 -6152
rect 74099 -6170 75246 -6152
rect 77443 -6170 78590 -6152
rect 80787 -6170 81934 -6152
rect 84131 -6170 85278 -6152
rect 87475 -6170 88622 -6152
rect 90819 -6170 91966 -6152
rect 94163 -6170 95310 -6152
rect 97507 -6170 98654 -6152
rect 100851 -6170 101998 -6152
rect 104195 -6170 105342 -6152
rect 107539 -6170 108686 -6152
rect 110883 -6170 112030 -6152
rect 114227 -6170 115374 -6152
rect 117571 -6170 118718 -6152
rect 120915 -6170 122062 -6152
rect 124259 -6170 125406 -6152
rect 127603 -6170 128750 -6152
rect 130947 -6170 132094 -6152
rect 134291 -6170 135438 -6152
rect 137635 -6170 138782 -6152
rect 140979 -6170 142126 -6152
rect 144323 -6170 145470 -6152
rect 147667 -6170 148814 -6152
rect 151011 -6170 152158 -6152
rect 154355 -6170 155502 -6152
rect 157699 -6170 158846 -6152
rect 161043 -6170 162190 -6152
rect 164387 -6170 165534 -6152
rect 167731 -6170 168878 -6152
rect 171075 -6170 172222 -6152
rect 174419 -6170 175566 -6152
rect 177763 -6170 178910 -6152
rect 181107 -6170 182254 -6152
rect 184451 -6170 185598 -6152
rect 187795 -6170 188942 -6152
rect 191139 -6170 192286 -6152
rect 194483 -6170 195630 -6152
rect 197827 -6170 198974 -6152
rect 201171 -6170 202318 -6152
rect 204515 -6170 205662 -6152
rect 207859 -6170 209006 -6152
rect 211203 -6170 211641 -6152
rect 4313 -6181 5022 -6170
rect 7657 -6181 8366 -6170
rect 11001 -6181 11710 -6170
rect 14345 -6181 15054 -6170
rect 17689 -6181 18398 -6170
rect 21033 -6181 21742 -6170
rect 24377 -6181 25086 -6170
rect 27721 -6181 28430 -6170
rect 31065 -6181 31774 -6170
rect 34409 -6181 35118 -6170
rect 37753 -6181 38462 -6170
rect 41097 -6181 41806 -6170
rect 44441 -6181 45150 -6170
rect 47785 -6181 48494 -6170
rect 51129 -6181 51838 -6170
rect 54473 -6181 55182 -6170
rect 57817 -6181 58526 -6170
rect 61161 -6181 61870 -6170
rect 64505 -6181 65214 -6170
rect 67849 -6181 68558 -6170
rect 71193 -6181 71902 -6170
rect 74537 -6181 75246 -6170
rect 77881 -6181 78590 -6170
rect 81225 -6181 81934 -6170
rect 84569 -6181 85278 -6170
rect 87913 -6181 88622 -6170
rect 91257 -6181 91966 -6170
rect 94601 -6181 95310 -6170
rect 97945 -6181 98654 -6170
rect 101289 -6181 101998 -6170
rect 104633 -6181 105342 -6170
rect 107977 -6181 108686 -6170
rect 111321 -6181 112030 -6170
rect 114665 -6181 115374 -6170
rect 118009 -6181 118718 -6170
rect 121353 -6181 122062 -6170
rect 124697 -6181 125406 -6170
rect 128041 -6181 128750 -6170
rect 131385 -6181 132094 -6170
rect 134729 -6181 135438 -6170
rect 138073 -6181 138782 -6170
rect 141417 -6181 142126 -6170
rect 144761 -6181 145470 -6170
rect 148105 -6181 148814 -6170
rect 151449 -6181 152158 -6170
rect 154793 -6181 155502 -6170
rect 158137 -6181 158846 -6170
rect 161481 -6181 162190 -6170
rect 164825 -6181 165534 -6170
rect 168169 -6181 168878 -6170
rect 171513 -6181 172222 -6170
rect 174857 -6181 175566 -6170
rect 178201 -6181 178910 -6170
rect 181545 -6181 182254 -6170
rect 184889 -6181 185598 -6170
rect 188233 -6181 188942 -6170
rect 191577 -6181 192286 -6170
rect 194921 -6181 195630 -6170
rect 198265 -6181 198974 -6170
rect 201609 -6181 202318 -6170
rect 204953 -6181 205662 -6170
rect 208297 -6181 209006 -6170
rect 4313 -6217 4987 -6181
rect 7657 -6217 8331 -6181
rect 11001 -6217 11675 -6181
rect 14345 -6217 15019 -6181
rect 17689 -6217 18363 -6181
rect 21033 -6217 21707 -6181
rect 24377 -6217 25051 -6181
rect 27721 -6217 28395 -6181
rect 31065 -6217 31739 -6181
rect 34409 -6217 35083 -6181
rect 37753 -6217 38427 -6181
rect 41097 -6217 41771 -6181
rect 44441 -6217 45115 -6181
rect 47785 -6217 48459 -6181
rect 51129 -6217 51803 -6181
rect 54473 -6217 55147 -6181
rect 57817 -6217 58491 -6181
rect 61161 -6217 61835 -6181
rect 64505 -6217 65179 -6181
rect 67849 -6217 68523 -6181
rect 71193 -6217 71867 -6181
rect 74537 -6217 75211 -6181
rect 77881 -6217 78555 -6181
rect 81225 -6217 81899 -6181
rect 84569 -6217 85243 -6181
rect 87913 -6217 88587 -6181
rect 91257 -6217 91931 -6181
rect 94601 -6217 95275 -6181
rect 97945 -6217 98619 -6181
rect 101289 -6217 101963 -6181
rect 104633 -6217 105307 -6181
rect 107977 -6217 108651 -6181
rect 111321 -6217 111995 -6181
rect 114665 -6217 115339 -6181
rect 118009 -6217 118683 -6181
rect 121353 -6217 122027 -6181
rect 124697 -6217 125371 -6181
rect 128041 -6217 128715 -6181
rect 131385 -6217 132059 -6181
rect 134729 -6217 135403 -6181
rect 138073 -6217 138747 -6181
rect 141417 -6217 142091 -6181
rect 144761 -6217 145435 -6181
rect 148105 -6217 148779 -6181
rect 151449 -6217 152123 -6181
rect 154793 -6217 155467 -6181
rect 158137 -6217 158811 -6181
rect 161481 -6217 162155 -6181
rect 164825 -6217 165499 -6181
rect 168169 -6217 168843 -6181
rect 171513 -6217 172187 -6181
rect 174857 -6217 175531 -6181
rect 178201 -6217 178875 -6181
rect 181545 -6217 182219 -6181
rect 184889 -6217 185563 -6181
rect 188233 -6217 188907 -6181
rect 191577 -6217 192251 -6181
rect 194921 -6217 195595 -6181
rect 198265 -6217 198939 -6181
rect 201609 -6217 202283 -6181
rect 204953 -6217 205627 -6181
rect 208297 -6217 208971 -6181
rect 212297 -6181 212350 -5067
rect 218280 -4943 218483 -4848
rect 220473 -4906 221827 -4848
rect 223817 -4906 225171 -4848
rect 227161 -4906 228515 -4848
rect 230505 -4906 231859 -4848
rect 233849 -4906 235203 -4848
rect 237193 -4906 238547 -4848
rect 240537 -4906 241891 -4848
rect 243881 -4906 245235 -4848
rect 247225 -4906 248579 -4848
rect 250569 -4906 251923 -4848
rect 253913 -4906 255267 -4848
rect 257257 -4906 258611 -4848
rect 260601 -4906 261955 -4848
rect 263945 -4906 265299 -4848
rect 267289 -4906 268643 -4848
rect 270633 -4906 271987 -4848
rect 273977 -4906 275331 -4848
rect 277321 -4906 278675 -4848
rect 280665 -4906 282019 -4848
rect 284009 -4906 285363 -4848
rect 287353 -4906 288707 -4848
rect 290697 -4906 292051 -4848
rect 294041 -4906 295395 -4848
rect 297385 -4906 298739 -4848
rect 300729 -4906 302083 -4848
rect 304073 -4906 305427 -4848
rect 307417 -4906 308771 -4848
rect 310761 -4906 312115 -4848
rect 314105 -4906 315459 -4848
rect 317449 -4906 318803 -4848
rect 320793 -4906 322147 -4848
rect 324137 -4906 325491 -4848
rect 327481 -4906 328835 -4848
rect 330825 -4906 332179 -4848
rect 334169 -4906 335523 -4848
rect 337513 -4906 338867 -4848
rect 340857 -4906 342211 -4848
rect 344201 -4906 345555 -4848
rect 347545 -4906 348899 -4848
rect 350889 -4906 352243 -4848
rect 354233 -4906 355587 -4848
rect 357577 -4906 358931 -4848
rect 360921 -4906 362275 -4848
rect 364265 -4906 365619 -4848
rect 367609 -4906 368963 -4848
rect 370953 -4906 372307 -4848
rect 374297 -4906 375651 -4848
rect 377641 -4906 378995 -4848
rect 380985 -4906 382339 -4848
rect 384329 -4906 385683 -4848
rect 387673 -4906 389027 -4848
rect 391017 -4906 392371 -4848
rect 394361 -4906 395715 -4848
rect 397705 -4906 399059 -4848
rect 401049 -4906 402403 -4848
rect 404393 -4906 405747 -4848
rect 407737 -4906 409091 -4848
rect 411081 -4906 412435 -4848
rect 414425 -4906 415779 -4848
rect 417769 -4906 419123 -4848
rect 421113 -4906 422467 -4848
rect 424457 -4906 425811 -4848
rect 427801 -4906 429155 -4848
rect 219900 -4943 221827 -4906
rect 223244 -4943 225171 -4906
rect 226588 -4943 228515 -4906
rect 229932 -4943 231859 -4906
rect 233276 -4943 235203 -4906
rect 236620 -4943 238547 -4906
rect 239964 -4943 241891 -4906
rect 243308 -4943 245235 -4906
rect 246652 -4943 248579 -4906
rect 249996 -4943 251923 -4906
rect 253340 -4943 255267 -4906
rect 256684 -4943 258611 -4906
rect 260028 -4943 261955 -4906
rect 263372 -4943 265299 -4906
rect 266716 -4943 268643 -4906
rect 270060 -4943 271987 -4906
rect 273404 -4943 275331 -4906
rect 276748 -4943 278675 -4906
rect 280092 -4943 282019 -4906
rect 283436 -4943 285363 -4906
rect 286780 -4943 288707 -4906
rect 290124 -4943 292051 -4906
rect 293468 -4943 295395 -4906
rect 296812 -4943 298739 -4906
rect 300156 -4943 302083 -4906
rect 303500 -4943 305427 -4906
rect 306844 -4943 308771 -4906
rect 310188 -4943 312115 -4906
rect 313532 -4943 315459 -4906
rect 316876 -4943 318803 -4906
rect 320220 -4943 322147 -4906
rect 323564 -4943 325491 -4906
rect 326908 -4943 328835 -4906
rect 330252 -4943 332179 -4906
rect 333596 -4943 335523 -4906
rect 336940 -4943 338867 -4906
rect 340284 -4943 342211 -4906
rect 343628 -4943 345555 -4906
rect 346972 -4943 348899 -4906
rect 350316 -4943 352243 -4906
rect 353660 -4943 355587 -4906
rect 357004 -4943 358931 -4906
rect 360348 -4943 362275 -4906
rect 363692 -4943 365619 -4906
rect 367036 -4943 368963 -4906
rect 370380 -4943 372307 -4906
rect 373724 -4943 375651 -4906
rect 377068 -4943 378995 -4906
rect 380412 -4943 382339 -4906
rect 383756 -4943 385683 -4906
rect 387100 -4943 389027 -4906
rect 390444 -4943 392371 -4906
rect 393788 -4943 395715 -4906
rect 397132 -4943 399059 -4906
rect 400476 -4943 402403 -4906
rect 403820 -4943 405747 -4906
rect 407164 -4943 409091 -4906
rect 410508 -4943 412435 -4906
rect 413852 -4943 415779 -4906
rect 417196 -4943 419123 -4906
rect 420540 -4943 422467 -4906
rect 423884 -4943 425811 -4906
rect 427228 -4943 429155 -4906
rect 218280 -5067 218985 -4943
rect 219900 -5067 222329 -4943
rect 223244 -5067 225673 -4943
rect 226588 -5067 229017 -4943
rect 229932 -5067 232361 -4943
rect 233276 -5067 235705 -4943
rect 236620 -5067 239049 -4943
rect 239964 -5067 242393 -4943
rect 243308 -5067 245737 -4943
rect 246652 -5067 249081 -4943
rect 249996 -5067 252425 -4943
rect 253340 -5067 255769 -4943
rect 256684 -5067 259113 -4943
rect 260028 -5067 262457 -4943
rect 263372 -5067 265801 -4943
rect 266716 -5067 269145 -4943
rect 270060 -5067 272489 -4943
rect 273404 -5067 275833 -4943
rect 276748 -5067 279177 -4943
rect 280092 -5067 282521 -4943
rect 283436 -5067 285865 -4943
rect 286780 -5067 289209 -4943
rect 290124 -5067 292553 -4943
rect 293468 -5067 295897 -4943
rect 296812 -5067 299241 -4943
rect 300156 -5067 302585 -4943
rect 303500 -5067 305929 -4943
rect 306844 -5067 309273 -4943
rect 310188 -5067 312617 -4943
rect 313532 -5067 315961 -4943
rect 316876 -5067 319305 -4943
rect 320220 -5067 322649 -4943
rect 323564 -5067 325993 -4943
rect 326908 -5067 329337 -4943
rect 330252 -5067 332681 -4943
rect 333596 -5067 336025 -4943
rect 336940 -5067 339369 -4943
rect 340284 -5067 342713 -4943
rect 343628 -5067 346057 -4943
rect 346972 -5067 349401 -4943
rect 350316 -5067 352745 -4943
rect 353660 -5067 356089 -4943
rect 357004 -5067 359433 -4943
rect 360348 -5067 362777 -4943
rect 363692 -5067 366121 -4943
rect 367036 -5067 369465 -4943
rect 370380 -5067 372809 -4943
rect 373724 -5067 376153 -4943
rect 377068 -5067 379497 -4943
rect 380412 -5067 382841 -4943
rect 383756 -5067 386185 -4943
rect 387100 -5067 389529 -4943
rect 390444 -5067 392873 -4943
rect 393788 -5067 396217 -4943
rect 397132 -5067 399561 -4943
rect 400476 -5067 402905 -4943
rect 403820 -5067 406249 -4943
rect 407164 -5067 409593 -4943
rect 410508 -5067 412937 -4943
rect 413852 -5067 416281 -4943
rect 417196 -5067 419625 -4943
rect 420540 -5067 422969 -4943
rect 423884 -5067 426313 -4943
rect 427228 -5067 429657 -4943
rect 218280 -6152 219038 -5067
rect 219900 -6022 222382 -5067
rect 223244 -6022 225726 -5067
rect 226588 -6022 229070 -5067
rect 229932 -6022 232414 -5067
rect 233276 -6022 235758 -5067
rect 236620 -6022 239102 -5067
rect 239964 -6022 242446 -5067
rect 243308 -6022 245790 -5067
rect 246652 -6022 249134 -5067
rect 249996 -6022 252478 -5067
rect 253340 -6022 255822 -5067
rect 256684 -6022 259166 -5067
rect 260028 -6022 262510 -5067
rect 263372 -6022 265854 -5067
rect 266716 -6022 269198 -5067
rect 270060 -6022 272542 -5067
rect 273404 -6022 275886 -5067
rect 276748 -6022 279230 -5067
rect 280092 -6022 282574 -5067
rect 283436 -6022 285918 -5067
rect 286780 -6022 289262 -5067
rect 290124 -6022 292606 -5067
rect 293468 -6022 295950 -5067
rect 296812 -6022 299294 -5067
rect 300156 -6022 302638 -5067
rect 303500 -6022 305982 -5067
rect 306844 -6022 309326 -5067
rect 310188 -6022 312670 -5067
rect 313532 -6022 316014 -5067
rect 316876 -6022 319358 -5067
rect 320220 -6022 322702 -5067
rect 323564 -6022 326046 -5067
rect 326908 -6022 329390 -5067
rect 330252 -6022 332734 -5067
rect 333596 -6022 336078 -5067
rect 336940 -6022 339422 -5067
rect 340284 -6022 342766 -5067
rect 343628 -6022 346110 -5067
rect 346972 -6022 349454 -5067
rect 350316 -6022 352798 -5067
rect 353660 -6022 356142 -5067
rect 357004 -6022 359486 -5067
rect 360348 -6022 362830 -5067
rect 363692 -6022 366174 -5067
rect 367036 -6022 369518 -5067
rect 370380 -6022 372862 -5067
rect 373724 -6022 376206 -5067
rect 377068 -6022 379550 -5067
rect 380412 -6022 382894 -5067
rect 383756 -6022 386238 -5067
rect 387100 -6022 389582 -5067
rect 390444 -6022 392926 -5067
rect 393788 -6022 396270 -5067
rect 397132 -6022 399614 -5067
rect 400476 -6022 402958 -5067
rect 403820 -6022 406302 -5067
rect 407164 -6022 409646 -5067
rect 410508 -6022 412990 -5067
rect 413852 -6022 416334 -5067
rect 417196 -6022 419678 -5067
rect 420540 -6022 423022 -5067
rect 423884 -6022 426366 -5067
rect 427228 -6022 429710 -5067
rect 220491 -6087 222382 -6022
rect 223835 -6087 225726 -6022
rect 227179 -6087 229070 -6022
rect 230523 -6087 232414 -6022
rect 233867 -6087 235758 -6022
rect 237211 -6087 239102 -6022
rect 240555 -6087 242446 -6022
rect 243899 -6087 245790 -6022
rect 247243 -6087 249134 -6022
rect 250587 -6087 252478 -6022
rect 253931 -6087 255822 -6022
rect 257275 -6087 259166 -6022
rect 260619 -6087 262510 -6022
rect 263963 -6087 265854 -6022
rect 267307 -6087 269198 -6022
rect 270651 -6087 272542 -6022
rect 273995 -6087 275886 -6022
rect 277339 -6087 279230 -6022
rect 280683 -6087 282574 -6022
rect 284027 -6087 285918 -6022
rect 287371 -6087 289262 -6022
rect 290715 -6087 292606 -6022
rect 294059 -6087 295950 -6022
rect 297403 -6087 299294 -6022
rect 300747 -6087 302638 -6022
rect 304091 -6087 305982 -6022
rect 307435 -6087 309326 -6022
rect 310779 -6087 312670 -6022
rect 314123 -6087 316014 -6022
rect 317467 -6087 319358 -6022
rect 320811 -6087 322702 -6022
rect 324155 -6087 326046 -6022
rect 327499 -6087 329390 -6022
rect 330843 -6087 332734 -6022
rect 334187 -6087 336078 -6022
rect 337531 -6087 339422 -6022
rect 340875 -6087 342766 -6022
rect 344219 -6087 346110 -6022
rect 347563 -6087 349454 -6022
rect 350907 -6087 352798 -6022
rect 354251 -6087 356142 -6022
rect 357595 -6087 359486 -6022
rect 360939 -6087 362830 -6022
rect 364283 -6087 366174 -6022
rect 367627 -6087 369518 -6022
rect 370971 -6087 372862 -6022
rect 374315 -6087 376206 -6022
rect 377659 -6087 379550 -6022
rect 381003 -6087 382894 -6022
rect 384347 -6087 386238 -6022
rect 387691 -6087 389582 -6022
rect 391035 -6087 392926 -6022
rect 394379 -6087 396270 -6022
rect 397723 -6087 399614 -6022
rect 401067 -6087 402958 -6022
rect 404411 -6087 406302 -6022
rect 407755 -6087 409646 -6022
rect 411099 -6087 412990 -6022
rect 414443 -6087 416334 -6022
rect 417787 -6087 419678 -6022
rect 421131 -6087 423022 -6022
rect 424475 -6087 426366 -6022
rect 427819 -6087 429710 -6022
rect 221082 -6147 222382 -6087
rect 224426 -6147 225726 -6087
rect 227770 -6147 229070 -6087
rect 231114 -6147 232414 -6087
rect 234458 -6147 235758 -6087
rect 237802 -6147 239102 -6087
rect 241146 -6147 242446 -6087
rect 244490 -6147 245790 -6087
rect 247834 -6147 249134 -6087
rect 251178 -6147 252478 -6087
rect 254522 -6147 255822 -6087
rect 257866 -6147 259166 -6087
rect 261210 -6147 262510 -6087
rect 264554 -6147 265854 -6087
rect 267898 -6147 269198 -6087
rect 271242 -6147 272542 -6087
rect 274586 -6147 275886 -6087
rect 277930 -6147 279230 -6087
rect 281274 -6147 282574 -6087
rect 284618 -6147 285918 -6087
rect 287962 -6147 289262 -6087
rect 291306 -6147 292606 -6087
rect 294650 -6147 295950 -6087
rect 297994 -6147 299294 -6087
rect 301338 -6147 302638 -6087
rect 304682 -6147 305982 -6087
rect 308026 -6147 309326 -6087
rect 311370 -6147 312670 -6087
rect 314714 -6147 316014 -6087
rect 318058 -6147 319358 -6087
rect 321402 -6147 322702 -6087
rect 324746 -6147 326046 -6087
rect 328090 -6147 329390 -6087
rect 331434 -6147 332734 -6087
rect 334778 -6147 336078 -6087
rect 338122 -6147 339422 -6087
rect 341466 -6147 342766 -6087
rect 344810 -6147 346110 -6087
rect 348154 -6147 349454 -6087
rect 351498 -6147 352798 -6087
rect 354842 -6147 356142 -6087
rect 358186 -6147 359486 -6087
rect 361530 -6147 362830 -6087
rect 364874 -6147 366174 -6087
rect 368218 -6147 369518 -6087
rect 371562 -6147 372862 -6087
rect 374906 -6147 376206 -6087
rect 378250 -6147 379550 -6087
rect 381594 -6147 382894 -6087
rect 384938 -6147 386238 -6087
rect 388282 -6147 389582 -6087
rect 391626 -6147 392926 -6087
rect 394970 -6147 396270 -6087
rect 398314 -6147 399614 -6087
rect 401658 -6147 402958 -6087
rect 405002 -6147 406302 -6087
rect 408346 -6147 409646 -6087
rect 411690 -6147 412990 -6087
rect 415034 -6147 416334 -6087
rect 418378 -6147 419678 -6087
rect 421722 -6147 423022 -6087
rect 425066 -6147 426366 -6087
rect 428410 -6147 429710 -6087
rect 221111 -6152 222382 -6147
rect 224455 -6152 225726 -6147
rect 227799 -6152 229070 -6147
rect 231143 -6152 232414 -6147
rect 234487 -6152 235758 -6147
rect 237831 -6152 239102 -6147
rect 241175 -6152 242446 -6147
rect 244519 -6152 245790 -6147
rect 247863 -6152 249134 -6147
rect 251207 -6152 252478 -6147
rect 254551 -6152 255822 -6147
rect 257895 -6152 259166 -6147
rect 261239 -6152 262510 -6147
rect 264583 -6152 265854 -6147
rect 267927 -6152 269198 -6147
rect 271271 -6152 272542 -6147
rect 274615 -6152 275886 -6147
rect 277959 -6152 279230 -6147
rect 281303 -6152 282574 -6147
rect 284647 -6152 285918 -6147
rect 287991 -6152 289262 -6147
rect 291335 -6152 292606 -6147
rect 294679 -6152 295950 -6147
rect 298023 -6152 299294 -6147
rect 301367 -6152 302638 -6147
rect 304711 -6152 305982 -6147
rect 308055 -6152 309326 -6147
rect 311399 -6152 312670 -6147
rect 314743 -6152 316014 -6147
rect 318087 -6152 319358 -6147
rect 321431 -6152 322702 -6147
rect 324775 -6152 326046 -6147
rect 328119 -6152 329390 -6147
rect 331463 -6152 332734 -6147
rect 334807 -6152 336078 -6147
rect 338151 -6152 339422 -6147
rect 341495 -6152 342766 -6147
rect 344839 -6152 346110 -6147
rect 348183 -6152 349454 -6147
rect 351527 -6152 352798 -6147
rect 354871 -6152 356142 -6147
rect 358215 -6152 359486 -6147
rect 361559 -6152 362830 -6147
rect 364903 -6152 366174 -6147
rect 368247 -6152 369518 -6147
rect 371591 -6152 372862 -6147
rect 374935 -6152 376206 -6147
rect 378279 -6152 379550 -6147
rect 381623 -6152 382894 -6147
rect 384967 -6152 386238 -6147
rect 388311 -6152 389582 -6147
rect 391655 -6152 392926 -6147
rect 394999 -6152 396270 -6147
rect 398343 -6152 399614 -6147
rect 401687 -6152 402958 -6147
rect 405031 -6152 406302 -6147
rect 408375 -6152 409646 -6147
rect 411719 -6152 412990 -6147
rect 415063 -6152 416334 -6147
rect 418407 -6152 419678 -6147
rect 421751 -6152 423022 -6147
rect 425095 -6152 426366 -6147
rect 428439 -6152 429710 -6147
rect 217891 -6170 219038 -6152
rect 221235 -6170 222382 -6152
rect 224579 -6170 225726 -6152
rect 227923 -6170 229070 -6152
rect 231267 -6170 232414 -6152
rect 234611 -6170 235758 -6152
rect 237955 -6170 239102 -6152
rect 241299 -6170 242446 -6152
rect 244643 -6170 245790 -6152
rect 247987 -6170 249134 -6152
rect 251331 -6170 252478 -6152
rect 254675 -6170 255822 -6152
rect 258019 -6170 259166 -6152
rect 261363 -6170 262510 -6152
rect 264707 -6170 265854 -6152
rect 268051 -6170 269198 -6152
rect 271395 -6170 272542 -6152
rect 274739 -6170 275886 -6152
rect 278083 -6170 279230 -6152
rect 281427 -6170 282574 -6152
rect 284771 -6170 285918 -6152
rect 288115 -6170 289262 -6152
rect 291459 -6170 292606 -6152
rect 294803 -6170 295950 -6152
rect 298147 -6170 299294 -6152
rect 301491 -6170 302638 -6152
rect 304835 -6170 305982 -6152
rect 308179 -6170 309326 -6152
rect 311523 -6170 312670 -6152
rect 314867 -6170 316014 -6152
rect 318211 -6170 319358 -6152
rect 321555 -6170 322702 -6152
rect 324899 -6170 326046 -6152
rect 328243 -6170 329390 -6152
rect 331587 -6170 332734 -6152
rect 334931 -6170 336078 -6152
rect 338275 -6170 339422 -6152
rect 341619 -6170 342766 -6152
rect 344963 -6170 346110 -6152
rect 348307 -6170 349454 -6152
rect 351651 -6170 352798 -6152
rect 354995 -6170 356142 -6152
rect 358339 -6170 359486 -6152
rect 361683 -6170 362830 -6152
rect 365027 -6170 366174 -6152
rect 368371 -6170 369518 -6152
rect 371715 -6170 372862 -6152
rect 375059 -6170 376206 -6152
rect 378403 -6170 379550 -6152
rect 381747 -6170 382894 -6152
rect 385091 -6170 386238 -6152
rect 388435 -6170 389582 -6152
rect 391779 -6170 392926 -6152
rect 395123 -6170 396270 -6152
rect 398467 -6170 399614 -6152
rect 401811 -6170 402958 -6152
rect 405155 -6170 406302 -6152
rect 408499 -6170 409646 -6152
rect 411843 -6170 412990 -6152
rect 415187 -6170 416334 -6152
rect 418531 -6170 419678 -6152
rect 421875 -6170 423022 -6152
rect 425219 -6170 426366 -6152
rect 428563 -6170 429710 -6152
rect 218329 -6181 219038 -6170
rect 221673 -6181 222382 -6170
rect 225017 -6181 225726 -6170
rect 228361 -6181 229070 -6170
rect 231705 -6181 232414 -6170
rect 235049 -6181 235758 -6170
rect 238393 -6181 239102 -6170
rect 241737 -6181 242446 -6170
rect 245081 -6181 245790 -6170
rect 248425 -6181 249134 -6170
rect 251769 -6181 252478 -6170
rect 255113 -6181 255822 -6170
rect 258457 -6181 259166 -6170
rect 261801 -6181 262510 -6170
rect 265145 -6181 265854 -6170
rect 268489 -6181 269198 -6170
rect 271833 -6181 272542 -6170
rect 275177 -6181 275886 -6170
rect 278521 -6181 279230 -6170
rect 281865 -6181 282574 -6170
rect 285209 -6181 285918 -6170
rect 288553 -6181 289262 -6170
rect 291897 -6181 292606 -6170
rect 295241 -6181 295950 -6170
rect 298585 -6181 299294 -6170
rect 301929 -6181 302638 -6170
rect 305273 -6181 305982 -6170
rect 308617 -6181 309326 -6170
rect 311961 -6181 312670 -6170
rect 315305 -6181 316014 -6170
rect 318649 -6181 319358 -6170
rect 321993 -6181 322702 -6170
rect 325337 -6181 326046 -6170
rect 328681 -6181 329390 -6170
rect 332025 -6181 332734 -6170
rect 335369 -6181 336078 -6170
rect 338713 -6181 339422 -6170
rect 342057 -6181 342766 -6170
rect 345401 -6181 346110 -6170
rect 348745 -6181 349454 -6170
rect 352089 -6181 352798 -6170
rect 355433 -6181 356142 -6170
rect 358777 -6181 359486 -6170
rect 362121 -6181 362830 -6170
rect 365465 -6181 366174 -6170
rect 368809 -6181 369518 -6170
rect 372153 -6181 372862 -6170
rect 375497 -6181 376206 -6170
rect 378841 -6181 379550 -6170
rect 382185 -6181 382894 -6170
rect 385529 -6181 386238 -6170
rect 388873 -6181 389582 -6170
rect 392217 -6181 392926 -6170
rect 395561 -6181 396270 -6170
rect 398905 -6181 399614 -6170
rect 402249 -6181 402958 -6170
rect 405593 -6181 406302 -6170
rect 408937 -6181 409646 -6170
rect 412281 -6181 412990 -6170
rect 415625 -6181 416334 -6170
rect 418969 -6181 419678 -6170
rect 422313 -6181 423022 -6170
rect 425657 -6181 426366 -6170
rect 429001 -6181 429710 -6170
rect 212297 -6217 212315 -6181
rect 218329 -6217 219003 -6181
rect 221673 -6217 222347 -6181
rect 225017 -6217 225691 -6181
rect 228361 -6217 229035 -6181
rect 231705 -6217 232379 -6181
rect 235049 -6217 235723 -6181
rect 238393 -6217 239067 -6181
rect 241737 -6217 242411 -6181
rect 245081 -6217 245755 -6181
rect 248425 -6217 249099 -6181
rect 251769 -6217 252443 -6181
rect 255113 -6217 255787 -6181
rect 258457 -6217 259131 -6181
rect 261801 -6217 262475 -6181
rect 265145 -6217 265819 -6181
rect 268489 -6217 269163 -6181
rect 271833 -6217 272507 -6181
rect 275177 -6217 275851 -6181
rect 278521 -6217 279195 -6181
rect 281865 -6217 282539 -6181
rect 285209 -6217 285883 -6181
rect 288553 -6217 289227 -6181
rect 291897 -6217 292571 -6181
rect 295241 -6217 295915 -6181
rect 298585 -6217 299259 -6181
rect 301929 -6217 302603 -6181
rect 305273 -6217 305947 -6181
rect 308617 -6217 309291 -6181
rect 311961 -6217 312635 -6181
rect 315305 -6217 315979 -6181
rect 318649 -6217 319323 -6181
rect 321993 -6217 322667 -6181
rect 325337 -6217 326011 -6181
rect 328681 -6217 329355 -6181
rect 332025 -6217 332699 -6181
rect 335369 -6217 336043 -6181
rect 338713 -6217 339387 -6181
rect 342057 -6217 342731 -6181
rect 345401 -6217 346075 -6181
rect 348745 -6217 349419 -6181
rect 352089 -6217 352763 -6181
rect 355433 -6217 356107 -6181
rect 358777 -6217 359451 -6181
rect 362121 -6217 362795 -6181
rect 365465 -6217 366139 -6181
rect 368809 -6217 369483 -6181
rect 372153 -6217 372827 -6181
rect 375497 -6217 376171 -6181
rect 378841 -6217 379515 -6181
rect 382185 -6217 382859 -6181
rect 385529 -6217 386203 -6181
rect 388873 -6217 389547 -6181
rect 392217 -6217 392891 -6181
rect 395561 -6217 396235 -6181
rect 398905 -6217 399579 -6181
rect 402249 -6217 402923 -6181
rect 405593 -6217 406267 -6181
rect 408937 -6217 409611 -6181
rect 412281 -6217 412955 -6181
rect 415625 -6217 416299 -6181
rect 418969 -6217 419643 -6181
rect 422313 -6217 422987 -6181
rect 425657 -6217 426331 -6181
rect 429001 -6217 429675 -6181
rect 4496 -6235 4987 -6217
rect 7840 -6235 8331 -6217
rect 11184 -6235 11675 -6217
rect 14528 -6235 15019 -6217
rect 17872 -6235 18363 -6217
rect 21216 -6235 21707 -6217
rect 24560 -6235 25051 -6217
rect 27904 -6235 28395 -6217
rect 31248 -6235 31739 -6217
rect 34592 -6235 35083 -6217
rect 37936 -6235 38427 -6217
rect 41280 -6235 41771 -6217
rect 44624 -6235 45115 -6217
rect 47968 -6235 48459 -6217
rect 51312 -6235 51803 -6217
rect 54656 -6235 55147 -6217
rect 58000 -6235 58491 -6217
rect 61344 -6235 61835 -6217
rect 64688 -6235 65179 -6217
rect 68032 -6235 68523 -6217
rect 71376 -6235 71867 -6217
rect 74720 -6235 75211 -6217
rect 78064 -6235 78555 -6217
rect 81408 -6235 81899 -6217
rect 84752 -6235 85243 -6217
rect 88096 -6235 88587 -6217
rect 91440 -6235 91931 -6217
rect 94784 -6235 95275 -6217
rect 98128 -6235 98619 -6217
rect 101472 -6235 101963 -6217
rect 104816 -6235 105307 -6217
rect 108160 -6235 108651 -6217
rect 111504 -6235 111995 -6217
rect 114848 -6235 115339 -6217
rect 118192 -6235 118683 -6217
rect 121536 -6235 122027 -6217
rect 124880 -6235 125371 -6217
rect 128224 -6235 128715 -6217
rect 131568 -6235 132059 -6217
rect 134912 -6235 135403 -6217
rect 138256 -6235 138747 -6217
rect 141600 -6235 142091 -6217
rect 144944 -6235 145435 -6217
rect 148288 -6235 148779 -6217
rect 151632 -6235 152123 -6217
rect 154976 -6235 155467 -6217
rect 158320 -6235 158811 -6217
rect 161664 -6235 162155 -6217
rect 165008 -6235 165499 -6217
rect 168352 -6235 168843 -6217
rect 171696 -6235 172187 -6217
rect 175040 -6235 175531 -6217
rect 178384 -6235 178875 -6217
rect 181728 -6235 182219 -6217
rect 185072 -6235 185563 -6217
rect 188416 -6235 188907 -6217
rect 191760 -6235 192251 -6217
rect 195104 -6235 195595 -6217
rect 198448 -6235 198939 -6217
rect 201792 -6235 202283 -6217
rect 205136 -6235 205627 -6217
rect 208480 -6235 208971 -6217
rect 211824 -6235 212315 -6217
rect 218512 -6235 219003 -6217
rect 221856 -6235 222347 -6217
rect 225200 -6235 225691 -6217
rect 228544 -6235 229035 -6217
rect 231888 -6235 232379 -6217
rect 235232 -6235 235723 -6217
rect 238576 -6235 239067 -6217
rect 241920 -6235 242411 -6217
rect 245264 -6235 245755 -6217
rect 248608 -6235 249099 -6217
rect 251952 -6235 252443 -6217
rect 255296 -6235 255787 -6217
rect 258640 -6235 259131 -6217
rect 261984 -6235 262475 -6217
rect 265328 -6235 265819 -6217
rect 268672 -6235 269163 -6217
rect 272016 -6235 272507 -6217
rect 275360 -6235 275851 -6217
rect 278704 -6235 279195 -6217
rect 282048 -6235 282539 -6217
rect 285392 -6235 285883 -6217
rect 288736 -6235 289227 -6217
rect 292080 -6235 292571 -6217
rect 295424 -6235 295915 -6217
rect 298768 -6235 299259 -6217
rect 302112 -6235 302603 -6217
rect 305456 -6235 305947 -6217
rect 308800 -6235 309291 -6217
rect 312144 -6235 312635 -6217
rect 315488 -6235 315979 -6217
rect 318832 -6235 319323 -6217
rect 322176 -6235 322667 -6217
rect 325520 -6235 326011 -6217
rect 328864 -6235 329355 -6217
rect 332208 -6235 332699 -6217
rect 335552 -6235 336043 -6217
rect 338896 -6235 339387 -6217
rect 342240 -6235 342731 -6217
rect 345584 -6235 346075 -6217
rect 348928 -6235 349419 -6217
rect 352272 -6235 352763 -6217
rect 355616 -6235 356107 -6217
rect 358960 -6235 359451 -6217
rect 362304 -6235 362795 -6217
rect 365648 -6235 366139 -6217
rect 368992 -6235 369483 -6217
rect 372336 -6235 372827 -6217
rect 375680 -6235 376171 -6217
rect 379024 -6235 379515 -6217
rect 382368 -6235 382859 -6217
rect 385712 -6235 386203 -6217
rect 389056 -6235 389547 -6217
rect 392400 -6235 392891 -6217
rect 395744 -6235 396235 -6217
rect 399088 -6235 399579 -6217
rect 402432 -6235 402923 -6217
rect 405776 -6235 406267 -6217
rect 409120 -6235 409611 -6217
rect 412464 -6235 412955 -6217
rect 415808 -6235 416299 -6217
rect 419152 -6235 419643 -6217
rect 422496 -6235 422987 -6217
rect 425840 -6235 426331 -6217
rect 429184 -6235 429675 -6217
<< error_s >>
rect 214016 -2965 214132 -2899
rect 214132 -3219 214518 -3153
rect 213868 -3232 213878 -3219
rect 213802 -3274 213878 -3232
rect 213930 -3274 214518 -3219
rect 213802 -3277 214518 -3274
rect 213802 -3514 213946 -3277
rect 214132 -3299 214518 -3277
rect 214056 -3385 214518 -3299
rect 214060 -3393 214260 -3385
rect 214076 -3397 214244 -3393
rect 213802 -3600 213976 -3514
rect 214002 -3574 214102 -3450
rect 214002 -3628 214004 -3574
rect 213687 -4371 213831 -4324
rect 213868 -4371 213885 -4270
rect 213687 -4382 214459 -4371
rect 213773 -4407 214459 -4382
rect 213785 -4436 214459 -4407
rect 213785 -4848 214518 -4436
rect 214967 -4848 215014 -4483
rect 215021 -4848 215068 -4537
rect 213785 -4906 215139 -4848
rect 213212 -4943 215139 -4906
rect 213212 -5067 215641 -4943
rect 213212 -6022 215694 -5067
rect 216556 -6022 217020 -4906
rect 213803 -6087 215694 -6022
rect 214394 -6147 215694 -6087
rect 214423 -6152 215694 -6147
rect 214547 -6170 215694 -6152
rect 214985 -6181 215694 -6170
rect 214985 -6217 215659 -6181
rect 215168 -6235 215659 -6217
<< error_ps >>
rect 217146 -3514 217290 -3274
rect 217476 -3299 217862 -3153
rect 217400 -3385 217862 -3299
rect 217146 -3600 217320 -3514
rect 2540 -6022 2720 -4906
rect 211496 -4943 211795 -4848
rect 217147 -4436 217803 -4371
rect 217147 -4848 217862 -4436
rect 217147 -4906 218280 -4848
rect 211496 -6152 212297 -4943
rect 211641 -6217 212297 -6152
rect 217020 -6022 218280 -4906
rect 217147 -6087 218280 -6022
rect 217738 -6147 218280 -6087
rect 217767 -6152 218280 -6147
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use icell64scs  x1
timestamp 1717439242
transform 1 0 0 0 1 0
box 0 -6337 215760 458
use icell64scs  x2
timestamp 1717439242
transform 1 0 214016 0 1 0
box 0 -6337 215760 458
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
