magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< nwell >>
rect -358 -183987 358 183987
<< mvpmos >>
rect -100 182490 100 183690
rect -100 181054 100 182254
rect -100 179618 100 180818
rect -100 178182 100 179382
rect -100 176746 100 177946
rect -100 175310 100 176510
rect -100 173874 100 175074
rect -100 172438 100 173638
rect -100 171002 100 172202
rect -100 169566 100 170766
rect -100 168130 100 169330
rect -100 166694 100 167894
rect -100 165258 100 166458
rect -100 163822 100 165022
rect -100 162386 100 163586
rect -100 160950 100 162150
rect -100 159514 100 160714
rect -100 158078 100 159278
rect -100 156642 100 157842
rect -100 155206 100 156406
rect -100 153770 100 154970
rect -100 152334 100 153534
rect -100 150898 100 152098
rect -100 149462 100 150662
rect -100 148026 100 149226
rect -100 146590 100 147790
rect -100 145154 100 146354
rect -100 143718 100 144918
rect -100 142282 100 143482
rect -100 140846 100 142046
rect -100 139410 100 140610
rect -100 137974 100 139174
rect -100 136538 100 137738
rect -100 135102 100 136302
rect -100 133666 100 134866
rect -100 132230 100 133430
rect -100 130794 100 131994
rect -100 129358 100 130558
rect -100 127922 100 129122
rect -100 126486 100 127686
rect -100 125050 100 126250
rect -100 123614 100 124814
rect -100 122178 100 123378
rect -100 120742 100 121942
rect -100 119306 100 120506
rect -100 117870 100 119070
rect -100 116434 100 117634
rect -100 114998 100 116198
rect -100 113562 100 114762
rect -100 112126 100 113326
rect -100 110690 100 111890
rect -100 109254 100 110454
rect -100 107818 100 109018
rect -100 106382 100 107582
rect -100 104946 100 106146
rect -100 103510 100 104710
rect -100 102074 100 103274
rect -100 100638 100 101838
rect -100 99202 100 100402
rect -100 97766 100 98966
rect -100 96330 100 97530
rect -100 94894 100 96094
rect -100 93458 100 94658
rect -100 92022 100 93222
rect -100 90586 100 91786
rect -100 89150 100 90350
rect -100 87714 100 88914
rect -100 86278 100 87478
rect -100 84842 100 86042
rect -100 83406 100 84606
rect -100 81970 100 83170
rect -100 80534 100 81734
rect -100 79098 100 80298
rect -100 77662 100 78862
rect -100 76226 100 77426
rect -100 74790 100 75990
rect -100 73354 100 74554
rect -100 71918 100 73118
rect -100 70482 100 71682
rect -100 69046 100 70246
rect -100 67610 100 68810
rect -100 66174 100 67374
rect -100 64738 100 65938
rect -100 63302 100 64502
rect -100 61866 100 63066
rect -100 60430 100 61630
rect -100 58994 100 60194
rect -100 57558 100 58758
rect -100 56122 100 57322
rect -100 54686 100 55886
rect -100 53250 100 54450
rect -100 51814 100 53014
rect -100 50378 100 51578
rect -100 48942 100 50142
rect -100 47506 100 48706
rect -100 46070 100 47270
rect -100 44634 100 45834
rect -100 43198 100 44398
rect -100 41762 100 42962
rect -100 40326 100 41526
rect -100 38890 100 40090
rect -100 37454 100 38654
rect -100 36018 100 37218
rect -100 34582 100 35782
rect -100 33146 100 34346
rect -100 31710 100 32910
rect -100 30274 100 31474
rect -100 28838 100 30038
rect -100 27402 100 28602
rect -100 25966 100 27166
rect -100 24530 100 25730
rect -100 23094 100 24294
rect -100 21658 100 22858
rect -100 20222 100 21422
rect -100 18786 100 19986
rect -100 17350 100 18550
rect -100 15914 100 17114
rect -100 14478 100 15678
rect -100 13042 100 14242
rect -100 11606 100 12806
rect -100 10170 100 11370
rect -100 8734 100 9934
rect -100 7298 100 8498
rect -100 5862 100 7062
rect -100 4426 100 5626
rect -100 2990 100 4190
rect -100 1554 100 2754
rect -100 118 100 1318
rect -100 -1318 100 -118
rect -100 -2754 100 -1554
rect -100 -4190 100 -2990
rect -100 -5626 100 -4426
rect -100 -7062 100 -5862
rect -100 -8498 100 -7298
rect -100 -9934 100 -8734
rect -100 -11370 100 -10170
rect -100 -12806 100 -11606
rect -100 -14242 100 -13042
rect -100 -15678 100 -14478
rect -100 -17114 100 -15914
rect -100 -18550 100 -17350
rect -100 -19986 100 -18786
rect -100 -21422 100 -20222
rect -100 -22858 100 -21658
rect -100 -24294 100 -23094
rect -100 -25730 100 -24530
rect -100 -27166 100 -25966
rect -100 -28602 100 -27402
rect -100 -30038 100 -28838
rect -100 -31474 100 -30274
rect -100 -32910 100 -31710
rect -100 -34346 100 -33146
rect -100 -35782 100 -34582
rect -100 -37218 100 -36018
rect -100 -38654 100 -37454
rect -100 -40090 100 -38890
rect -100 -41526 100 -40326
rect -100 -42962 100 -41762
rect -100 -44398 100 -43198
rect -100 -45834 100 -44634
rect -100 -47270 100 -46070
rect -100 -48706 100 -47506
rect -100 -50142 100 -48942
rect -100 -51578 100 -50378
rect -100 -53014 100 -51814
rect -100 -54450 100 -53250
rect -100 -55886 100 -54686
rect -100 -57322 100 -56122
rect -100 -58758 100 -57558
rect -100 -60194 100 -58994
rect -100 -61630 100 -60430
rect -100 -63066 100 -61866
rect -100 -64502 100 -63302
rect -100 -65938 100 -64738
rect -100 -67374 100 -66174
rect -100 -68810 100 -67610
rect -100 -70246 100 -69046
rect -100 -71682 100 -70482
rect -100 -73118 100 -71918
rect -100 -74554 100 -73354
rect -100 -75990 100 -74790
rect -100 -77426 100 -76226
rect -100 -78862 100 -77662
rect -100 -80298 100 -79098
rect -100 -81734 100 -80534
rect -100 -83170 100 -81970
rect -100 -84606 100 -83406
rect -100 -86042 100 -84842
rect -100 -87478 100 -86278
rect -100 -88914 100 -87714
rect -100 -90350 100 -89150
rect -100 -91786 100 -90586
rect -100 -93222 100 -92022
rect -100 -94658 100 -93458
rect -100 -96094 100 -94894
rect -100 -97530 100 -96330
rect -100 -98966 100 -97766
rect -100 -100402 100 -99202
rect -100 -101838 100 -100638
rect -100 -103274 100 -102074
rect -100 -104710 100 -103510
rect -100 -106146 100 -104946
rect -100 -107582 100 -106382
rect -100 -109018 100 -107818
rect -100 -110454 100 -109254
rect -100 -111890 100 -110690
rect -100 -113326 100 -112126
rect -100 -114762 100 -113562
rect -100 -116198 100 -114998
rect -100 -117634 100 -116434
rect -100 -119070 100 -117870
rect -100 -120506 100 -119306
rect -100 -121942 100 -120742
rect -100 -123378 100 -122178
rect -100 -124814 100 -123614
rect -100 -126250 100 -125050
rect -100 -127686 100 -126486
rect -100 -129122 100 -127922
rect -100 -130558 100 -129358
rect -100 -131994 100 -130794
rect -100 -133430 100 -132230
rect -100 -134866 100 -133666
rect -100 -136302 100 -135102
rect -100 -137738 100 -136538
rect -100 -139174 100 -137974
rect -100 -140610 100 -139410
rect -100 -142046 100 -140846
rect -100 -143482 100 -142282
rect -100 -144918 100 -143718
rect -100 -146354 100 -145154
rect -100 -147790 100 -146590
rect -100 -149226 100 -148026
rect -100 -150662 100 -149462
rect -100 -152098 100 -150898
rect -100 -153534 100 -152334
rect -100 -154970 100 -153770
rect -100 -156406 100 -155206
rect -100 -157842 100 -156642
rect -100 -159278 100 -158078
rect -100 -160714 100 -159514
rect -100 -162150 100 -160950
rect -100 -163586 100 -162386
rect -100 -165022 100 -163822
rect -100 -166458 100 -165258
rect -100 -167894 100 -166694
rect -100 -169330 100 -168130
rect -100 -170766 100 -169566
rect -100 -172202 100 -171002
rect -100 -173638 100 -172438
rect -100 -175074 100 -173874
rect -100 -176510 100 -175310
rect -100 -177946 100 -176746
rect -100 -179382 100 -178182
rect -100 -180818 100 -179618
rect -100 -182254 100 -181054
rect -100 -183690 100 -182490
<< mvpdiff >>
rect -158 183678 -100 183690
rect -158 182502 -146 183678
rect -112 182502 -100 183678
rect -158 182490 -100 182502
rect 100 183678 158 183690
rect 100 182502 112 183678
rect 146 182502 158 183678
rect 100 182490 158 182502
rect -158 182242 -100 182254
rect -158 181066 -146 182242
rect -112 181066 -100 182242
rect -158 181054 -100 181066
rect 100 182242 158 182254
rect 100 181066 112 182242
rect 146 181066 158 182242
rect 100 181054 158 181066
rect -158 180806 -100 180818
rect -158 179630 -146 180806
rect -112 179630 -100 180806
rect -158 179618 -100 179630
rect 100 180806 158 180818
rect 100 179630 112 180806
rect 146 179630 158 180806
rect 100 179618 158 179630
rect -158 179370 -100 179382
rect -158 178194 -146 179370
rect -112 178194 -100 179370
rect -158 178182 -100 178194
rect 100 179370 158 179382
rect 100 178194 112 179370
rect 146 178194 158 179370
rect 100 178182 158 178194
rect -158 177934 -100 177946
rect -158 176758 -146 177934
rect -112 176758 -100 177934
rect -158 176746 -100 176758
rect 100 177934 158 177946
rect 100 176758 112 177934
rect 146 176758 158 177934
rect 100 176746 158 176758
rect -158 176498 -100 176510
rect -158 175322 -146 176498
rect -112 175322 -100 176498
rect -158 175310 -100 175322
rect 100 176498 158 176510
rect 100 175322 112 176498
rect 146 175322 158 176498
rect 100 175310 158 175322
rect -158 175062 -100 175074
rect -158 173886 -146 175062
rect -112 173886 -100 175062
rect -158 173874 -100 173886
rect 100 175062 158 175074
rect 100 173886 112 175062
rect 146 173886 158 175062
rect 100 173874 158 173886
rect -158 173626 -100 173638
rect -158 172450 -146 173626
rect -112 172450 -100 173626
rect -158 172438 -100 172450
rect 100 173626 158 173638
rect 100 172450 112 173626
rect 146 172450 158 173626
rect 100 172438 158 172450
rect -158 172190 -100 172202
rect -158 171014 -146 172190
rect -112 171014 -100 172190
rect -158 171002 -100 171014
rect 100 172190 158 172202
rect 100 171014 112 172190
rect 146 171014 158 172190
rect 100 171002 158 171014
rect -158 170754 -100 170766
rect -158 169578 -146 170754
rect -112 169578 -100 170754
rect -158 169566 -100 169578
rect 100 170754 158 170766
rect 100 169578 112 170754
rect 146 169578 158 170754
rect 100 169566 158 169578
rect -158 169318 -100 169330
rect -158 168142 -146 169318
rect -112 168142 -100 169318
rect -158 168130 -100 168142
rect 100 169318 158 169330
rect 100 168142 112 169318
rect 146 168142 158 169318
rect 100 168130 158 168142
rect -158 167882 -100 167894
rect -158 166706 -146 167882
rect -112 166706 -100 167882
rect -158 166694 -100 166706
rect 100 167882 158 167894
rect 100 166706 112 167882
rect 146 166706 158 167882
rect 100 166694 158 166706
rect -158 166446 -100 166458
rect -158 165270 -146 166446
rect -112 165270 -100 166446
rect -158 165258 -100 165270
rect 100 166446 158 166458
rect 100 165270 112 166446
rect 146 165270 158 166446
rect 100 165258 158 165270
rect -158 165010 -100 165022
rect -158 163834 -146 165010
rect -112 163834 -100 165010
rect -158 163822 -100 163834
rect 100 165010 158 165022
rect 100 163834 112 165010
rect 146 163834 158 165010
rect 100 163822 158 163834
rect -158 163574 -100 163586
rect -158 162398 -146 163574
rect -112 162398 -100 163574
rect -158 162386 -100 162398
rect 100 163574 158 163586
rect 100 162398 112 163574
rect 146 162398 158 163574
rect 100 162386 158 162398
rect -158 162138 -100 162150
rect -158 160962 -146 162138
rect -112 160962 -100 162138
rect -158 160950 -100 160962
rect 100 162138 158 162150
rect 100 160962 112 162138
rect 146 160962 158 162138
rect 100 160950 158 160962
rect -158 160702 -100 160714
rect -158 159526 -146 160702
rect -112 159526 -100 160702
rect -158 159514 -100 159526
rect 100 160702 158 160714
rect 100 159526 112 160702
rect 146 159526 158 160702
rect 100 159514 158 159526
rect -158 159266 -100 159278
rect -158 158090 -146 159266
rect -112 158090 -100 159266
rect -158 158078 -100 158090
rect 100 159266 158 159278
rect 100 158090 112 159266
rect 146 158090 158 159266
rect 100 158078 158 158090
rect -158 157830 -100 157842
rect -158 156654 -146 157830
rect -112 156654 -100 157830
rect -158 156642 -100 156654
rect 100 157830 158 157842
rect 100 156654 112 157830
rect 146 156654 158 157830
rect 100 156642 158 156654
rect -158 156394 -100 156406
rect -158 155218 -146 156394
rect -112 155218 -100 156394
rect -158 155206 -100 155218
rect 100 156394 158 156406
rect 100 155218 112 156394
rect 146 155218 158 156394
rect 100 155206 158 155218
rect -158 154958 -100 154970
rect -158 153782 -146 154958
rect -112 153782 -100 154958
rect -158 153770 -100 153782
rect 100 154958 158 154970
rect 100 153782 112 154958
rect 146 153782 158 154958
rect 100 153770 158 153782
rect -158 153522 -100 153534
rect -158 152346 -146 153522
rect -112 152346 -100 153522
rect -158 152334 -100 152346
rect 100 153522 158 153534
rect 100 152346 112 153522
rect 146 152346 158 153522
rect 100 152334 158 152346
rect -158 152086 -100 152098
rect -158 150910 -146 152086
rect -112 150910 -100 152086
rect -158 150898 -100 150910
rect 100 152086 158 152098
rect 100 150910 112 152086
rect 146 150910 158 152086
rect 100 150898 158 150910
rect -158 150650 -100 150662
rect -158 149474 -146 150650
rect -112 149474 -100 150650
rect -158 149462 -100 149474
rect 100 150650 158 150662
rect 100 149474 112 150650
rect 146 149474 158 150650
rect 100 149462 158 149474
rect -158 149214 -100 149226
rect -158 148038 -146 149214
rect -112 148038 -100 149214
rect -158 148026 -100 148038
rect 100 149214 158 149226
rect 100 148038 112 149214
rect 146 148038 158 149214
rect 100 148026 158 148038
rect -158 147778 -100 147790
rect -158 146602 -146 147778
rect -112 146602 -100 147778
rect -158 146590 -100 146602
rect 100 147778 158 147790
rect 100 146602 112 147778
rect 146 146602 158 147778
rect 100 146590 158 146602
rect -158 146342 -100 146354
rect -158 145166 -146 146342
rect -112 145166 -100 146342
rect -158 145154 -100 145166
rect 100 146342 158 146354
rect 100 145166 112 146342
rect 146 145166 158 146342
rect 100 145154 158 145166
rect -158 144906 -100 144918
rect -158 143730 -146 144906
rect -112 143730 -100 144906
rect -158 143718 -100 143730
rect 100 144906 158 144918
rect 100 143730 112 144906
rect 146 143730 158 144906
rect 100 143718 158 143730
rect -158 143470 -100 143482
rect -158 142294 -146 143470
rect -112 142294 -100 143470
rect -158 142282 -100 142294
rect 100 143470 158 143482
rect 100 142294 112 143470
rect 146 142294 158 143470
rect 100 142282 158 142294
rect -158 142034 -100 142046
rect -158 140858 -146 142034
rect -112 140858 -100 142034
rect -158 140846 -100 140858
rect 100 142034 158 142046
rect 100 140858 112 142034
rect 146 140858 158 142034
rect 100 140846 158 140858
rect -158 140598 -100 140610
rect -158 139422 -146 140598
rect -112 139422 -100 140598
rect -158 139410 -100 139422
rect 100 140598 158 140610
rect 100 139422 112 140598
rect 146 139422 158 140598
rect 100 139410 158 139422
rect -158 139162 -100 139174
rect -158 137986 -146 139162
rect -112 137986 -100 139162
rect -158 137974 -100 137986
rect 100 139162 158 139174
rect 100 137986 112 139162
rect 146 137986 158 139162
rect 100 137974 158 137986
rect -158 137726 -100 137738
rect -158 136550 -146 137726
rect -112 136550 -100 137726
rect -158 136538 -100 136550
rect 100 137726 158 137738
rect 100 136550 112 137726
rect 146 136550 158 137726
rect 100 136538 158 136550
rect -158 136290 -100 136302
rect -158 135114 -146 136290
rect -112 135114 -100 136290
rect -158 135102 -100 135114
rect 100 136290 158 136302
rect 100 135114 112 136290
rect 146 135114 158 136290
rect 100 135102 158 135114
rect -158 134854 -100 134866
rect -158 133678 -146 134854
rect -112 133678 -100 134854
rect -158 133666 -100 133678
rect 100 134854 158 134866
rect 100 133678 112 134854
rect 146 133678 158 134854
rect 100 133666 158 133678
rect -158 133418 -100 133430
rect -158 132242 -146 133418
rect -112 132242 -100 133418
rect -158 132230 -100 132242
rect 100 133418 158 133430
rect 100 132242 112 133418
rect 146 132242 158 133418
rect 100 132230 158 132242
rect -158 131982 -100 131994
rect -158 130806 -146 131982
rect -112 130806 -100 131982
rect -158 130794 -100 130806
rect 100 131982 158 131994
rect 100 130806 112 131982
rect 146 130806 158 131982
rect 100 130794 158 130806
rect -158 130546 -100 130558
rect -158 129370 -146 130546
rect -112 129370 -100 130546
rect -158 129358 -100 129370
rect 100 130546 158 130558
rect 100 129370 112 130546
rect 146 129370 158 130546
rect 100 129358 158 129370
rect -158 129110 -100 129122
rect -158 127934 -146 129110
rect -112 127934 -100 129110
rect -158 127922 -100 127934
rect 100 129110 158 129122
rect 100 127934 112 129110
rect 146 127934 158 129110
rect 100 127922 158 127934
rect -158 127674 -100 127686
rect -158 126498 -146 127674
rect -112 126498 -100 127674
rect -158 126486 -100 126498
rect 100 127674 158 127686
rect 100 126498 112 127674
rect 146 126498 158 127674
rect 100 126486 158 126498
rect -158 126238 -100 126250
rect -158 125062 -146 126238
rect -112 125062 -100 126238
rect -158 125050 -100 125062
rect 100 126238 158 126250
rect 100 125062 112 126238
rect 146 125062 158 126238
rect 100 125050 158 125062
rect -158 124802 -100 124814
rect -158 123626 -146 124802
rect -112 123626 -100 124802
rect -158 123614 -100 123626
rect 100 124802 158 124814
rect 100 123626 112 124802
rect 146 123626 158 124802
rect 100 123614 158 123626
rect -158 123366 -100 123378
rect -158 122190 -146 123366
rect -112 122190 -100 123366
rect -158 122178 -100 122190
rect 100 123366 158 123378
rect 100 122190 112 123366
rect 146 122190 158 123366
rect 100 122178 158 122190
rect -158 121930 -100 121942
rect -158 120754 -146 121930
rect -112 120754 -100 121930
rect -158 120742 -100 120754
rect 100 121930 158 121942
rect 100 120754 112 121930
rect 146 120754 158 121930
rect 100 120742 158 120754
rect -158 120494 -100 120506
rect -158 119318 -146 120494
rect -112 119318 -100 120494
rect -158 119306 -100 119318
rect 100 120494 158 120506
rect 100 119318 112 120494
rect 146 119318 158 120494
rect 100 119306 158 119318
rect -158 119058 -100 119070
rect -158 117882 -146 119058
rect -112 117882 -100 119058
rect -158 117870 -100 117882
rect 100 119058 158 119070
rect 100 117882 112 119058
rect 146 117882 158 119058
rect 100 117870 158 117882
rect -158 117622 -100 117634
rect -158 116446 -146 117622
rect -112 116446 -100 117622
rect -158 116434 -100 116446
rect 100 117622 158 117634
rect 100 116446 112 117622
rect 146 116446 158 117622
rect 100 116434 158 116446
rect -158 116186 -100 116198
rect -158 115010 -146 116186
rect -112 115010 -100 116186
rect -158 114998 -100 115010
rect 100 116186 158 116198
rect 100 115010 112 116186
rect 146 115010 158 116186
rect 100 114998 158 115010
rect -158 114750 -100 114762
rect -158 113574 -146 114750
rect -112 113574 -100 114750
rect -158 113562 -100 113574
rect 100 114750 158 114762
rect 100 113574 112 114750
rect 146 113574 158 114750
rect 100 113562 158 113574
rect -158 113314 -100 113326
rect -158 112138 -146 113314
rect -112 112138 -100 113314
rect -158 112126 -100 112138
rect 100 113314 158 113326
rect 100 112138 112 113314
rect 146 112138 158 113314
rect 100 112126 158 112138
rect -158 111878 -100 111890
rect -158 110702 -146 111878
rect -112 110702 -100 111878
rect -158 110690 -100 110702
rect 100 111878 158 111890
rect 100 110702 112 111878
rect 146 110702 158 111878
rect 100 110690 158 110702
rect -158 110442 -100 110454
rect -158 109266 -146 110442
rect -112 109266 -100 110442
rect -158 109254 -100 109266
rect 100 110442 158 110454
rect 100 109266 112 110442
rect 146 109266 158 110442
rect 100 109254 158 109266
rect -158 109006 -100 109018
rect -158 107830 -146 109006
rect -112 107830 -100 109006
rect -158 107818 -100 107830
rect 100 109006 158 109018
rect 100 107830 112 109006
rect 146 107830 158 109006
rect 100 107818 158 107830
rect -158 107570 -100 107582
rect -158 106394 -146 107570
rect -112 106394 -100 107570
rect -158 106382 -100 106394
rect 100 107570 158 107582
rect 100 106394 112 107570
rect 146 106394 158 107570
rect 100 106382 158 106394
rect -158 106134 -100 106146
rect -158 104958 -146 106134
rect -112 104958 -100 106134
rect -158 104946 -100 104958
rect 100 106134 158 106146
rect 100 104958 112 106134
rect 146 104958 158 106134
rect 100 104946 158 104958
rect -158 104698 -100 104710
rect -158 103522 -146 104698
rect -112 103522 -100 104698
rect -158 103510 -100 103522
rect 100 104698 158 104710
rect 100 103522 112 104698
rect 146 103522 158 104698
rect 100 103510 158 103522
rect -158 103262 -100 103274
rect -158 102086 -146 103262
rect -112 102086 -100 103262
rect -158 102074 -100 102086
rect 100 103262 158 103274
rect 100 102086 112 103262
rect 146 102086 158 103262
rect 100 102074 158 102086
rect -158 101826 -100 101838
rect -158 100650 -146 101826
rect -112 100650 -100 101826
rect -158 100638 -100 100650
rect 100 101826 158 101838
rect 100 100650 112 101826
rect 146 100650 158 101826
rect 100 100638 158 100650
rect -158 100390 -100 100402
rect -158 99214 -146 100390
rect -112 99214 -100 100390
rect -158 99202 -100 99214
rect 100 100390 158 100402
rect 100 99214 112 100390
rect 146 99214 158 100390
rect 100 99202 158 99214
rect -158 98954 -100 98966
rect -158 97778 -146 98954
rect -112 97778 -100 98954
rect -158 97766 -100 97778
rect 100 98954 158 98966
rect 100 97778 112 98954
rect 146 97778 158 98954
rect 100 97766 158 97778
rect -158 97518 -100 97530
rect -158 96342 -146 97518
rect -112 96342 -100 97518
rect -158 96330 -100 96342
rect 100 97518 158 97530
rect 100 96342 112 97518
rect 146 96342 158 97518
rect 100 96330 158 96342
rect -158 96082 -100 96094
rect -158 94906 -146 96082
rect -112 94906 -100 96082
rect -158 94894 -100 94906
rect 100 96082 158 96094
rect 100 94906 112 96082
rect 146 94906 158 96082
rect 100 94894 158 94906
rect -158 94646 -100 94658
rect -158 93470 -146 94646
rect -112 93470 -100 94646
rect -158 93458 -100 93470
rect 100 94646 158 94658
rect 100 93470 112 94646
rect 146 93470 158 94646
rect 100 93458 158 93470
rect -158 93210 -100 93222
rect -158 92034 -146 93210
rect -112 92034 -100 93210
rect -158 92022 -100 92034
rect 100 93210 158 93222
rect 100 92034 112 93210
rect 146 92034 158 93210
rect 100 92022 158 92034
rect -158 91774 -100 91786
rect -158 90598 -146 91774
rect -112 90598 -100 91774
rect -158 90586 -100 90598
rect 100 91774 158 91786
rect 100 90598 112 91774
rect 146 90598 158 91774
rect 100 90586 158 90598
rect -158 90338 -100 90350
rect -158 89162 -146 90338
rect -112 89162 -100 90338
rect -158 89150 -100 89162
rect 100 90338 158 90350
rect 100 89162 112 90338
rect 146 89162 158 90338
rect 100 89150 158 89162
rect -158 88902 -100 88914
rect -158 87726 -146 88902
rect -112 87726 -100 88902
rect -158 87714 -100 87726
rect 100 88902 158 88914
rect 100 87726 112 88902
rect 146 87726 158 88902
rect 100 87714 158 87726
rect -158 87466 -100 87478
rect -158 86290 -146 87466
rect -112 86290 -100 87466
rect -158 86278 -100 86290
rect 100 87466 158 87478
rect 100 86290 112 87466
rect 146 86290 158 87466
rect 100 86278 158 86290
rect -158 86030 -100 86042
rect -158 84854 -146 86030
rect -112 84854 -100 86030
rect -158 84842 -100 84854
rect 100 86030 158 86042
rect 100 84854 112 86030
rect 146 84854 158 86030
rect 100 84842 158 84854
rect -158 84594 -100 84606
rect -158 83418 -146 84594
rect -112 83418 -100 84594
rect -158 83406 -100 83418
rect 100 84594 158 84606
rect 100 83418 112 84594
rect 146 83418 158 84594
rect 100 83406 158 83418
rect -158 83158 -100 83170
rect -158 81982 -146 83158
rect -112 81982 -100 83158
rect -158 81970 -100 81982
rect 100 83158 158 83170
rect 100 81982 112 83158
rect 146 81982 158 83158
rect 100 81970 158 81982
rect -158 81722 -100 81734
rect -158 80546 -146 81722
rect -112 80546 -100 81722
rect -158 80534 -100 80546
rect 100 81722 158 81734
rect 100 80546 112 81722
rect 146 80546 158 81722
rect 100 80534 158 80546
rect -158 80286 -100 80298
rect -158 79110 -146 80286
rect -112 79110 -100 80286
rect -158 79098 -100 79110
rect 100 80286 158 80298
rect 100 79110 112 80286
rect 146 79110 158 80286
rect 100 79098 158 79110
rect -158 78850 -100 78862
rect -158 77674 -146 78850
rect -112 77674 -100 78850
rect -158 77662 -100 77674
rect 100 78850 158 78862
rect 100 77674 112 78850
rect 146 77674 158 78850
rect 100 77662 158 77674
rect -158 77414 -100 77426
rect -158 76238 -146 77414
rect -112 76238 -100 77414
rect -158 76226 -100 76238
rect 100 77414 158 77426
rect 100 76238 112 77414
rect 146 76238 158 77414
rect 100 76226 158 76238
rect -158 75978 -100 75990
rect -158 74802 -146 75978
rect -112 74802 -100 75978
rect -158 74790 -100 74802
rect 100 75978 158 75990
rect 100 74802 112 75978
rect 146 74802 158 75978
rect 100 74790 158 74802
rect -158 74542 -100 74554
rect -158 73366 -146 74542
rect -112 73366 -100 74542
rect -158 73354 -100 73366
rect 100 74542 158 74554
rect 100 73366 112 74542
rect 146 73366 158 74542
rect 100 73354 158 73366
rect -158 73106 -100 73118
rect -158 71930 -146 73106
rect -112 71930 -100 73106
rect -158 71918 -100 71930
rect 100 73106 158 73118
rect 100 71930 112 73106
rect 146 71930 158 73106
rect 100 71918 158 71930
rect -158 71670 -100 71682
rect -158 70494 -146 71670
rect -112 70494 -100 71670
rect -158 70482 -100 70494
rect 100 71670 158 71682
rect 100 70494 112 71670
rect 146 70494 158 71670
rect 100 70482 158 70494
rect -158 70234 -100 70246
rect -158 69058 -146 70234
rect -112 69058 -100 70234
rect -158 69046 -100 69058
rect 100 70234 158 70246
rect 100 69058 112 70234
rect 146 69058 158 70234
rect 100 69046 158 69058
rect -158 68798 -100 68810
rect -158 67622 -146 68798
rect -112 67622 -100 68798
rect -158 67610 -100 67622
rect 100 68798 158 68810
rect 100 67622 112 68798
rect 146 67622 158 68798
rect 100 67610 158 67622
rect -158 67362 -100 67374
rect -158 66186 -146 67362
rect -112 66186 -100 67362
rect -158 66174 -100 66186
rect 100 67362 158 67374
rect 100 66186 112 67362
rect 146 66186 158 67362
rect 100 66174 158 66186
rect -158 65926 -100 65938
rect -158 64750 -146 65926
rect -112 64750 -100 65926
rect -158 64738 -100 64750
rect 100 65926 158 65938
rect 100 64750 112 65926
rect 146 64750 158 65926
rect 100 64738 158 64750
rect -158 64490 -100 64502
rect -158 63314 -146 64490
rect -112 63314 -100 64490
rect -158 63302 -100 63314
rect 100 64490 158 64502
rect 100 63314 112 64490
rect 146 63314 158 64490
rect 100 63302 158 63314
rect -158 63054 -100 63066
rect -158 61878 -146 63054
rect -112 61878 -100 63054
rect -158 61866 -100 61878
rect 100 63054 158 63066
rect 100 61878 112 63054
rect 146 61878 158 63054
rect 100 61866 158 61878
rect -158 61618 -100 61630
rect -158 60442 -146 61618
rect -112 60442 -100 61618
rect -158 60430 -100 60442
rect 100 61618 158 61630
rect 100 60442 112 61618
rect 146 60442 158 61618
rect 100 60430 158 60442
rect -158 60182 -100 60194
rect -158 59006 -146 60182
rect -112 59006 -100 60182
rect -158 58994 -100 59006
rect 100 60182 158 60194
rect 100 59006 112 60182
rect 146 59006 158 60182
rect 100 58994 158 59006
rect -158 58746 -100 58758
rect -158 57570 -146 58746
rect -112 57570 -100 58746
rect -158 57558 -100 57570
rect 100 58746 158 58758
rect 100 57570 112 58746
rect 146 57570 158 58746
rect 100 57558 158 57570
rect -158 57310 -100 57322
rect -158 56134 -146 57310
rect -112 56134 -100 57310
rect -158 56122 -100 56134
rect 100 57310 158 57322
rect 100 56134 112 57310
rect 146 56134 158 57310
rect 100 56122 158 56134
rect -158 55874 -100 55886
rect -158 54698 -146 55874
rect -112 54698 -100 55874
rect -158 54686 -100 54698
rect 100 55874 158 55886
rect 100 54698 112 55874
rect 146 54698 158 55874
rect 100 54686 158 54698
rect -158 54438 -100 54450
rect -158 53262 -146 54438
rect -112 53262 -100 54438
rect -158 53250 -100 53262
rect 100 54438 158 54450
rect 100 53262 112 54438
rect 146 53262 158 54438
rect 100 53250 158 53262
rect -158 53002 -100 53014
rect -158 51826 -146 53002
rect -112 51826 -100 53002
rect -158 51814 -100 51826
rect 100 53002 158 53014
rect 100 51826 112 53002
rect 146 51826 158 53002
rect 100 51814 158 51826
rect -158 51566 -100 51578
rect -158 50390 -146 51566
rect -112 50390 -100 51566
rect -158 50378 -100 50390
rect 100 51566 158 51578
rect 100 50390 112 51566
rect 146 50390 158 51566
rect 100 50378 158 50390
rect -158 50130 -100 50142
rect -158 48954 -146 50130
rect -112 48954 -100 50130
rect -158 48942 -100 48954
rect 100 50130 158 50142
rect 100 48954 112 50130
rect 146 48954 158 50130
rect 100 48942 158 48954
rect -158 48694 -100 48706
rect -158 47518 -146 48694
rect -112 47518 -100 48694
rect -158 47506 -100 47518
rect 100 48694 158 48706
rect 100 47518 112 48694
rect 146 47518 158 48694
rect 100 47506 158 47518
rect -158 47258 -100 47270
rect -158 46082 -146 47258
rect -112 46082 -100 47258
rect -158 46070 -100 46082
rect 100 47258 158 47270
rect 100 46082 112 47258
rect 146 46082 158 47258
rect 100 46070 158 46082
rect -158 45822 -100 45834
rect -158 44646 -146 45822
rect -112 44646 -100 45822
rect -158 44634 -100 44646
rect 100 45822 158 45834
rect 100 44646 112 45822
rect 146 44646 158 45822
rect 100 44634 158 44646
rect -158 44386 -100 44398
rect -158 43210 -146 44386
rect -112 43210 -100 44386
rect -158 43198 -100 43210
rect 100 44386 158 44398
rect 100 43210 112 44386
rect 146 43210 158 44386
rect 100 43198 158 43210
rect -158 42950 -100 42962
rect -158 41774 -146 42950
rect -112 41774 -100 42950
rect -158 41762 -100 41774
rect 100 42950 158 42962
rect 100 41774 112 42950
rect 146 41774 158 42950
rect 100 41762 158 41774
rect -158 41514 -100 41526
rect -158 40338 -146 41514
rect -112 40338 -100 41514
rect -158 40326 -100 40338
rect 100 41514 158 41526
rect 100 40338 112 41514
rect 146 40338 158 41514
rect 100 40326 158 40338
rect -158 40078 -100 40090
rect -158 38902 -146 40078
rect -112 38902 -100 40078
rect -158 38890 -100 38902
rect 100 40078 158 40090
rect 100 38902 112 40078
rect 146 38902 158 40078
rect 100 38890 158 38902
rect -158 38642 -100 38654
rect -158 37466 -146 38642
rect -112 37466 -100 38642
rect -158 37454 -100 37466
rect 100 38642 158 38654
rect 100 37466 112 38642
rect 146 37466 158 38642
rect 100 37454 158 37466
rect -158 37206 -100 37218
rect -158 36030 -146 37206
rect -112 36030 -100 37206
rect -158 36018 -100 36030
rect 100 37206 158 37218
rect 100 36030 112 37206
rect 146 36030 158 37206
rect 100 36018 158 36030
rect -158 35770 -100 35782
rect -158 34594 -146 35770
rect -112 34594 -100 35770
rect -158 34582 -100 34594
rect 100 35770 158 35782
rect 100 34594 112 35770
rect 146 34594 158 35770
rect 100 34582 158 34594
rect -158 34334 -100 34346
rect -158 33158 -146 34334
rect -112 33158 -100 34334
rect -158 33146 -100 33158
rect 100 34334 158 34346
rect 100 33158 112 34334
rect 146 33158 158 34334
rect 100 33146 158 33158
rect -158 32898 -100 32910
rect -158 31722 -146 32898
rect -112 31722 -100 32898
rect -158 31710 -100 31722
rect 100 32898 158 32910
rect 100 31722 112 32898
rect 146 31722 158 32898
rect 100 31710 158 31722
rect -158 31462 -100 31474
rect -158 30286 -146 31462
rect -112 30286 -100 31462
rect -158 30274 -100 30286
rect 100 31462 158 31474
rect 100 30286 112 31462
rect 146 30286 158 31462
rect 100 30274 158 30286
rect -158 30026 -100 30038
rect -158 28850 -146 30026
rect -112 28850 -100 30026
rect -158 28838 -100 28850
rect 100 30026 158 30038
rect 100 28850 112 30026
rect 146 28850 158 30026
rect 100 28838 158 28850
rect -158 28590 -100 28602
rect -158 27414 -146 28590
rect -112 27414 -100 28590
rect -158 27402 -100 27414
rect 100 28590 158 28602
rect 100 27414 112 28590
rect 146 27414 158 28590
rect 100 27402 158 27414
rect -158 27154 -100 27166
rect -158 25978 -146 27154
rect -112 25978 -100 27154
rect -158 25966 -100 25978
rect 100 27154 158 27166
rect 100 25978 112 27154
rect 146 25978 158 27154
rect 100 25966 158 25978
rect -158 25718 -100 25730
rect -158 24542 -146 25718
rect -112 24542 -100 25718
rect -158 24530 -100 24542
rect 100 25718 158 25730
rect 100 24542 112 25718
rect 146 24542 158 25718
rect 100 24530 158 24542
rect -158 24282 -100 24294
rect -158 23106 -146 24282
rect -112 23106 -100 24282
rect -158 23094 -100 23106
rect 100 24282 158 24294
rect 100 23106 112 24282
rect 146 23106 158 24282
rect 100 23094 158 23106
rect -158 22846 -100 22858
rect -158 21670 -146 22846
rect -112 21670 -100 22846
rect -158 21658 -100 21670
rect 100 22846 158 22858
rect 100 21670 112 22846
rect 146 21670 158 22846
rect 100 21658 158 21670
rect -158 21410 -100 21422
rect -158 20234 -146 21410
rect -112 20234 -100 21410
rect -158 20222 -100 20234
rect 100 21410 158 21422
rect 100 20234 112 21410
rect 146 20234 158 21410
rect 100 20222 158 20234
rect -158 19974 -100 19986
rect -158 18798 -146 19974
rect -112 18798 -100 19974
rect -158 18786 -100 18798
rect 100 19974 158 19986
rect 100 18798 112 19974
rect 146 18798 158 19974
rect 100 18786 158 18798
rect -158 18538 -100 18550
rect -158 17362 -146 18538
rect -112 17362 -100 18538
rect -158 17350 -100 17362
rect 100 18538 158 18550
rect 100 17362 112 18538
rect 146 17362 158 18538
rect 100 17350 158 17362
rect -158 17102 -100 17114
rect -158 15926 -146 17102
rect -112 15926 -100 17102
rect -158 15914 -100 15926
rect 100 17102 158 17114
rect 100 15926 112 17102
rect 146 15926 158 17102
rect 100 15914 158 15926
rect -158 15666 -100 15678
rect -158 14490 -146 15666
rect -112 14490 -100 15666
rect -158 14478 -100 14490
rect 100 15666 158 15678
rect 100 14490 112 15666
rect 146 14490 158 15666
rect 100 14478 158 14490
rect -158 14230 -100 14242
rect -158 13054 -146 14230
rect -112 13054 -100 14230
rect -158 13042 -100 13054
rect 100 14230 158 14242
rect 100 13054 112 14230
rect 146 13054 158 14230
rect 100 13042 158 13054
rect -158 12794 -100 12806
rect -158 11618 -146 12794
rect -112 11618 -100 12794
rect -158 11606 -100 11618
rect 100 12794 158 12806
rect 100 11618 112 12794
rect 146 11618 158 12794
rect 100 11606 158 11618
rect -158 11358 -100 11370
rect -158 10182 -146 11358
rect -112 10182 -100 11358
rect -158 10170 -100 10182
rect 100 11358 158 11370
rect 100 10182 112 11358
rect 146 10182 158 11358
rect 100 10170 158 10182
rect -158 9922 -100 9934
rect -158 8746 -146 9922
rect -112 8746 -100 9922
rect -158 8734 -100 8746
rect 100 9922 158 9934
rect 100 8746 112 9922
rect 146 8746 158 9922
rect 100 8734 158 8746
rect -158 8486 -100 8498
rect -158 7310 -146 8486
rect -112 7310 -100 8486
rect -158 7298 -100 7310
rect 100 8486 158 8498
rect 100 7310 112 8486
rect 146 7310 158 8486
rect 100 7298 158 7310
rect -158 7050 -100 7062
rect -158 5874 -146 7050
rect -112 5874 -100 7050
rect -158 5862 -100 5874
rect 100 7050 158 7062
rect 100 5874 112 7050
rect 146 5874 158 7050
rect 100 5862 158 5874
rect -158 5614 -100 5626
rect -158 4438 -146 5614
rect -112 4438 -100 5614
rect -158 4426 -100 4438
rect 100 5614 158 5626
rect 100 4438 112 5614
rect 146 4438 158 5614
rect 100 4426 158 4438
rect -158 4178 -100 4190
rect -158 3002 -146 4178
rect -112 3002 -100 4178
rect -158 2990 -100 3002
rect 100 4178 158 4190
rect 100 3002 112 4178
rect 146 3002 158 4178
rect 100 2990 158 3002
rect -158 2742 -100 2754
rect -158 1566 -146 2742
rect -112 1566 -100 2742
rect -158 1554 -100 1566
rect 100 2742 158 2754
rect 100 1566 112 2742
rect 146 1566 158 2742
rect 100 1554 158 1566
rect -158 1306 -100 1318
rect -158 130 -146 1306
rect -112 130 -100 1306
rect -158 118 -100 130
rect 100 1306 158 1318
rect 100 130 112 1306
rect 146 130 158 1306
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -1306 -146 -130
rect -112 -1306 -100 -130
rect -158 -1318 -100 -1306
rect 100 -130 158 -118
rect 100 -1306 112 -130
rect 146 -1306 158 -130
rect 100 -1318 158 -1306
rect -158 -1566 -100 -1554
rect -158 -2742 -146 -1566
rect -112 -2742 -100 -1566
rect -158 -2754 -100 -2742
rect 100 -1566 158 -1554
rect 100 -2742 112 -1566
rect 146 -2742 158 -1566
rect 100 -2754 158 -2742
rect -158 -3002 -100 -2990
rect -158 -4178 -146 -3002
rect -112 -4178 -100 -3002
rect -158 -4190 -100 -4178
rect 100 -3002 158 -2990
rect 100 -4178 112 -3002
rect 146 -4178 158 -3002
rect 100 -4190 158 -4178
rect -158 -4438 -100 -4426
rect -158 -5614 -146 -4438
rect -112 -5614 -100 -4438
rect -158 -5626 -100 -5614
rect 100 -4438 158 -4426
rect 100 -5614 112 -4438
rect 146 -5614 158 -4438
rect 100 -5626 158 -5614
rect -158 -5874 -100 -5862
rect -158 -7050 -146 -5874
rect -112 -7050 -100 -5874
rect -158 -7062 -100 -7050
rect 100 -5874 158 -5862
rect 100 -7050 112 -5874
rect 146 -7050 158 -5874
rect 100 -7062 158 -7050
rect -158 -7310 -100 -7298
rect -158 -8486 -146 -7310
rect -112 -8486 -100 -7310
rect -158 -8498 -100 -8486
rect 100 -7310 158 -7298
rect 100 -8486 112 -7310
rect 146 -8486 158 -7310
rect 100 -8498 158 -8486
rect -158 -8746 -100 -8734
rect -158 -9922 -146 -8746
rect -112 -9922 -100 -8746
rect -158 -9934 -100 -9922
rect 100 -8746 158 -8734
rect 100 -9922 112 -8746
rect 146 -9922 158 -8746
rect 100 -9934 158 -9922
rect -158 -10182 -100 -10170
rect -158 -11358 -146 -10182
rect -112 -11358 -100 -10182
rect -158 -11370 -100 -11358
rect 100 -10182 158 -10170
rect 100 -11358 112 -10182
rect 146 -11358 158 -10182
rect 100 -11370 158 -11358
rect -158 -11618 -100 -11606
rect -158 -12794 -146 -11618
rect -112 -12794 -100 -11618
rect -158 -12806 -100 -12794
rect 100 -11618 158 -11606
rect 100 -12794 112 -11618
rect 146 -12794 158 -11618
rect 100 -12806 158 -12794
rect -158 -13054 -100 -13042
rect -158 -14230 -146 -13054
rect -112 -14230 -100 -13054
rect -158 -14242 -100 -14230
rect 100 -13054 158 -13042
rect 100 -14230 112 -13054
rect 146 -14230 158 -13054
rect 100 -14242 158 -14230
rect -158 -14490 -100 -14478
rect -158 -15666 -146 -14490
rect -112 -15666 -100 -14490
rect -158 -15678 -100 -15666
rect 100 -14490 158 -14478
rect 100 -15666 112 -14490
rect 146 -15666 158 -14490
rect 100 -15678 158 -15666
rect -158 -15926 -100 -15914
rect -158 -17102 -146 -15926
rect -112 -17102 -100 -15926
rect -158 -17114 -100 -17102
rect 100 -15926 158 -15914
rect 100 -17102 112 -15926
rect 146 -17102 158 -15926
rect 100 -17114 158 -17102
rect -158 -17362 -100 -17350
rect -158 -18538 -146 -17362
rect -112 -18538 -100 -17362
rect -158 -18550 -100 -18538
rect 100 -17362 158 -17350
rect 100 -18538 112 -17362
rect 146 -18538 158 -17362
rect 100 -18550 158 -18538
rect -158 -18798 -100 -18786
rect -158 -19974 -146 -18798
rect -112 -19974 -100 -18798
rect -158 -19986 -100 -19974
rect 100 -18798 158 -18786
rect 100 -19974 112 -18798
rect 146 -19974 158 -18798
rect 100 -19986 158 -19974
rect -158 -20234 -100 -20222
rect -158 -21410 -146 -20234
rect -112 -21410 -100 -20234
rect -158 -21422 -100 -21410
rect 100 -20234 158 -20222
rect 100 -21410 112 -20234
rect 146 -21410 158 -20234
rect 100 -21422 158 -21410
rect -158 -21670 -100 -21658
rect -158 -22846 -146 -21670
rect -112 -22846 -100 -21670
rect -158 -22858 -100 -22846
rect 100 -21670 158 -21658
rect 100 -22846 112 -21670
rect 146 -22846 158 -21670
rect 100 -22858 158 -22846
rect -158 -23106 -100 -23094
rect -158 -24282 -146 -23106
rect -112 -24282 -100 -23106
rect -158 -24294 -100 -24282
rect 100 -23106 158 -23094
rect 100 -24282 112 -23106
rect 146 -24282 158 -23106
rect 100 -24294 158 -24282
rect -158 -24542 -100 -24530
rect -158 -25718 -146 -24542
rect -112 -25718 -100 -24542
rect -158 -25730 -100 -25718
rect 100 -24542 158 -24530
rect 100 -25718 112 -24542
rect 146 -25718 158 -24542
rect 100 -25730 158 -25718
rect -158 -25978 -100 -25966
rect -158 -27154 -146 -25978
rect -112 -27154 -100 -25978
rect -158 -27166 -100 -27154
rect 100 -25978 158 -25966
rect 100 -27154 112 -25978
rect 146 -27154 158 -25978
rect 100 -27166 158 -27154
rect -158 -27414 -100 -27402
rect -158 -28590 -146 -27414
rect -112 -28590 -100 -27414
rect -158 -28602 -100 -28590
rect 100 -27414 158 -27402
rect 100 -28590 112 -27414
rect 146 -28590 158 -27414
rect 100 -28602 158 -28590
rect -158 -28850 -100 -28838
rect -158 -30026 -146 -28850
rect -112 -30026 -100 -28850
rect -158 -30038 -100 -30026
rect 100 -28850 158 -28838
rect 100 -30026 112 -28850
rect 146 -30026 158 -28850
rect 100 -30038 158 -30026
rect -158 -30286 -100 -30274
rect -158 -31462 -146 -30286
rect -112 -31462 -100 -30286
rect -158 -31474 -100 -31462
rect 100 -30286 158 -30274
rect 100 -31462 112 -30286
rect 146 -31462 158 -30286
rect 100 -31474 158 -31462
rect -158 -31722 -100 -31710
rect -158 -32898 -146 -31722
rect -112 -32898 -100 -31722
rect -158 -32910 -100 -32898
rect 100 -31722 158 -31710
rect 100 -32898 112 -31722
rect 146 -32898 158 -31722
rect 100 -32910 158 -32898
rect -158 -33158 -100 -33146
rect -158 -34334 -146 -33158
rect -112 -34334 -100 -33158
rect -158 -34346 -100 -34334
rect 100 -33158 158 -33146
rect 100 -34334 112 -33158
rect 146 -34334 158 -33158
rect 100 -34346 158 -34334
rect -158 -34594 -100 -34582
rect -158 -35770 -146 -34594
rect -112 -35770 -100 -34594
rect -158 -35782 -100 -35770
rect 100 -34594 158 -34582
rect 100 -35770 112 -34594
rect 146 -35770 158 -34594
rect 100 -35782 158 -35770
rect -158 -36030 -100 -36018
rect -158 -37206 -146 -36030
rect -112 -37206 -100 -36030
rect -158 -37218 -100 -37206
rect 100 -36030 158 -36018
rect 100 -37206 112 -36030
rect 146 -37206 158 -36030
rect 100 -37218 158 -37206
rect -158 -37466 -100 -37454
rect -158 -38642 -146 -37466
rect -112 -38642 -100 -37466
rect -158 -38654 -100 -38642
rect 100 -37466 158 -37454
rect 100 -38642 112 -37466
rect 146 -38642 158 -37466
rect 100 -38654 158 -38642
rect -158 -38902 -100 -38890
rect -158 -40078 -146 -38902
rect -112 -40078 -100 -38902
rect -158 -40090 -100 -40078
rect 100 -38902 158 -38890
rect 100 -40078 112 -38902
rect 146 -40078 158 -38902
rect 100 -40090 158 -40078
rect -158 -40338 -100 -40326
rect -158 -41514 -146 -40338
rect -112 -41514 -100 -40338
rect -158 -41526 -100 -41514
rect 100 -40338 158 -40326
rect 100 -41514 112 -40338
rect 146 -41514 158 -40338
rect 100 -41526 158 -41514
rect -158 -41774 -100 -41762
rect -158 -42950 -146 -41774
rect -112 -42950 -100 -41774
rect -158 -42962 -100 -42950
rect 100 -41774 158 -41762
rect 100 -42950 112 -41774
rect 146 -42950 158 -41774
rect 100 -42962 158 -42950
rect -158 -43210 -100 -43198
rect -158 -44386 -146 -43210
rect -112 -44386 -100 -43210
rect -158 -44398 -100 -44386
rect 100 -43210 158 -43198
rect 100 -44386 112 -43210
rect 146 -44386 158 -43210
rect 100 -44398 158 -44386
rect -158 -44646 -100 -44634
rect -158 -45822 -146 -44646
rect -112 -45822 -100 -44646
rect -158 -45834 -100 -45822
rect 100 -44646 158 -44634
rect 100 -45822 112 -44646
rect 146 -45822 158 -44646
rect 100 -45834 158 -45822
rect -158 -46082 -100 -46070
rect -158 -47258 -146 -46082
rect -112 -47258 -100 -46082
rect -158 -47270 -100 -47258
rect 100 -46082 158 -46070
rect 100 -47258 112 -46082
rect 146 -47258 158 -46082
rect 100 -47270 158 -47258
rect -158 -47518 -100 -47506
rect -158 -48694 -146 -47518
rect -112 -48694 -100 -47518
rect -158 -48706 -100 -48694
rect 100 -47518 158 -47506
rect 100 -48694 112 -47518
rect 146 -48694 158 -47518
rect 100 -48706 158 -48694
rect -158 -48954 -100 -48942
rect -158 -50130 -146 -48954
rect -112 -50130 -100 -48954
rect -158 -50142 -100 -50130
rect 100 -48954 158 -48942
rect 100 -50130 112 -48954
rect 146 -50130 158 -48954
rect 100 -50142 158 -50130
rect -158 -50390 -100 -50378
rect -158 -51566 -146 -50390
rect -112 -51566 -100 -50390
rect -158 -51578 -100 -51566
rect 100 -50390 158 -50378
rect 100 -51566 112 -50390
rect 146 -51566 158 -50390
rect 100 -51578 158 -51566
rect -158 -51826 -100 -51814
rect -158 -53002 -146 -51826
rect -112 -53002 -100 -51826
rect -158 -53014 -100 -53002
rect 100 -51826 158 -51814
rect 100 -53002 112 -51826
rect 146 -53002 158 -51826
rect 100 -53014 158 -53002
rect -158 -53262 -100 -53250
rect -158 -54438 -146 -53262
rect -112 -54438 -100 -53262
rect -158 -54450 -100 -54438
rect 100 -53262 158 -53250
rect 100 -54438 112 -53262
rect 146 -54438 158 -53262
rect 100 -54450 158 -54438
rect -158 -54698 -100 -54686
rect -158 -55874 -146 -54698
rect -112 -55874 -100 -54698
rect -158 -55886 -100 -55874
rect 100 -54698 158 -54686
rect 100 -55874 112 -54698
rect 146 -55874 158 -54698
rect 100 -55886 158 -55874
rect -158 -56134 -100 -56122
rect -158 -57310 -146 -56134
rect -112 -57310 -100 -56134
rect -158 -57322 -100 -57310
rect 100 -56134 158 -56122
rect 100 -57310 112 -56134
rect 146 -57310 158 -56134
rect 100 -57322 158 -57310
rect -158 -57570 -100 -57558
rect -158 -58746 -146 -57570
rect -112 -58746 -100 -57570
rect -158 -58758 -100 -58746
rect 100 -57570 158 -57558
rect 100 -58746 112 -57570
rect 146 -58746 158 -57570
rect 100 -58758 158 -58746
rect -158 -59006 -100 -58994
rect -158 -60182 -146 -59006
rect -112 -60182 -100 -59006
rect -158 -60194 -100 -60182
rect 100 -59006 158 -58994
rect 100 -60182 112 -59006
rect 146 -60182 158 -59006
rect 100 -60194 158 -60182
rect -158 -60442 -100 -60430
rect -158 -61618 -146 -60442
rect -112 -61618 -100 -60442
rect -158 -61630 -100 -61618
rect 100 -60442 158 -60430
rect 100 -61618 112 -60442
rect 146 -61618 158 -60442
rect 100 -61630 158 -61618
rect -158 -61878 -100 -61866
rect -158 -63054 -146 -61878
rect -112 -63054 -100 -61878
rect -158 -63066 -100 -63054
rect 100 -61878 158 -61866
rect 100 -63054 112 -61878
rect 146 -63054 158 -61878
rect 100 -63066 158 -63054
rect -158 -63314 -100 -63302
rect -158 -64490 -146 -63314
rect -112 -64490 -100 -63314
rect -158 -64502 -100 -64490
rect 100 -63314 158 -63302
rect 100 -64490 112 -63314
rect 146 -64490 158 -63314
rect 100 -64502 158 -64490
rect -158 -64750 -100 -64738
rect -158 -65926 -146 -64750
rect -112 -65926 -100 -64750
rect -158 -65938 -100 -65926
rect 100 -64750 158 -64738
rect 100 -65926 112 -64750
rect 146 -65926 158 -64750
rect 100 -65938 158 -65926
rect -158 -66186 -100 -66174
rect -158 -67362 -146 -66186
rect -112 -67362 -100 -66186
rect -158 -67374 -100 -67362
rect 100 -66186 158 -66174
rect 100 -67362 112 -66186
rect 146 -67362 158 -66186
rect 100 -67374 158 -67362
rect -158 -67622 -100 -67610
rect -158 -68798 -146 -67622
rect -112 -68798 -100 -67622
rect -158 -68810 -100 -68798
rect 100 -67622 158 -67610
rect 100 -68798 112 -67622
rect 146 -68798 158 -67622
rect 100 -68810 158 -68798
rect -158 -69058 -100 -69046
rect -158 -70234 -146 -69058
rect -112 -70234 -100 -69058
rect -158 -70246 -100 -70234
rect 100 -69058 158 -69046
rect 100 -70234 112 -69058
rect 146 -70234 158 -69058
rect 100 -70246 158 -70234
rect -158 -70494 -100 -70482
rect -158 -71670 -146 -70494
rect -112 -71670 -100 -70494
rect -158 -71682 -100 -71670
rect 100 -70494 158 -70482
rect 100 -71670 112 -70494
rect 146 -71670 158 -70494
rect 100 -71682 158 -71670
rect -158 -71930 -100 -71918
rect -158 -73106 -146 -71930
rect -112 -73106 -100 -71930
rect -158 -73118 -100 -73106
rect 100 -71930 158 -71918
rect 100 -73106 112 -71930
rect 146 -73106 158 -71930
rect 100 -73118 158 -73106
rect -158 -73366 -100 -73354
rect -158 -74542 -146 -73366
rect -112 -74542 -100 -73366
rect -158 -74554 -100 -74542
rect 100 -73366 158 -73354
rect 100 -74542 112 -73366
rect 146 -74542 158 -73366
rect 100 -74554 158 -74542
rect -158 -74802 -100 -74790
rect -158 -75978 -146 -74802
rect -112 -75978 -100 -74802
rect -158 -75990 -100 -75978
rect 100 -74802 158 -74790
rect 100 -75978 112 -74802
rect 146 -75978 158 -74802
rect 100 -75990 158 -75978
rect -158 -76238 -100 -76226
rect -158 -77414 -146 -76238
rect -112 -77414 -100 -76238
rect -158 -77426 -100 -77414
rect 100 -76238 158 -76226
rect 100 -77414 112 -76238
rect 146 -77414 158 -76238
rect 100 -77426 158 -77414
rect -158 -77674 -100 -77662
rect -158 -78850 -146 -77674
rect -112 -78850 -100 -77674
rect -158 -78862 -100 -78850
rect 100 -77674 158 -77662
rect 100 -78850 112 -77674
rect 146 -78850 158 -77674
rect 100 -78862 158 -78850
rect -158 -79110 -100 -79098
rect -158 -80286 -146 -79110
rect -112 -80286 -100 -79110
rect -158 -80298 -100 -80286
rect 100 -79110 158 -79098
rect 100 -80286 112 -79110
rect 146 -80286 158 -79110
rect 100 -80298 158 -80286
rect -158 -80546 -100 -80534
rect -158 -81722 -146 -80546
rect -112 -81722 -100 -80546
rect -158 -81734 -100 -81722
rect 100 -80546 158 -80534
rect 100 -81722 112 -80546
rect 146 -81722 158 -80546
rect 100 -81734 158 -81722
rect -158 -81982 -100 -81970
rect -158 -83158 -146 -81982
rect -112 -83158 -100 -81982
rect -158 -83170 -100 -83158
rect 100 -81982 158 -81970
rect 100 -83158 112 -81982
rect 146 -83158 158 -81982
rect 100 -83170 158 -83158
rect -158 -83418 -100 -83406
rect -158 -84594 -146 -83418
rect -112 -84594 -100 -83418
rect -158 -84606 -100 -84594
rect 100 -83418 158 -83406
rect 100 -84594 112 -83418
rect 146 -84594 158 -83418
rect 100 -84606 158 -84594
rect -158 -84854 -100 -84842
rect -158 -86030 -146 -84854
rect -112 -86030 -100 -84854
rect -158 -86042 -100 -86030
rect 100 -84854 158 -84842
rect 100 -86030 112 -84854
rect 146 -86030 158 -84854
rect 100 -86042 158 -86030
rect -158 -86290 -100 -86278
rect -158 -87466 -146 -86290
rect -112 -87466 -100 -86290
rect -158 -87478 -100 -87466
rect 100 -86290 158 -86278
rect 100 -87466 112 -86290
rect 146 -87466 158 -86290
rect 100 -87478 158 -87466
rect -158 -87726 -100 -87714
rect -158 -88902 -146 -87726
rect -112 -88902 -100 -87726
rect -158 -88914 -100 -88902
rect 100 -87726 158 -87714
rect 100 -88902 112 -87726
rect 146 -88902 158 -87726
rect 100 -88914 158 -88902
rect -158 -89162 -100 -89150
rect -158 -90338 -146 -89162
rect -112 -90338 -100 -89162
rect -158 -90350 -100 -90338
rect 100 -89162 158 -89150
rect 100 -90338 112 -89162
rect 146 -90338 158 -89162
rect 100 -90350 158 -90338
rect -158 -90598 -100 -90586
rect -158 -91774 -146 -90598
rect -112 -91774 -100 -90598
rect -158 -91786 -100 -91774
rect 100 -90598 158 -90586
rect 100 -91774 112 -90598
rect 146 -91774 158 -90598
rect 100 -91786 158 -91774
rect -158 -92034 -100 -92022
rect -158 -93210 -146 -92034
rect -112 -93210 -100 -92034
rect -158 -93222 -100 -93210
rect 100 -92034 158 -92022
rect 100 -93210 112 -92034
rect 146 -93210 158 -92034
rect 100 -93222 158 -93210
rect -158 -93470 -100 -93458
rect -158 -94646 -146 -93470
rect -112 -94646 -100 -93470
rect -158 -94658 -100 -94646
rect 100 -93470 158 -93458
rect 100 -94646 112 -93470
rect 146 -94646 158 -93470
rect 100 -94658 158 -94646
rect -158 -94906 -100 -94894
rect -158 -96082 -146 -94906
rect -112 -96082 -100 -94906
rect -158 -96094 -100 -96082
rect 100 -94906 158 -94894
rect 100 -96082 112 -94906
rect 146 -96082 158 -94906
rect 100 -96094 158 -96082
rect -158 -96342 -100 -96330
rect -158 -97518 -146 -96342
rect -112 -97518 -100 -96342
rect -158 -97530 -100 -97518
rect 100 -96342 158 -96330
rect 100 -97518 112 -96342
rect 146 -97518 158 -96342
rect 100 -97530 158 -97518
rect -158 -97778 -100 -97766
rect -158 -98954 -146 -97778
rect -112 -98954 -100 -97778
rect -158 -98966 -100 -98954
rect 100 -97778 158 -97766
rect 100 -98954 112 -97778
rect 146 -98954 158 -97778
rect 100 -98966 158 -98954
rect -158 -99214 -100 -99202
rect -158 -100390 -146 -99214
rect -112 -100390 -100 -99214
rect -158 -100402 -100 -100390
rect 100 -99214 158 -99202
rect 100 -100390 112 -99214
rect 146 -100390 158 -99214
rect 100 -100402 158 -100390
rect -158 -100650 -100 -100638
rect -158 -101826 -146 -100650
rect -112 -101826 -100 -100650
rect -158 -101838 -100 -101826
rect 100 -100650 158 -100638
rect 100 -101826 112 -100650
rect 146 -101826 158 -100650
rect 100 -101838 158 -101826
rect -158 -102086 -100 -102074
rect -158 -103262 -146 -102086
rect -112 -103262 -100 -102086
rect -158 -103274 -100 -103262
rect 100 -102086 158 -102074
rect 100 -103262 112 -102086
rect 146 -103262 158 -102086
rect 100 -103274 158 -103262
rect -158 -103522 -100 -103510
rect -158 -104698 -146 -103522
rect -112 -104698 -100 -103522
rect -158 -104710 -100 -104698
rect 100 -103522 158 -103510
rect 100 -104698 112 -103522
rect 146 -104698 158 -103522
rect 100 -104710 158 -104698
rect -158 -104958 -100 -104946
rect -158 -106134 -146 -104958
rect -112 -106134 -100 -104958
rect -158 -106146 -100 -106134
rect 100 -104958 158 -104946
rect 100 -106134 112 -104958
rect 146 -106134 158 -104958
rect 100 -106146 158 -106134
rect -158 -106394 -100 -106382
rect -158 -107570 -146 -106394
rect -112 -107570 -100 -106394
rect -158 -107582 -100 -107570
rect 100 -106394 158 -106382
rect 100 -107570 112 -106394
rect 146 -107570 158 -106394
rect 100 -107582 158 -107570
rect -158 -107830 -100 -107818
rect -158 -109006 -146 -107830
rect -112 -109006 -100 -107830
rect -158 -109018 -100 -109006
rect 100 -107830 158 -107818
rect 100 -109006 112 -107830
rect 146 -109006 158 -107830
rect 100 -109018 158 -109006
rect -158 -109266 -100 -109254
rect -158 -110442 -146 -109266
rect -112 -110442 -100 -109266
rect -158 -110454 -100 -110442
rect 100 -109266 158 -109254
rect 100 -110442 112 -109266
rect 146 -110442 158 -109266
rect 100 -110454 158 -110442
rect -158 -110702 -100 -110690
rect -158 -111878 -146 -110702
rect -112 -111878 -100 -110702
rect -158 -111890 -100 -111878
rect 100 -110702 158 -110690
rect 100 -111878 112 -110702
rect 146 -111878 158 -110702
rect 100 -111890 158 -111878
rect -158 -112138 -100 -112126
rect -158 -113314 -146 -112138
rect -112 -113314 -100 -112138
rect -158 -113326 -100 -113314
rect 100 -112138 158 -112126
rect 100 -113314 112 -112138
rect 146 -113314 158 -112138
rect 100 -113326 158 -113314
rect -158 -113574 -100 -113562
rect -158 -114750 -146 -113574
rect -112 -114750 -100 -113574
rect -158 -114762 -100 -114750
rect 100 -113574 158 -113562
rect 100 -114750 112 -113574
rect 146 -114750 158 -113574
rect 100 -114762 158 -114750
rect -158 -115010 -100 -114998
rect -158 -116186 -146 -115010
rect -112 -116186 -100 -115010
rect -158 -116198 -100 -116186
rect 100 -115010 158 -114998
rect 100 -116186 112 -115010
rect 146 -116186 158 -115010
rect 100 -116198 158 -116186
rect -158 -116446 -100 -116434
rect -158 -117622 -146 -116446
rect -112 -117622 -100 -116446
rect -158 -117634 -100 -117622
rect 100 -116446 158 -116434
rect 100 -117622 112 -116446
rect 146 -117622 158 -116446
rect 100 -117634 158 -117622
rect -158 -117882 -100 -117870
rect -158 -119058 -146 -117882
rect -112 -119058 -100 -117882
rect -158 -119070 -100 -119058
rect 100 -117882 158 -117870
rect 100 -119058 112 -117882
rect 146 -119058 158 -117882
rect 100 -119070 158 -119058
rect -158 -119318 -100 -119306
rect -158 -120494 -146 -119318
rect -112 -120494 -100 -119318
rect -158 -120506 -100 -120494
rect 100 -119318 158 -119306
rect 100 -120494 112 -119318
rect 146 -120494 158 -119318
rect 100 -120506 158 -120494
rect -158 -120754 -100 -120742
rect -158 -121930 -146 -120754
rect -112 -121930 -100 -120754
rect -158 -121942 -100 -121930
rect 100 -120754 158 -120742
rect 100 -121930 112 -120754
rect 146 -121930 158 -120754
rect 100 -121942 158 -121930
rect -158 -122190 -100 -122178
rect -158 -123366 -146 -122190
rect -112 -123366 -100 -122190
rect -158 -123378 -100 -123366
rect 100 -122190 158 -122178
rect 100 -123366 112 -122190
rect 146 -123366 158 -122190
rect 100 -123378 158 -123366
rect -158 -123626 -100 -123614
rect -158 -124802 -146 -123626
rect -112 -124802 -100 -123626
rect -158 -124814 -100 -124802
rect 100 -123626 158 -123614
rect 100 -124802 112 -123626
rect 146 -124802 158 -123626
rect 100 -124814 158 -124802
rect -158 -125062 -100 -125050
rect -158 -126238 -146 -125062
rect -112 -126238 -100 -125062
rect -158 -126250 -100 -126238
rect 100 -125062 158 -125050
rect 100 -126238 112 -125062
rect 146 -126238 158 -125062
rect 100 -126250 158 -126238
rect -158 -126498 -100 -126486
rect -158 -127674 -146 -126498
rect -112 -127674 -100 -126498
rect -158 -127686 -100 -127674
rect 100 -126498 158 -126486
rect 100 -127674 112 -126498
rect 146 -127674 158 -126498
rect 100 -127686 158 -127674
rect -158 -127934 -100 -127922
rect -158 -129110 -146 -127934
rect -112 -129110 -100 -127934
rect -158 -129122 -100 -129110
rect 100 -127934 158 -127922
rect 100 -129110 112 -127934
rect 146 -129110 158 -127934
rect 100 -129122 158 -129110
rect -158 -129370 -100 -129358
rect -158 -130546 -146 -129370
rect -112 -130546 -100 -129370
rect -158 -130558 -100 -130546
rect 100 -129370 158 -129358
rect 100 -130546 112 -129370
rect 146 -130546 158 -129370
rect 100 -130558 158 -130546
rect -158 -130806 -100 -130794
rect -158 -131982 -146 -130806
rect -112 -131982 -100 -130806
rect -158 -131994 -100 -131982
rect 100 -130806 158 -130794
rect 100 -131982 112 -130806
rect 146 -131982 158 -130806
rect 100 -131994 158 -131982
rect -158 -132242 -100 -132230
rect -158 -133418 -146 -132242
rect -112 -133418 -100 -132242
rect -158 -133430 -100 -133418
rect 100 -132242 158 -132230
rect 100 -133418 112 -132242
rect 146 -133418 158 -132242
rect 100 -133430 158 -133418
rect -158 -133678 -100 -133666
rect -158 -134854 -146 -133678
rect -112 -134854 -100 -133678
rect -158 -134866 -100 -134854
rect 100 -133678 158 -133666
rect 100 -134854 112 -133678
rect 146 -134854 158 -133678
rect 100 -134866 158 -134854
rect -158 -135114 -100 -135102
rect -158 -136290 -146 -135114
rect -112 -136290 -100 -135114
rect -158 -136302 -100 -136290
rect 100 -135114 158 -135102
rect 100 -136290 112 -135114
rect 146 -136290 158 -135114
rect 100 -136302 158 -136290
rect -158 -136550 -100 -136538
rect -158 -137726 -146 -136550
rect -112 -137726 -100 -136550
rect -158 -137738 -100 -137726
rect 100 -136550 158 -136538
rect 100 -137726 112 -136550
rect 146 -137726 158 -136550
rect 100 -137738 158 -137726
rect -158 -137986 -100 -137974
rect -158 -139162 -146 -137986
rect -112 -139162 -100 -137986
rect -158 -139174 -100 -139162
rect 100 -137986 158 -137974
rect 100 -139162 112 -137986
rect 146 -139162 158 -137986
rect 100 -139174 158 -139162
rect -158 -139422 -100 -139410
rect -158 -140598 -146 -139422
rect -112 -140598 -100 -139422
rect -158 -140610 -100 -140598
rect 100 -139422 158 -139410
rect 100 -140598 112 -139422
rect 146 -140598 158 -139422
rect 100 -140610 158 -140598
rect -158 -140858 -100 -140846
rect -158 -142034 -146 -140858
rect -112 -142034 -100 -140858
rect -158 -142046 -100 -142034
rect 100 -140858 158 -140846
rect 100 -142034 112 -140858
rect 146 -142034 158 -140858
rect 100 -142046 158 -142034
rect -158 -142294 -100 -142282
rect -158 -143470 -146 -142294
rect -112 -143470 -100 -142294
rect -158 -143482 -100 -143470
rect 100 -142294 158 -142282
rect 100 -143470 112 -142294
rect 146 -143470 158 -142294
rect 100 -143482 158 -143470
rect -158 -143730 -100 -143718
rect -158 -144906 -146 -143730
rect -112 -144906 -100 -143730
rect -158 -144918 -100 -144906
rect 100 -143730 158 -143718
rect 100 -144906 112 -143730
rect 146 -144906 158 -143730
rect 100 -144918 158 -144906
rect -158 -145166 -100 -145154
rect -158 -146342 -146 -145166
rect -112 -146342 -100 -145166
rect -158 -146354 -100 -146342
rect 100 -145166 158 -145154
rect 100 -146342 112 -145166
rect 146 -146342 158 -145166
rect 100 -146354 158 -146342
rect -158 -146602 -100 -146590
rect -158 -147778 -146 -146602
rect -112 -147778 -100 -146602
rect -158 -147790 -100 -147778
rect 100 -146602 158 -146590
rect 100 -147778 112 -146602
rect 146 -147778 158 -146602
rect 100 -147790 158 -147778
rect -158 -148038 -100 -148026
rect -158 -149214 -146 -148038
rect -112 -149214 -100 -148038
rect -158 -149226 -100 -149214
rect 100 -148038 158 -148026
rect 100 -149214 112 -148038
rect 146 -149214 158 -148038
rect 100 -149226 158 -149214
rect -158 -149474 -100 -149462
rect -158 -150650 -146 -149474
rect -112 -150650 -100 -149474
rect -158 -150662 -100 -150650
rect 100 -149474 158 -149462
rect 100 -150650 112 -149474
rect 146 -150650 158 -149474
rect 100 -150662 158 -150650
rect -158 -150910 -100 -150898
rect -158 -152086 -146 -150910
rect -112 -152086 -100 -150910
rect -158 -152098 -100 -152086
rect 100 -150910 158 -150898
rect 100 -152086 112 -150910
rect 146 -152086 158 -150910
rect 100 -152098 158 -152086
rect -158 -152346 -100 -152334
rect -158 -153522 -146 -152346
rect -112 -153522 -100 -152346
rect -158 -153534 -100 -153522
rect 100 -152346 158 -152334
rect 100 -153522 112 -152346
rect 146 -153522 158 -152346
rect 100 -153534 158 -153522
rect -158 -153782 -100 -153770
rect -158 -154958 -146 -153782
rect -112 -154958 -100 -153782
rect -158 -154970 -100 -154958
rect 100 -153782 158 -153770
rect 100 -154958 112 -153782
rect 146 -154958 158 -153782
rect 100 -154970 158 -154958
rect -158 -155218 -100 -155206
rect -158 -156394 -146 -155218
rect -112 -156394 -100 -155218
rect -158 -156406 -100 -156394
rect 100 -155218 158 -155206
rect 100 -156394 112 -155218
rect 146 -156394 158 -155218
rect 100 -156406 158 -156394
rect -158 -156654 -100 -156642
rect -158 -157830 -146 -156654
rect -112 -157830 -100 -156654
rect -158 -157842 -100 -157830
rect 100 -156654 158 -156642
rect 100 -157830 112 -156654
rect 146 -157830 158 -156654
rect 100 -157842 158 -157830
rect -158 -158090 -100 -158078
rect -158 -159266 -146 -158090
rect -112 -159266 -100 -158090
rect -158 -159278 -100 -159266
rect 100 -158090 158 -158078
rect 100 -159266 112 -158090
rect 146 -159266 158 -158090
rect 100 -159278 158 -159266
rect -158 -159526 -100 -159514
rect -158 -160702 -146 -159526
rect -112 -160702 -100 -159526
rect -158 -160714 -100 -160702
rect 100 -159526 158 -159514
rect 100 -160702 112 -159526
rect 146 -160702 158 -159526
rect 100 -160714 158 -160702
rect -158 -160962 -100 -160950
rect -158 -162138 -146 -160962
rect -112 -162138 -100 -160962
rect -158 -162150 -100 -162138
rect 100 -160962 158 -160950
rect 100 -162138 112 -160962
rect 146 -162138 158 -160962
rect 100 -162150 158 -162138
rect -158 -162398 -100 -162386
rect -158 -163574 -146 -162398
rect -112 -163574 -100 -162398
rect -158 -163586 -100 -163574
rect 100 -162398 158 -162386
rect 100 -163574 112 -162398
rect 146 -163574 158 -162398
rect 100 -163586 158 -163574
rect -158 -163834 -100 -163822
rect -158 -165010 -146 -163834
rect -112 -165010 -100 -163834
rect -158 -165022 -100 -165010
rect 100 -163834 158 -163822
rect 100 -165010 112 -163834
rect 146 -165010 158 -163834
rect 100 -165022 158 -165010
rect -158 -165270 -100 -165258
rect -158 -166446 -146 -165270
rect -112 -166446 -100 -165270
rect -158 -166458 -100 -166446
rect 100 -165270 158 -165258
rect 100 -166446 112 -165270
rect 146 -166446 158 -165270
rect 100 -166458 158 -166446
rect -158 -166706 -100 -166694
rect -158 -167882 -146 -166706
rect -112 -167882 -100 -166706
rect -158 -167894 -100 -167882
rect 100 -166706 158 -166694
rect 100 -167882 112 -166706
rect 146 -167882 158 -166706
rect 100 -167894 158 -167882
rect -158 -168142 -100 -168130
rect -158 -169318 -146 -168142
rect -112 -169318 -100 -168142
rect -158 -169330 -100 -169318
rect 100 -168142 158 -168130
rect 100 -169318 112 -168142
rect 146 -169318 158 -168142
rect 100 -169330 158 -169318
rect -158 -169578 -100 -169566
rect -158 -170754 -146 -169578
rect -112 -170754 -100 -169578
rect -158 -170766 -100 -170754
rect 100 -169578 158 -169566
rect 100 -170754 112 -169578
rect 146 -170754 158 -169578
rect 100 -170766 158 -170754
rect -158 -171014 -100 -171002
rect -158 -172190 -146 -171014
rect -112 -172190 -100 -171014
rect -158 -172202 -100 -172190
rect 100 -171014 158 -171002
rect 100 -172190 112 -171014
rect 146 -172190 158 -171014
rect 100 -172202 158 -172190
rect -158 -172450 -100 -172438
rect -158 -173626 -146 -172450
rect -112 -173626 -100 -172450
rect -158 -173638 -100 -173626
rect 100 -172450 158 -172438
rect 100 -173626 112 -172450
rect 146 -173626 158 -172450
rect 100 -173638 158 -173626
rect -158 -173886 -100 -173874
rect -158 -175062 -146 -173886
rect -112 -175062 -100 -173886
rect -158 -175074 -100 -175062
rect 100 -173886 158 -173874
rect 100 -175062 112 -173886
rect 146 -175062 158 -173886
rect 100 -175074 158 -175062
rect -158 -175322 -100 -175310
rect -158 -176498 -146 -175322
rect -112 -176498 -100 -175322
rect -158 -176510 -100 -176498
rect 100 -175322 158 -175310
rect 100 -176498 112 -175322
rect 146 -176498 158 -175322
rect 100 -176510 158 -176498
rect -158 -176758 -100 -176746
rect -158 -177934 -146 -176758
rect -112 -177934 -100 -176758
rect -158 -177946 -100 -177934
rect 100 -176758 158 -176746
rect 100 -177934 112 -176758
rect 146 -177934 158 -176758
rect 100 -177946 158 -177934
rect -158 -178194 -100 -178182
rect -158 -179370 -146 -178194
rect -112 -179370 -100 -178194
rect -158 -179382 -100 -179370
rect 100 -178194 158 -178182
rect 100 -179370 112 -178194
rect 146 -179370 158 -178194
rect 100 -179382 158 -179370
rect -158 -179630 -100 -179618
rect -158 -180806 -146 -179630
rect -112 -180806 -100 -179630
rect -158 -180818 -100 -180806
rect 100 -179630 158 -179618
rect 100 -180806 112 -179630
rect 146 -180806 158 -179630
rect 100 -180818 158 -180806
rect -158 -181066 -100 -181054
rect -158 -182242 -146 -181066
rect -112 -182242 -100 -181066
rect -158 -182254 -100 -182242
rect 100 -181066 158 -181054
rect 100 -182242 112 -181066
rect 146 -182242 158 -181066
rect 100 -182254 158 -182242
rect -158 -182502 -100 -182490
rect -158 -183678 -146 -182502
rect -112 -183678 -100 -182502
rect -158 -183690 -100 -183678
rect 100 -182502 158 -182490
rect 100 -183678 112 -182502
rect 146 -183678 158 -182502
rect 100 -183690 158 -183678
<< mvpdiffc >>
rect -146 182502 -112 183678
rect 112 182502 146 183678
rect -146 181066 -112 182242
rect 112 181066 146 182242
rect -146 179630 -112 180806
rect 112 179630 146 180806
rect -146 178194 -112 179370
rect 112 178194 146 179370
rect -146 176758 -112 177934
rect 112 176758 146 177934
rect -146 175322 -112 176498
rect 112 175322 146 176498
rect -146 173886 -112 175062
rect 112 173886 146 175062
rect -146 172450 -112 173626
rect 112 172450 146 173626
rect -146 171014 -112 172190
rect 112 171014 146 172190
rect -146 169578 -112 170754
rect 112 169578 146 170754
rect -146 168142 -112 169318
rect 112 168142 146 169318
rect -146 166706 -112 167882
rect 112 166706 146 167882
rect -146 165270 -112 166446
rect 112 165270 146 166446
rect -146 163834 -112 165010
rect 112 163834 146 165010
rect -146 162398 -112 163574
rect 112 162398 146 163574
rect -146 160962 -112 162138
rect 112 160962 146 162138
rect -146 159526 -112 160702
rect 112 159526 146 160702
rect -146 158090 -112 159266
rect 112 158090 146 159266
rect -146 156654 -112 157830
rect 112 156654 146 157830
rect -146 155218 -112 156394
rect 112 155218 146 156394
rect -146 153782 -112 154958
rect 112 153782 146 154958
rect -146 152346 -112 153522
rect 112 152346 146 153522
rect -146 150910 -112 152086
rect 112 150910 146 152086
rect -146 149474 -112 150650
rect 112 149474 146 150650
rect -146 148038 -112 149214
rect 112 148038 146 149214
rect -146 146602 -112 147778
rect 112 146602 146 147778
rect -146 145166 -112 146342
rect 112 145166 146 146342
rect -146 143730 -112 144906
rect 112 143730 146 144906
rect -146 142294 -112 143470
rect 112 142294 146 143470
rect -146 140858 -112 142034
rect 112 140858 146 142034
rect -146 139422 -112 140598
rect 112 139422 146 140598
rect -146 137986 -112 139162
rect 112 137986 146 139162
rect -146 136550 -112 137726
rect 112 136550 146 137726
rect -146 135114 -112 136290
rect 112 135114 146 136290
rect -146 133678 -112 134854
rect 112 133678 146 134854
rect -146 132242 -112 133418
rect 112 132242 146 133418
rect -146 130806 -112 131982
rect 112 130806 146 131982
rect -146 129370 -112 130546
rect 112 129370 146 130546
rect -146 127934 -112 129110
rect 112 127934 146 129110
rect -146 126498 -112 127674
rect 112 126498 146 127674
rect -146 125062 -112 126238
rect 112 125062 146 126238
rect -146 123626 -112 124802
rect 112 123626 146 124802
rect -146 122190 -112 123366
rect 112 122190 146 123366
rect -146 120754 -112 121930
rect 112 120754 146 121930
rect -146 119318 -112 120494
rect 112 119318 146 120494
rect -146 117882 -112 119058
rect 112 117882 146 119058
rect -146 116446 -112 117622
rect 112 116446 146 117622
rect -146 115010 -112 116186
rect 112 115010 146 116186
rect -146 113574 -112 114750
rect 112 113574 146 114750
rect -146 112138 -112 113314
rect 112 112138 146 113314
rect -146 110702 -112 111878
rect 112 110702 146 111878
rect -146 109266 -112 110442
rect 112 109266 146 110442
rect -146 107830 -112 109006
rect 112 107830 146 109006
rect -146 106394 -112 107570
rect 112 106394 146 107570
rect -146 104958 -112 106134
rect 112 104958 146 106134
rect -146 103522 -112 104698
rect 112 103522 146 104698
rect -146 102086 -112 103262
rect 112 102086 146 103262
rect -146 100650 -112 101826
rect 112 100650 146 101826
rect -146 99214 -112 100390
rect 112 99214 146 100390
rect -146 97778 -112 98954
rect 112 97778 146 98954
rect -146 96342 -112 97518
rect 112 96342 146 97518
rect -146 94906 -112 96082
rect 112 94906 146 96082
rect -146 93470 -112 94646
rect 112 93470 146 94646
rect -146 92034 -112 93210
rect 112 92034 146 93210
rect -146 90598 -112 91774
rect 112 90598 146 91774
rect -146 89162 -112 90338
rect 112 89162 146 90338
rect -146 87726 -112 88902
rect 112 87726 146 88902
rect -146 86290 -112 87466
rect 112 86290 146 87466
rect -146 84854 -112 86030
rect 112 84854 146 86030
rect -146 83418 -112 84594
rect 112 83418 146 84594
rect -146 81982 -112 83158
rect 112 81982 146 83158
rect -146 80546 -112 81722
rect 112 80546 146 81722
rect -146 79110 -112 80286
rect 112 79110 146 80286
rect -146 77674 -112 78850
rect 112 77674 146 78850
rect -146 76238 -112 77414
rect 112 76238 146 77414
rect -146 74802 -112 75978
rect 112 74802 146 75978
rect -146 73366 -112 74542
rect 112 73366 146 74542
rect -146 71930 -112 73106
rect 112 71930 146 73106
rect -146 70494 -112 71670
rect 112 70494 146 71670
rect -146 69058 -112 70234
rect 112 69058 146 70234
rect -146 67622 -112 68798
rect 112 67622 146 68798
rect -146 66186 -112 67362
rect 112 66186 146 67362
rect -146 64750 -112 65926
rect 112 64750 146 65926
rect -146 63314 -112 64490
rect 112 63314 146 64490
rect -146 61878 -112 63054
rect 112 61878 146 63054
rect -146 60442 -112 61618
rect 112 60442 146 61618
rect -146 59006 -112 60182
rect 112 59006 146 60182
rect -146 57570 -112 58746
rect 112 57570 146 58746
rect -146 56134 -112 57310
rect 112 56134 146 57310
rect -146 54698 -112 55874
rect 112 54698 146 55874
rect -146 53262 -112 54438
rect 112 53262 146 54438
rect -146 51826 -112 53002
rect 112 51826 146 53002
rect -146 50390 -112 51566
rect 112 50390 146 51566
rect -146 48954 -112 50130
rect 112 48954 146 50130
rect -146 47518 -112 48694
rect 112 47518 146 48694
rect -146 46082 -112 47258
rect 112 46082 146 47258
rect -146 44646 -112 45822
rect 112 44646 146 45822
rect -146 43210 -112 44386
rect 112 43210 146 44386
rect -146 41774 -112 42950
rect 112 41774 146 42950
rect -146 40338 -112 41514
rect 112 40338 146 41514
rect -146 38902 -112 40078
rect 112 38902 146 40078
rect -146 37466 -112 38642
rect 112 37466 146 38642
rect -146 36030 -112 37206
rect 112 36030 146 37206
rect -146 34594 -112 35770
rect 112 34594 146 35770
rect -146 33158 -112 34334
rect 112 33158 146 34334
rect -146 31722 -112 32898
rect 112 31722 146 32898
rect -146 30286 -112 31462
rect 112 30286 146 31462
rect -146 28850 -112 30026
rect 112 28850 146 30026
rect -146 27414 -112 28590
rect 112 27414 146 28590
rect -146 25978 -112 27154
rect 112 25978 146 27154
rect -146 24542 -112 25718
rect 112 24542 146 25718
rect -146 23106 -112 24282
rect 112 23106 146 24282
rect -146 21670 -112 22846
rect 112 21670 146 22846
rect -146 20234 -112 21410
rect 112 20234 146 21410
rect -146 18798 -112 19974
rect 112 18798 146 19974
rect -146 17362 -112 18538
rect 112 17362 146 18538
rect -146 15926 -112 17102
rect 112 15926 146 17102
rect -146 14490 -112 15666
rect 112 14490 146 15666
rect -146 13054 -112 14230
rect 112 13054 146 14230
rect -146 11618 -112 12794
rect 112 11618 146 12794
rect -146 10182 -112 11358
rect 112 10182 146 11358
rect -146 8746 -112 9922
rect 112 8746 146 9922
rect -146 7310 -112 8486
rect 112 7310 146 8486
rect -146 5874 -112 7050
rect 112 5874 146 7050
rect -146 4438 -112 5614
rect 112 4438 146 5614
rect -146 3002 -112 4178
rect 112 3002 146 4178
rect -146 1566 -112 2742
rect 112 1566 146 2742
rect -146 130 -112 1306
rect 112 130 146 1306
rect -146 -1306 -112 -130
rect 112 -1306 146 -130
rect -146 -2742 -112 -1566
rect 112 -2742 146 -1566
rect -146 -4178 -112 -3002
rect 112 -4178 146 -3002
rect -146 -5614 -112 -4438
rect 112 -5614 146 -4438
rect -146 -7050 -112 -5874
rect 112 -7050 146 -5874
rect -146 -8486 -112 -7310
rect 112 -8486 146 -7310
rect -146 -9922 -112 -8746
rect 112 -9922 146 -8746
rect -146 -11358 -112 -10182
rect 112 -11358 146 -10182
rect -146 -12794 -112 -11618
rect 112 -12794 146 -11618
rect -146 -14230 -112 -13054
rect 112 -14230 146 -13054
rect -146 -15666 -112 -14490
rect 112 -15666 146 -14490
rect -146 -17102 -112 -15926
rect 112 -17102 146 -15926
rect -146 -18538 -112 -17362
rect 112 -18538 146 -17362
rect -146 -19974 -112 -18798
rect 112 -19974 146 -18798
rect -146 -21410 -112 -20234
rect 112 -21410 146 -20234
rect -146 -22846 -112 -21670
rect 112 -22846 146 -21670
rect -146 -24282 -112 -23106
rect 112 -24282 146 -23106
rect -146 -25718 -112 -24542
rect 112 -25718 146 -24542
rect -146 -27154 -112 -25978
rect 112 -27154 146 -25978
rect -146 -28590 -112 -27414
rect 112 -28590 146 -27414
rect -146 -30026 -112 -28850
rect 112 -30026 146 -28850
rect -146 -31462 -112 -30286
rect 112 -31462 146 -30286
rect -146 -32898 -112 -31722
rect 112 -32898 146 -31722
rect -146 -34334 -112 -33158
rect 112 -34334 146 -33158
rect -146 -35770 -112 -34594
rect 112 -35770 146 -34594
rect -146 -37206 -112 -36030
rect 112 -37206 146 -36030
rect -146 -38642 -112 -37466
rect 112 -38642 146 -37466
rect -146 -40078 -112 -38902
rect 112 -40078 146 -38902
rect -146 -41514 -112 -40338
rect 112 -41514 146 -40338
rect -146 -42950 -112 -41774
rect 112 -42950 146 -41774
rect -146 -44386 -112 -43210
rect 112 -44386 146 -43210
rect -146 -45822 -112 -44646
rect 112 -45822 146 -44646
rect -146 -47258 -112 -46082
rect 112 -47258 146 -46082
rect -146 -48694 -112 -47518
rect 112 -48694 146 -47518
rect -146 -50130 -112 -48954
rect 112 -50130 146 -48954
rect -146 -51566 -112 -50390
rect 112 -51566 146 -50390
rect -146 -53002 -112 -51826
rect 112 -53002 146 -51826
rect -146 -54438 -112 -53262
rect 112 -54438 146 -53262
rect -146 -55874 -112 -54698
rect 112 -55874 146 -54698
rect -146 -57310 -112 -56134
rect 112 -57310 146 -56134
rect -146 -58746 -112 -57570
rect 112 -58746 146 -57570
rect -146 -60182 -112 -59006
rect 112 -60182 146 -59006
rect -146 -61618 -112 -60442
rect 112 -61618 146 -60442
rect -146 -63054 -112 -61878
rect 112 -63054 146 -61878
rect -146 -64490 -112 -63314
rect 112 -64490 146 -63314
rect -146 -65926 -112 -64750
rect 112 -65926 146 -64750
rect -146 -67362 -112 -66186
rect 112 -67362 146 -66186
rect -146 -68798 -112 -67622
rect 112 -68798 146 -67622
rect -146 -70234 -112 -69058
rect 112 -70234 146 -69058
rect -146 -71670 -112 -70494
rect 112 -71670 146 -70494
rect -146 -73106 -112 -71930
rect 112 -73106 146 -71930
rect -146 -74542 -112 -73366
rect 112 -74542 146 -73366
rect -146 -75978 -112 -74802
rect 112 -75978 146 -74802
rect -146 -77414 -112 -76238
rect 112 -77414 146 -76238
rect -146 -78850 -112 -77674
rect 112 -78850 146 -77674
rect -146 -80286 -112 -79110
rect 112 -80286 146 -79110
rect -146 -81722 -112 -80546
rect 112 -81722 146 -80546
rect -146 -83158 -112 -81982
rect 112 -83158 146 -81982
rect -146 -84594 -112 -83418
rect 112 -84594 146 -83418
rect -146 -86030 -112 -84854
rect 112 -86030 146 -84854
rect -146 -87466 -112 -86290
rect 112 -87466 146 -86290
rect -146 -88902 -112 -87726
rect 112 -88902 146 -87726
rect -146 -90338 -112 -89162
rect 112 -90338 146 -89162
rect -146 -91774 -112 -90598
rect 112 -91774 146 -90598
rect -146 -93210 -112 -92034
rect 112 -93210 146 -92034
rect -146 -94646 -112 -93470
rect 112 -94646 146 -93470
rect -146 -96082 -112 -94906
rect 112 -96082 146 -94906
rect -146 -97518 -112 -96342
rect 112 -97518 146 -96342
rect -146 -98954 -112 -97778
rect 112 -98954 146 -97778
rect -146 -100390 -112 -99214
rect 112 -100390 146 -99214
rect -146 -101826 -112 -100650
rect 112 -101826 146 -100650
rect -146 -103262 -112 -102086
rect 112 -103262 146 -102086
rect -146 -104698 -112 -103522
rect 112 -104698 146 -103522
rect -146 -106134 -112 -104958
rect 112 -106134 146 -104958
rect -146 -107570 -112 -106394
rect 112 -107570 146 -106394
rect -146 -109006 -112 -107830
rect 112 -109006 146 -107830
rect -146 -110442 -112 -109266
rect 112 -110442 146 -109266
rect -146 -111878 -112 -110702
rect 112 -111878 146 -110702
rect -146 -113314 -112 -112138
rect 112 -113314 146 -112138
rect -146 -114750 -112 -113574
rect 112 -114750 146 -113574
rect -146 -116186 -112 -115010
rect 112 -116186 146 -115010
rect -146 -117622 -112 -116446
rect 112 -117622 146 -116446
rect -146 -119058 -112 -117882
rect 112 -119058 146 -117882
rect -146 -120494 -112 -119318
rect 112 -120494 146 -119318
rect -146 -121930 -112 -120754
rect 112 -121930 146 -120754
rect -146 -123366 -112 -122190
rect 112 -123366 146 -122190
rect -146 -124802 -112 -123626
rect 112 -124802 146 -123626
rect -146 -126238 -112 -125062
rect 112 -126238 146 -125062
rect -146 -127674 -112 -126498
rect 112 -127674 146 -126498
rect -146 -129110 -112 -127934
rect 112 -129110 146 -127934
rect -146 -130546 -112 -129370
rect 112 -130546 146 -129370
rect -146 -131982 -112 -130806
rect 112 -131982 146 -130806
rect -146 -133418 -112 -132242
rect 112 -133418 146 -132242
rect -146 -134854 -112 -133678
rect 112 -134854 146 -133678
rect -146 -136290 -112 -135114
rect 112 -136290 146 -135114
rect -146 -137726 -112 -136550
rect 112 -137726 146 -136550
rect -146 -139162 -112 -137986
rect 112 -139162 146 -137986
rect -146 -140598 -112 -139422
rect 112 -140598 146 -139422
rect -146 -142034 -112 -140858
rect 112 -142034 146 -140858
rect -146 -143470 -112 -142294
rect 112 -143470 146 -142294
rect -146 -144906 -112 -143730
rect 112 -144906 146 -143730
rect -146 -146342 -112 -145166
rect 112 -146342 146 -145166
rect -146 -147778 -112 -146602
rect 112 -147778 146 -146602
rect -146 -149214 -112 -148038
rect 112 -149214 146 -148038
rect -146 -150650 -112 -149474
rect 112 -150650 146 -149474
rect -146 -152086 -112 -150910
rect 112 -152086 146 -150910
rect -146 -153522 -112 -152346
rect 112 -153522 146 -152346
rect -146 -154958 -112 -153782
rect 112 -154958 146 -153782
rect -146 -156394 -112 -155218
rect 112 -156394 146 -155218
rect -146 -157830 -112 -156654
rect 112 -157830 146 -156654
rect -146 -159266 -112 -158090
rect 112 -159266 146 -158090
rect -146 -160702 -112 -159526
rect 112 -160702 146 -159526
rect -146 -162138 -112 -160962
rect 112 -162138 146 -160962
rect -146 -163574 -112 -162398
rect 112 -163574 146 -162398
rect -146 -165010 -112 -163834
rect 112 -165010 146 -163834
rect -146 -166446 -112 -165270
rect 112 -166446 146 -165270
rect -146 -167882 -112 -166706
rect 112 -167882 146 -166706
rect -146 -169318 -112 -168142
rect 112 -169318 146 -168142
rect -146 -170754 -112 -169578
rect 112 -170754 146 -169578
rect -146 -172190 -112 -171014
rect 112 -172190 146 -171014
rect -146 -173626 -112 -172450
rect 112 -173626 146 -172450
rect -146 -175062 -112 -173886
rect 112 -175062 146 -173886
rect -146 -176498 -112 -175322
rect 112 -176498 146 -175322
rect -146 -177934 -112 -176758
rect 112 -177934 146 -176758
rect -146 -179370 -112 -178194
rect 112 -179370 146 -178194
rect -146 -180806 -112 -179630
rect 112 -180806 146 -179630
rect -146 -182242 -112 -181066
rect 112 -182242 146 -181066
rect -146 -183678 -112 -182502
rect 112 -183678 146 -182502
<< mvnsubdiff >>
rect -292 183909 292 183921
rect -292 183875 -184 183909
rect 184 183875 292 183909
rect -292 183863 292 183875
rect -292 183813 -234 183863
rect -292 -183813 -280 183813
rect -246 -183813 -234 183813
rect 234 183813 292 183863
rect -292 -183863 -234 -183813
rect 234 -183813 246 183813
rect 280 -183813 292 183813
rect 234 -183863 292 -183813
rect -292 -183875 292 -183863
rect -292 -183909 -184 -183875
rect 184 -183909 292 -183875
rect -292 -183921 292 -183909
<< mvnsubdiffcont >>
rect -184 183875 184 183909
rect -280 -183813 -246 183813
rect 246 -183813 280 183813
rect -184 -183909 184 -183875
<< poly >>
rect -100 183771 100 183787
rect -100 183737 -84 183771
rect 84 183737 100 183771
rect -100 183690 100 183737
rect -100 182443 100 182490
rect -100 182409 -84 182443
rect 84 182409 100 182443
rect -100 182393 100 182409
rect -100 182335 100 182351
rect -100 182301 -84 182335
rect 84 182301 100 182335
rect -100 182254 100 182301
rect -100 181007 100 181054
rect -100 180973 -84 181007
rect 84 180973 100 181007
rect -100 180957 100 180973
rect -100 180899 100 180915
rect -100 180865 -84 180899
rect 84 180865 100 180899
rect -100 180818 100 180865
rect -100 179571 100 179618
rect -100 179537 -84 179571
rect 84 179537 100 179571
rect -100 179521 100 179537
rect -100 179463 100 179479
rect -100 179429 -84 179463
rect 84 179429 100 179463
rect -100 179382 100 179429
rect -100 178135 100 178182
rect -100 178101 -84 178135
rect 84 178101 100 178135
rect -100 178085 100 178101
rect -100 178027 100 178043
rect -100 177993 -84 178027
rect 84 177993 100 178027
rect -100 177946 100 177993
rect -100 176699 100 176746
rect -100 176665 -84 176699
rect 84 176665 100 176699
rect -100 176649 100 176665
rect -100 176591 100 176607
rect -100 176557 -84 176591
rect 84 176557 100 176591
rect -100 176510 100 176557
rect -100 175263 100 175310
rect -100 175229 -84 175263
rect 84 175229 100 175263
rect -100 175213 100 175229
rect -100 175155 100 175171
rect -100 175121 -84 175155
rect 84 175121 100 175155
rect -100 175074 100 175121
rect -100 173827 100 173874
rect -100 173793 -84 173827
rect 84 173793 100 173827
rect -100 173777 100 173793
rect -100 173719 100 173735
rect -100 173685 -84 173719
rect 84 173685 100 173719
rect -100 173638 100 173685
rect -100 172391 100 172438
rect -100 172357 -84 172391
rect 84 172357 100 172391
rect -100 172341 100 172357
rect -100 172283 100 172299
rect -100 172249 -84 172283
rect 84 172249 100 172283
rect -100 172202 100 172249
rect -100 170955 100 171002
rect -100 170921 -84 170955
rect 84 170921 100 170955
rect -100 170905 100 170921
rect -100 170847 100 170863
rect -100 170813 -84 170847
rect 84 170813 100 170847
rect -100 170766 100 170813
rect -100 169519 100 169566
rect -100 169485 -84 169519
rect 84 169485 100 169519
rect -100 169469 100 169485
rect -100 169411 100 169427
rect -100 169377 -84 169411
rect 84 169377 100 169411
rect -100 169330 100 169377
rect -100 168083 100 168130
rect -100 168049 -84 168083
rect 84 168049 100 168083
rect -100 168033 100 168049
rect -100 167975 100 167991
rect -100 167941 -84 167975
rect 84 167941 100 167975
rect -100 167894 100 167941
rect -100 166647 100 166694
rect -100 166613 -84 166647
rect 84 166613 100 166647
rect -100 166597 100 166613
rect -100 166539 100 166555
rect -100 166505 -84 166539
rect 84 166505 100 166539
rect -100 166458 100 166505
rect -100 165211 100 165258
rect -100 165177 -84 165211
rect 84 165177 100 165211
rect -100 165161 100 165177
rect -100 165103 100 165119
rect -100 165069 -84 165103
rect 84 165069 100 165103
rect -100 165022 100 165069
rect -100 163775 100 163822
rect -100 163741 -84 163775
rect 84 163741 100 163775
rect -100 163725 100 163741
rect -100 163667 100 163683
rect -100 163633 -84 163667
rect 84 163633 100 163667
rect -100 163586 100 163633
rect -100 162339 100 162386
rect -100 162305 -84 162339
rect 84 162305 100 162339
rect -100 162289 100 162305
rect -100 162231 100 162247
rect -100 162197 -84 162231
rect 84 162197 100 162231
rect -100 162150 100 162197
rect -100 160903 100 160950
rect -100 160869 -84 160903
rect 84 160869 100 160903
rect -100 160853 100 160869
rect -100 160795 100 160811
rect -100 160761 -84 160795
rect 84 160761 100 160795
rect -100 160714 100 160761
rect -100 159467 100 159514
rect -100 159433 -84 159467
rect 84 159433 100 159467
rect -100 159417 100 159433
rect -100 159359 100 159375
rect -100 159325 -84 159359
rect 84 159325 100 159359
rect -100 159278 100 159325
rect -100 158031 100 158078
rect -100 157997 -84 158031
rect 84 157997 100 158031
rect -100 157981 100 157997
rect -100 157923 100 157939
rect -100 157889 -84 157923
rect 84 157889 100 157923
rect -100 157842 100 157889
rect -100 156595 100 156642
rect -100 156561 -84 156595
rect 84 156561 100 156595
rect -100 156545 100 156561
rect -100 156487 100 156503
rect -100 156453 -84 156487
rect 84 156453 100 156487
rect -100 156406 100 156453
rect -100 155159 100 155206
rect -100 155125 -84 155159
rect 84 155125 100 155159
rect -100 155109 100 155125
rect -100 155051 100 155067
rect -100 155017 -84 155051
rect 84 155017 100 155051
rect -100 154970 100 155017
rect -100 153723 100 153770
rect -100 153689 -84 153723
rect 84 153689 100 153723
rect -100 153673 100 153689
rect -100 153615 100 153631
rect -100 153581 -84 153615
rect 84 153581 100 153615
rect -100 153534 100 153581
rect -100 152287 100 152334
rect -100 152253 -84 152287
rect 84 152253 100 152287
rect -100 152237 100 152253
rect -100 152179 100 152195
rect -100 152145 -84 152179
rect 84 152145 100 152179
rect -100 152098 100 152145
rect -100 150851 100 150898
rect -100 150817 -84 150851
rect 84 150817 100 150851
rect -100 150801 100 150817
rect -100 150743 100 150759
rect -100 150709 -84 150743
rect 84 150709 100 150743
rect -100 150662 100 150709
rect -100 149415 100 149462
rect -100 149381 -84 149415
rect 84 149381 100 149415
rect -100 149365 100 149381
rect -100 149307 100 149323
rect -100 149273 -84 149307
rect 84 149273 100 149307
rect -100 149226 100 149273
rect -100 147979 100 148026
rect -100 147945 -84 147979
rect 84 147945 100 147979
rect -100 147929 100 147945
rect -100 147871 100 147887
rect -100 147837 -84 147871
rect 84 147837 100 147871
rect -100 147790 100 147837
rect -100 146543 100 146590
rect -100 146509 -84 146543
rect 84 146509 100 146543
rect -100 146493 100 146509
rect -100 146435 100 146451
rect -100 146401 -84 146435
rect 84 146401 100 146435
rect -100 146354 100 146401
rect -100 145107 100 145154
rect -100 145073 -84 145107
rect 84 145073 100 145107
rect -100 145057 100 145073
rect -100 144999 100 145015
rect -100 144965 -84 144999
rect 84 144965 100 144999
rect -100 144918 100 144965
rect -100 143671 100 143718
rect -100 143637 -84 143671
rect 84 143637 100 143671
rect -100 143621 100 143637
rect -100 143563 100 143579
rect -100 143529 -84 143563
rect 84 143529 100 143563
rect -100 143482 100 143529
rect -100 142235 100 142282
rect -100 142201 -84 142235
rect 84 142201 100 142235
rect -100 142185 100 142201
rect -100 142127 100 142143
rect -100 142093 -84 142127
rect 84 142093 100 142127
rect -100 142046 100 142093
rect -100 140799 100 140846
rect -100 140765 -84 140799
rect 84 140765 100 140799
rect -100 140749 100 140765
rect -100 140691 100 140707
rect -100 140657 -84 140691
rect 84 140657 100 140691
rect -100 140610 100 140657
rect -100 139363 100 139410
rect -100 139329 -84 139363
rect 84 139329 100 139363
rect -100 139313 100 139329
rect -100 139255 100 139271
rect -100 139221 -84 139255
rect 84 139221 100 139255
rect -100 139174 100 139221
rect -100 137927 100 137974
rect -100 137893 -84 137927
rect 84 137893 100 137927
rect -100 137877 100 137893
rect -100 137819 100 137835
rect -100 137785 -84 137819
rect 84 137785 100 137819
rect -100 137738 100 137785
rect -100 136491 100 136538
rect -100 136457 -84 136491
rect 84 136457 100 136491
rect -100 136441 100 136457
rect -100 136383 100 136399
rect -100 136349 -84 136383
rect 84 136349 100 136383
rect -100 136302 100 136349
rect -100 135055 100 135102
rect -100 135021 -84 135055
rect 84 135021 100 135055
rect -100 135005 100 135021
rect -100 134947 100 134963
rect -100 134913 -84 134947
rect 84 134913 100 134947
rect -100 134866 100 134913
rect -100 133619 100 133666
rect -100 133585 -84 133619
rect 84 133585 100 133619
rect -100 133569 100 133585
rect -100 133511 100 133527
rect -100 133477 -84 133511
rect 84 133477 100 133511
rect -100 133430 100 133477
rect -100 132183 100 132230
rect -100 132149 -84 132183
rect 84 132149 100 132183
rect -100 132133 100 132149
rect -100 132075 100 132091
rect -100 132041 -84 132075
rect 84 132041 100 132075
rect -100 131994 100 132041
rect -100 130747 100 130794
rect -100 130713 -84 130747
rect 84 130713 100 130747
rect -100 130697 100 130713
rect -100 130639 100 130655
rect -100 130605 -84 130639
rect 84 130605 100 130639
rect -100 130558 100 130605
rect -100 129311 100 129358
rect -100 129277 -84 129311
rect 84 129277 100 129311
rect -100 129261 100 129277
rect -100 129203 100 129219
rect -100 129169 -84 129203
rect 84 129169 100 129203
rect -100 129122 100 129169
rect -100 127875 100 127922
rect -100 127841 -84 127875
rect 84 127841 100 127875
rect -100 127825 100 127841
rect -100 127767 100 127783
rect -100 127733 -84 127767
rect 84 127733 100 127767
rect -100 127686 100 127733
rect -100 126439 100 126486
rect -100 126405 -84 126439
rect 84 126405 100 126439
rect -100 126389 100 126405
rect -100 126331 100 126347
rect -100 126297 -84 126331
rect 84 126297 100 126331
rect -100 126250 100 126297
rect -100 125003 100 125050
rect -100 124969 -84 125003
rect 84 124969 100 125003
rect -100 124953 100 124969
rect -100 124895 100 124911
rect -100 124861 -84 124895
rect 84 124861 100 124895
rect -100 124814 100 124861
rect -100 123567 100 123614
rect -100 123533 -84 123567
rect 84 123533 100 123567
rect -100 123517 100 123533
rect -100 123459 100 123475
rect -100 123425 -84 123459
rect 84 123425 100 123459
rect -100 123378 100 123425
rect -100 122131 100 122178
rect -100 122097 -84 122131
rect 84 122097 100 122131
rect -100 122081 100 122097
rect -100 122023 100 122039
rect -100 121989 -84 122023
rect 84 121989 100 122023
rect -100 121942 100 121989
rect -100 120695 100 120742
rect -100 120661 -84 120695
rect 84 120661 100 120695
rect -100 120645 100 120661
rect -100 120587 100 120603
rect -100 120553 -84 120587
rect 84 120553 100 120587
rect -100 120506 100 120553
rect -100 119259 100 119306
rect -100 119225 -84 119259
rect 84 119225 100 119259
rect -100 119209 100 119225
rect -100 119151 100 119167
rect -100 119117 -84 119151
rect 84 119117 100 119151
rect -100 119070 100 119117
rect -100 117823 100 117870
rect -100 117789 -84 117823
rect 84 117789 100 117823
rect -100 117773 100 117789
rect -100 117715 100 117731
rect -100 117681 -84 117715
rect 84 117681 100 117715
rect -100 117634 100 117681
rect -100 116387 100 116434
rect -100 116353 -84 116387
rect 84 116353 100 116387
rect -100 116337 100 116353
rect -100 116279 100 116295
rect -100 116245 -84 116279
rect 84 116245 100 116279
rect -100 116198 100 116245
rect -100 114951 100 114998
rect -100 114917 -84 114951
rect 84 114917 100 114951
rect -100 114901 100 114917
rect -100 114843 100 114859
rect -100 114809 -84 114843
rect 84 114809 100 114843
rect -100 114762 100 114809
rect -100 113515 100 113562
rect -100 113481 -84 113515
rect 84 113481 100 113515
rect -100 113465 100 113481
rect -100 113407 100 113423
rect -100 113373 -84 113407
rect 84 113373 100 113407
rect -100 113326 100 113373
rect -100 112079 100 112126
rect -100 112045 -84 112079
rect 84 112045 100 112079
rect -100 112029 100 112045
rect -100 111971 100 111987
rect -100 111937 -84 111971
rect 84 111937 100 111971
rect -100 111890 100 111937
rect -100 110643 100 110690
rect -100 110609 -84 110643
rect 84 110609 100 110643
rect -100 110593 100 110609
rect -100 110535 100 110551
rect -100 110501 -84 110535
rect 84 110501 100 110535
rect -100 110454 100 110501
rect -100 109207 100 109254
rect -100 109173 -84 109207
rect 84 109173 100 109207
rect -100 109157 100 109173
rect -100 109099 100 109115
rect -100 109065 -84 109099
rect 84 109065 100 109099
rect -100 109018 100 109065
rect -100 107771 100 107818
rect -100 107737 -84 107771
rect 84 107737 100 107771
rect -100 107721 100 107737
rect -100 107663 100 107679
rect -100 107629 -84 107663
rect 84 107629 100 107663
rect -100 107582 100 107629
rect -100 106335 100 106382
rect -100 106301 -84 106335
rect 84 106301 100 106335
rect -100 106285 100 106301
rect -100 106227 100 106243
rect -100 106193 -84 106227
rect 84 106193 100 106227
rect -100 106146 100 106193
rect -100 104899 100 104946
rect -100 104865 -84 104899
rect 84 104865 100 104899
rect -100 104849 100 104865
rect -100 104791 100 104807
rect -100 104757 -84 104791
rect 84 104757 100 104791
rect -100 104710 100 104757
rect -100 103463 100 103510
rect -100 103429 -84 103463
rect 84 103429 100 103463
rect -100 103413 100 103429
rect -100 103355 100 103371
rect -100 103321 -84 103355
rect 84 103321 100 103355
rect -100 103274 100 103321
rect -100 102027 100 102074
rect -100 101993 -84 102027
rect 84 101993 100 102027
rect -100 101977 100 101993
rect -100 101919 100 101935
rect -100 101885 -84 101919
rect 84 101885 100 101919
rect -100 101838 100 101885
rect -100 100591 100 100638
rect -100 100557 -84 100591
rect 84 100557 100 100591
rect -100 100541 100 100557
rect -100 100483 100 100499
rect -100 100449 -84 100483
rect 84 100449 100 100483
rect -100 100402 100 100449
rect -100 99155 100 99202
rect -100 99121 -84 99155
rect 84 99121 100 99155
rect -100 99105 100 99121
rect -100 99047 100 99063
rect -100 99013 -84 99047
rect 84 99013 100 99047
rect -100 98966 100 99013
rect -100 97719 100 97766
rect -100 97685 -84 97719
rect 84 97685 100 97719
rect -100 97669 100 97685
rect -100 97611 100 97627
rect -100 97577 -84 97611
rect 84 97577 100 97611
rect -100 97530 100 97577
rect -100 96283 100 96330
rect -100 96249 -84 96283
rect 84 96249 100 96283
rect -100 96233 100 96249
rect -100 96175 100 96191
rect -100 96141 -84 96175
rect 84 96141 100 96175
rect -100 96094 100 96141
rect -100 94847 100 94894
rect -100 94813 -84 94847
rect 84 94813 100 94847
rect -100 94797 100 94813
rect -100 94739 100 94755
rect -100 94705 -84 94739
rect 84 94705 100 94739
rect -100 94658 100 94705
rect -100 93411 100 93458
rect -100 93377 -84 93411
rect 84 93377 100 93411
rect -100 93361 100 93377
rect -100 93303 100 93319
rect -100 93269 -84 93303
rect 84 93269 100 93303
rect -100 93222 100 93269
rect -100 91975 100 92022
rect -100 91941 -84 91975
rect 84 91941 100 91975
rect -100 91925 100 91941
rect -100 91867 100 91883
rect -100 91833 -84 91867
rect 84 91833 100 91867
rect -100 91786 100 91833
rect -100 90539 100 90586
rect -100 90505 -84 90539
rect 84 90505 100 90539
rect -100 90489 100 90505
rect -100 90431 100 90447
rect -100 90397 -84 90431
rect 84 90397 100 90431
rect -100 90350 100 90397
rect -100 89103 100 89150
rect -100 89069 -84 89103
rect 84 89069 100 89103
rect -100 89053 100 89069
rect -100 88995 100 89011
rect -100 88961 -84 88995
rect 84 88961 100 88995
rect -100 88914 100 88961
rect -100 87667 100 87714
rect -100 87633 -84 87667
rect 84 87633 100 87667
rect -100 87617 100 87633
rect -100 87559 100 87575
rect -100 87525 -84 87559
rect 84 87525 100 87559
rect -100 87478 100 87525
rect -100 86231 100 86278
rect -100 86197 -84 86231
rect 84 86197 100 86231
rect -100 86181 100 86197
rect -100 86123 100 86139
rect -100 86089 -84 86123
rect 84 86089 100 86123
rect -100 86042 100 86089
rect -100 84795 100 84842
rect -100 84761 -84 84795
rect 84 84761 100 84795
rect -100 84745 100 84761
rect -100 84687 100 84703
rect -100 84653 -84 84687
rect 84 84653 100 84687
rect -100 84606 100 84653
rect -100 83359 100 83406
rect -100 83325 -84 83359
rect 84 83325 100 83359
rect -100 83309 100 83325
rect -100 83251 100 83267
rect -100 83217 -84 83251
rect 84 83217 100 83251
rect -100 83170 100 83217
rect -100 81923 100 81970
rect -100 81889 -84 81923
rect 84 81889 100 81923
rect -100 81873 100 81889
rect -100 81815 100 81831
rect -100 81781 -84 81815
rect 84 81781 100 81815
rect -100 81734 100 81781
rect -100 80487 100 80534
rect -100 80453 -84 80487
rect 84 80453 100 80487
rect -100 80437 100 80453
rect -100 80379 100 80395
rect -100 80345 -84 80379
rect 84 80345 100 80379
rect -100 80298 100 80345
rect -100 79051 100 79098
rect -100 79017 -84 79051
rect 84 79017 100 79051
rect -100 79001 100 79017
rect -100 78943 100 78959
rect -100 78909 -84 78943
rect 84 78909 100 78943
rect -100 78862 100 78909
rect -100 77615 100 77662
rect -100 77581 -84 77615
rect 84 77581 100 77615
rect -100 77565 100 77581
rect -100 77507 100 77523
rect -100 77473 -84 77507
rect 84 77473 100 77507
rect -100 77426 100 77473
rect -100 76179 100 76226
rect -100 76145 -84 76179
rect 84 76145 100 76179
rect -100 76129 100 76145
rect -100 76071 100 76087
rect -100 76037 -84 76071
rect 84 76037 100 76071
rect -100 75990 100 76037
rect -100 74743 100 74790
rect -100 74709 -84 74743
rect 84 74709 100 74743
rect -100 74693 100 74709
rect -100 74635 100 74651
rect -100 74601 -84 74635
rect 84 74601 100 74635
rect -100 74554 100 74601
rect -100 73307 100 73354
rect -100 73273 -84 73307
rect 84 73273 100 73307
rect -100 73257 100 73273
rect -100 73199 100 73215
rect -100 73165 -84 73199
rect 84 73165 100 73199
rect -100 73118 100 73165
rect -100 71871 100 71918
rect -100 71837 -84 71871
rect 84 71837 100 71871
rect -100 71821 100 71837
rect -100 71763 100 71779
rect -100 71729 -84 71763
rect 84 71729 100 71763
rect -100 71682 100 71729
rect -100 70435 100 70482
rect -100 70401 -84 70435
rect 84 70401 100 70435
rect -100 70385 100 70401
rect -100 70327 100 70343
rect -100 70293 -84 70327
rect 84 70293 100 70327
rect -100 70246 100 70293
rect -100 68999 100 69046
rect -100 68965 -84 68999
rect 84 68965 100 68999
rect -100 68949 100 68965
rect -100 68891 100 68907
rect -100 68857 -84 68891
rect 84 68857 100 68891
rect -100 68810 100 68857
rect -100 67563 100 67610
rect -100 67529 -84 67563
rect 84 67529 100 67563
rect -100 67513 100 67529
rect -100 67455 100 67471
rect -100 67421 -84 67455
rect 84 67421 100 67455
rect -100 67374 100 67421
rect -100 66127 100 66174
rect -100 66093 -84 66127
rect 84 66093 100 66127
rect -100 66077 100 66093
rect -100 66019 100 66035
rect -100 65985 -84 66019
rect 84 65985 100 66019
rect -100 65938 100 65985
rect -100 64691 100 64738
rect -100 64657 -84 64691
rect 84 64657 100 64691
rect -100 64641 100 64657
rect -100 64583 100 64599
rect -100 64549 -84 64583
rect 84 64549 100 64583
rect -100 64502 100 64549
rect -100 63255 100 63302
rect -100 63221 -84 63255
rect 84 63221 100 63255
rect -100 63205 100 63221
rect -100 63147 100 63163
rect -100 63113 -84 63147
rect 84 63113 100 63147
rect -100 63066 100 63113
rect -100 61819 100 61866
rect -100 61785 -84 61819
rect 84 61785 100 61819
rect -100 61769 100 61785
rect -100 61711 100 61727
rect -100 61677 -84 61711
rect 84 61677 100 61711
rect -100 61630 100 61677
rect -100 60383 100 60430
rect -100 60349 -84 60383
rect 84 60349 100 60383
rect -100 60333 100 60349
rect -100 60275 100 60291
rect -100 60241 -84 60275
rect 84 60241 100 60275
rect -100 60194 100 60241
rect -100 58947 100 58994
rect -100 58913 -84 58947
rect 84 58913 100 58947
rect -100 58897 100 58913
rect -100 58839 100 58855
rect -100 58805 -84 58839
rect 84 58805 100 58839
rect -100 58758 100 58805
rect -100 57511 100 57558
rect -100 57477 -84 57511
rect 84 57477 100 57511
rect -100 57461 100 57477
rect -100 57403 100 57419
rect -100 57369 -84 57403
rect 84 57369 100 57403
rect -100 57322 100 57369
rect -100 56075 100 56122
rect -100 56041 -84 56075
rect 84 56041 100 56075
rect -100 56025 100 56041
rect -100 55967 100 55983
rect -100 55933 -84 55967
rect 84 55933 100 55967
rect -100 55886 100 55933
rect -100 54639 100 54686
rect -100 54605 -84 54639
rect 84 54605 100 54639
rect -100 54589 100 54605
rect -100 54531 100 54547
rect -100 54497 -84 54531
rect 84 54497 100 54531
rect -100 54450 100 54497
rect -100 53203 100 53250
rect -100 53169 -84 53203
rect 84 53169 100 53203
rect -100 53153 100 53169
rect -100 53095 100 53111
rect -100 53061 -84 53095
rect 84 53061 100 53095
rect -100 53014 100 53061
rect -100 51767 100 51814
rect -100 51733 -84 51767
rect 84 51733 100 51767
rect -100 51717 100 51733
rect -100 51659 100 51675
rect -100 51625 -84 51659
rect 84 51625 100 51659
rect -100 51578 100 51625
rect -100 50331 100 50378
rect -100 50297 -84 50331
rect 84 50297 100 50331
rect -100 50281 100 50297
rect -100 50223 100 50239
rect -100 50189 -84 50223
rect 84 50189 100 50223
rect -100 50142 100 50189
rect -100 48895 100 48942
rect -100 48861 -84 48895
rect 84 48861 100 48895
rect -100 48845 100 48861
rect -100 48787 100 48803
rect -100 48753 -84 48787
rect 84 48753 100 48787
rect -100 48706 100 48753
rect -100 47459 100 47506
rect -100 47425 -84 47459
rect 84 47425 100 47459
rect -100 47409 100 47425
rect -100 47351 100 47367
rect -100 47317 -84 47351
rect 84 47317 100 47351
rect -100 47270 100 47317
rect -100 46023 100 46070
rect -100 45989 -84 46023
rect 84 45989 100 46023
rect -100 45973 100 45989
rect -100 45915 100 45931
rect -100 45881 -84 45915
rect 84 45881 100 45915
rect -100 45834 100 45881
rect -100 44587 100 44634
rect -100 44553 -84 44587
rect 84 44553 100 44587
rect -100 44537 100 44553
rect -100 44479 100 44495
rect -100 44445 -84 44479
rect 84 44445 100 44479
rect -100 44398 100 44445
rect -100 43151 100 43198
rect -100 43117 -84 43151
rect 84 43117 100 43151
rect -100 43101 100 43117
rect -100 43043 100 43059
rect -100 43009 -84 43043
rect 84 43009 100 43043
rect -100 42962 100 43009
rect -100 41715 100 41762
rect -100 41681 -84 41715
rect 84 41681 100 41715
rect -100 41665 100 41681
rect -100 41607 100 41623
rect -100 41573 -84 41607
rect 84 41573 100 41607
rect -100 41526 100 41573
rect -100 40279 100 40326
rect -100 40245 -84 40279
rect 84 40245 100 40279
rect -100 40229 100 40245
rect -100 40171 100 40187
rect -100 40137 -84 40171
rect 84 40137 100 40171
rect -100 40090 100 40137
rect -100 38843 100 38890
rect -100 38809 -84 38843
rect 84 38809 100 38843
rect -100 38793 100 38809
rect -100 38735 100 38751
rect -100 38701 -84 38735
rect 84 38701 100 38735
rect -100 38654 100 38701
rect -100 37407 100 37454
rect -100 37373 -84 37407
rect 84 37373 100 37407
rect -100 37357 100 37373
rect -100 37299 100 37315
rect -100 37265 -84 37299
rect 84 37265 100 37299
rect -100 37218 100 37265
rect -100 35971 100 36018
rect -100 35937 -84 35971
rect 84 35937 100 35971
rect -100 35921 100 35937
rect -100 35863 100 35879
rect -100 35829 -84 35863
rect 84 35829 100 35863
rect -100 35782 100 35829
rect -100 34535 100 34582
rect -100 34501 -84 34535
rect 84 34501 100 34535
rect -100 34485 100 34501
rect -100 34427 100 34443
rect -100 34393 -84 34427
rect 84 34393 100 34427
rect -100 34346 100 34393
rect -100 33099 100 33146
rect -100 33065 -84 33099
rect 84 33065 100 33099
rect -100 33049 100 33065
rect -100 32991 100 33007
rect -100 32957 -84 32991
rect 84 32957 100 32991
rect -100 32910 100 32957
rect -100 31663 100 31710
rect -100 31629 -84 31663
rect 84 31629 100 31663
rect -100 31613 100 31629
rect -100 31555 100 31571
rect -100 31521 -84 31555
rect 84 31521 100 31555
rect -100 31474 100 31521
rect -100 30227 100 30274
rect -100 30193 -84 30227
rect 84 30193 100 30227
rect -100 30177 100 30193
rect -100 30119 100 30135
rect -100 30085 -84 30119
rect 84 30085 100 30119
rect -100 30038 100 30085
rect -100 28791 100 28838
rect -100 28757 -84 28791
rect 84 28757 100 28791
rect -100 28741 100 28757
rect -100 28683 100 28699
rect -100 28649 -84 28683
rect 84 28649 100 28683
rect -100 28602 100 28649
rect -100 27355 100 27402
rect -100 27321 -84 27355
rect 84 27321 100 27355
rect -100 27305 100 27321
rect -100 27247 100 27263
rect -100 27213 -84 27247
rect 84 27213 100 27247
rect -100 27166 100 27213
rect -100 25919 100 25966
rect -100 25885 -84 25919
rect 84 25885 100 25919
rect -100 25869 100 25885
rect -100 25811 100 25827
rect -100 25777 -84 25811
rect 84 25777 100 25811
rect -100 25730 100 25777
rect -100 24483 100 24530
rect -100 24449 -84 24483
rect 84 24449 100 24483
rect -100 24433 100 24449
rect -100 24375 100 24391
rect -100 24341 -84 24375
rect 84 24341 100 24375
rect -100 24294 100 24341
rect -100 23047 100 23094
rect -100 23013 -84 23047
rect 84 23013 100 23047
rect -100 22997 100 23013
rect -100 22939 100 22955
rect -100 22905 -84 22939
rect 84 22905 100 22939
rect -100 22858 100 22905
rect -100 21611 100 21658
rect -100 21577 -84 21611
rect 84 21577 100 21611
rect -100 21561 100 21577
rect -100 21503 100 21519
rect -100 21469 -84 21503
rect 84 21469 100 21503
rect -100 21422 100 21469
rect -100 20175 100 20222
rect -100 20141 -84 20175
rect 84 20141 100 20175
rect -100 20125 100 20141
rect -100 20067 100 20083
rect -100 20033 -84 20067
rect 84 20033 100 20067
rect -100 19986 100 20033
rect -100 18739 100 18786
rect -100 18705 -84 18739
rect 84 18705 100 18739
rect -100 18689 100 18705
rect -100 18631 100 18647
rect -100 18597 -84 18631
rect 84 18597 100 18631
rect -100 18550 100 18597
rect -100 17303 100 17350
rect -100 17269 -84 17303
rect 84 17269 100 17303
rect -100 17253 100 17269
rect -100 17195 100 17211
rect -100 17161 -84 17195
rect 84 17161 100 17195
rect -100 17114 100 17161
rect -100 15867 100 15914
rect -100 15833 -84 15867
rect 84 15833 100 15867
rect -100 15817 100 15833
rect -100 15759 100 15775
rect -100 15725 -84 15759
rect 84 15725 100 15759
rect -100 15678 100 15725
rect -100 14431 100 14478
rect -100 14397 -84 14431
rect 84 14397 100 14431
rect -100 14381 100 14397
rect -100 14323 100 14339
rect -100 14289 -84 14323
rect 84 14289 100 14323
rect -100 14242 100 14289
rect -100 12995 100 13042
rect -100 12961 -84 12995
rect 84 12961 100 12995
rect -100 12945 100 12961
rect -100 12887 100 12903
rect -100 12853 -84 12887
rect 84 12853 100 12887
rect -100 12806 100 12853
rect -100 11559 100 11606
rect -100 11525 -84 11559
rect 84 11525 100 11559
rect -100 11509 100 11525
rect -100 11451 100 11467
rect -100 11417 -84 11451
rect 84 11417 100 11451
rect -100 11370 100 11417
rect -100 10123 100 10170
rect -100 10089 -84 10123
rect 84 10089 100 10123
rect -100 10073 100 10089
rect -100 10015 100 10031
rect -100 9981 -84 10015
rect 84 9981 100 10015
rect -100 9934 100 9981
rect -100 8687 100 8734
rect -100 8653 -84 8687
rect 84 8653 100 8687
rect -100 8637 100 8653
rect -100 8579 100 8595
rect -100 8545 -84 8579
rect 84 8545 100 8579
rect -100 8498 100 8545
rect -100 7251 100 7298
rect -100 7217 -84 7251
rect 84 7217 100 7251
rect -100 7201 100 7217
rect -100 7143 100 7159
rect -100 7109 -84 7143
rect 84 7109 100 7143
rect -100 7062 100 7109
rect -100 5815 100 5862
rect -100 5781 -84 5815
rect 84 5781 100 5815
rect -100 5765 100 5781
rect -100 5707 100 5723
rect -100 5673 -84 5707
rect 84 5673 100 5707
rect -100 5626 100 5673
rect -100 4379 100 4426
rect -100 4345 -84 4379
rect 84 4345 100 4379
rect -100 4329 100 4345
rect -100 4271 100 4287
rect -100 4237 -84 4271
rect 84 4237 100 4271
rect -100 4190 100 4237
rect -100 2943 100 2990
rect -100 2909 -84 2943
rect 84 2909 100 2943
rect -100 2893 100 2909
rect -100 2835 100 2851
rect -100 2801 -84 2835
rect 84 2801 100 2835
rect -100 2754 100 2801
rect -100 1507 100 1554
rect -100 1473 -84 1507
rect 84 1473 100 1507
rect -100 1457 100 1473
rect -100 1399 100 1415
rect -100 1365 -84 1399
rect 84 1365 100 1399
rect -100 1318 100 1365
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -1365 100 -1318
rect -100 -1399 -84 -1365
rect 84 -1399 100 -1365
rect -100 -1415 100 -1399
rect -100 -1473 100 -1457
rect -100 -1507 -84 -1473
rect 84 -1507 100 -1473
rect -100 -1554 100 -1507
rect -100 -2801 100 -2754
rect -100 -2835 -84 -2801
rect 84 -2835 100 -2801
rect -100 -2851 100 -2835
rect -100 -2909 100 -2893
rect -100 -2943 -84 -2909
rect 84 -2943 100 -2909
rect -100 -2990 100 -2943
rect -100 -4237 100 -4190
rect -100 -4271 -84 -4237
rect 84 -4271 100 -4237
rect -100 -4287 100 -4271
rect -100 -4345 100 -4329
rect -100 -4379 -84 -4345
rect 84 -4379 100 -4345
rect -100 -4426 100 -4379
rect -100 -5673 100 -5626
rect -100 -5707 -84 -5673
rect 84 -5707 100 -5673
rect -100 -5723 100 -5707
rect -100 -5781 100 -5765
rect -100 -5815 -84 -5781
rect 84 -5815 100 -5781
rect -100 -5862 100 -5815
rect -100 -7109 100 -7062
rect -100 -7143 -84 -7109
rect 84 -7143 100 -7109
rect -100 -7159 100 -7143
rect -100 -7217 100 -7201
rect -100 -7251 -84 -7217
rect 84 -7251 100 -7217
rect -100 -7298 100 -7251
rect -100 -8545 100 -8498
rect -100 -8579 -84 -8545
rect 84 -8579 100 -8545
rect -100 -8595 100 -8579
rect -100 -8653 100 -8637
rect -100 -8687 -84 -8653
rect 84 -8687 100 -8653
rect -100 -8734 100 -8687
rect -100 -9981 100 -9934
rect -100 -10015 -84 -9981
rect 84 -10015 100 -9981
rect -100 -10031 100 -10015
rect -100 -10089 100 -10073
rect -100 -10123 -84 -10089
rect 84 -10123 100 -10089
rect -100 -10170 100 -10123
rect -100 -11417 100 -11370
rect -100 -11451 -84 -11417
rect 84 -11451 100 -11417
rect -100 -11467 100 -11451
rect -100 -11525 100 -11509
rect -100 -11559 -84 -11525
rect 84 -11559 100 -11525
rect -100 -11606 100 -11559
rect -100 -12853 100 -12806
rect -100 -12887 -84 -12853
rect 84 -12887 100 -12853
rect -100 -12903 100 -12887
rect -100 -12961 100 -12945
rect -100 -12995 -84 -12961
rect 84 -12995 100 -12961
rect -100 -13042 100 -12995
rect -100 -14289 100 -14242
rect -100 -14323 -84 -14289
rect 84 -14323 100 -14289
rect -100 -14339 100 -14323
rect -100 -14397 100 -14381
rect -100 -14431 -84 -14397
rect 84 -14431 100 -14397
rect -100 -14478 100 -14431
rect -100 -15725 100 -15678
rect -100 -15759 -84 -15725
rect 84 -15759 100 -15725
rect -100 -15775 100 -15759
rect -100 -15833 100 -15817
rect -100 -15867 -84 -15833
rect 84 -15867 100 -15833
rect -100 -15914 100 -15867
rect -100 -17161 100 -17114
rect -100 -17195 -84 -17161
rect 84 -17195 100 -17161
rect -100 -17211 100 -17195
rect -100 -17269 100 -17253
rect -100 -17303 -84 -17269
rect 84 -17303 100 -17269
rect -100 -17350 100 -17303
rect -100 -18597 100 -18550
rect -100 -18631 -84 -18597
rect 84 -18631 100 -18597
rect -100 -18647 100 -18631
rect -100 -18705 100 -18689
rect -100 -18739 -84 -18705
rect 84 -18739 100 -18705
rect -100 -18786 100 -18739
rect -100 -20033 100 -19986
rect -100 -20067 -84 -20033
rect 84 -20067 100 -20033
rect -100 -20083 100 -20067
rect -100 -20141 100 -20125
rect -100 -20175 -84 -20141
rect 84 -20175 100 -20141
rect -100 -20222 100 -20175
rect -100 -21469 100 -21422
rect -100 -21503 -84 -21469
rect 84 -21503 100 -21469
rect -100 -21519 100 -21503
rect -100 -21577 100 -21561
rect -100 -21611 -84 -21577
rect 84 -21611 100 -21577
rect -100 -21658 100 -21611
rect -100 -22905 100 -22858
rect -100 -22939 -84 -22905
rect 84 -22939 100 -22905
rect -100 -22955 100 -22939
rect -100 -23013 100 -22997
rect -100 -23047 -84 -23013
rect 84 -23047 100 -23013
rect -100 -23094 100 -23047
rect -100 -24341 100 -24294
rect -100 -24375 -84 -24341
rect 84 -24375 100 -24341
rect -100 -24391 100 -24375
rect -100 -24449 100 -24433
rect -100 -24483 -84 -24449
rect 84 -24483 100 -24449
rect -100 -24530 100 -24483
rect -100 -25777 100 -25730
rect -100 -25811 -84 -25777
rect 84 -25811 100 -25777
rect -100 -25827 100 -25811
rect -100 -25885 100 -25869
rect -100 -25919 -84 -25885
rect 84 -25919 100 -25885
rect -100 -25966 100 -25919
rect -100 -27213 100 -27166
rect -100 -27247 -84 -27213
rect 84 -27247 100 -27213
rect -100 -27263 100 -27247
rect -100 -27321 100 -27305
rect -100 -27355 -84 -27321
rect 84 -27355 100 -27321
rect -100 -27402 100 -27355
rect -100 -28649 100 -28602
rect -100 -28683 -84 -28649
rect 84 -28683 100 -28649
rect -100 -28699 100 -28683
rect -100 -28757 100 -28741
rect -100 -28791 -84 -28757
rect 84 -28791 100 -28757
rect -100 -28838 100 -28791
rect -100 -30085 100 -30038
rect -100 -30119 -84 -30085
rect 84 -30119 100 -30085
rect -100 -30135 100 -30119
rect -100 -30193 100 -30177
rect -100 -30227 -84 -30193
rect 84 -30227 100 -30193
rect -100 -30274 100 -30227
rect -100 -31521 100 -31474
rect -100 -31555 -84 -31521
rect 84 -31555 100 -31521
rect -100 -31571 100 -31555
rect -100 -31629 100 -31613
rect -100 -31663 -84 -31629
rect 84 -31663 100 -31629
rect -100 -31710 100 -31663
rect -100 -32957 100 -32910
rect -100 -32991 -84 -32957
rect 84 -32991 100 -32957
rect -100 -33007 100 -32991
rect -100 -33065 100 -33049
rect -100 -33099 -84 -33065
rect 84 -33099 100 -33065
rect -100 -33146 100 -33099
rect -100 -34393 100 -34346
rect -100 -34427 -84 -34393
rect 84 -34427 100 -34393
rect -100 -34443 100 -34427
rect -100 -34501 100 -34485
rect -100 -34535 -84 -34501
rect 84 -34535 100 -34501
rect -100 -34582 100 -34535
rect -100 -35829 100 -35782
rect -100 -35863 -84 -35829
rect 84 -35863 100 -35829
rect -100 -35879 100 -35863
rect -100 -35937 100 -35921
rect -100 -35971 -84 -35937
rect 84 -35971 100 -35937
rect -100 -36018 100 -35971
rect -100 -37265 100 -37218
rect -100 -37299 -84 -37265
rect 84 -37299 100 -37265
rect -100 -37315 100 -37299
rect -100 -37373 100 -37357
rect -100 -37407 -84 -37373
rect 84 -37407 100 -37373
rect -100 -37454 100 -37407
rect -100 -38701 100 -38654
rect -100 -38735 -84 -38701
rect 84 -38735 100 -38701
rect -100 -38751 100 -38735
rect -100 -38809 100 -38793
rect -100 -38843 -84 -38809
rect 84 -38843 100 -38809
rect -100 -38890 100 -38843
rect -100 -40137 100 -40090
rect -100 -40171 -84 -40137
rect 84 -40171 100 -40137
rect -100 -40187 100 -40171
rect -100 -40245 100 -40229
rect -100 -40279 -84 -40245
rect 84 -40279 100 -40245
rect -100 -40326 100 -40279
rect -100 -41573 100 -41526
rect -100 -41607 -84 -41573
rect 84 -41607 100 -41573
rect -100 -41623 100 -41607
rect -100 -41681 100 -41665
rect -100 -41715 -84 -41681
rect 84 -41715 100 -41681
rect -100 -41762 100 -41715
rect -100 -43009 100 -42962
rect -100 -43043 -84 -43009
rect 84 -43043 100 -43009
rect -100 -43059 100 -43043
rect -100 -43117 100 -43101
rect -100 -43151 -84 -43117
rect 84 -43151 100 -43117
rect -100 -43198 100 -43151
rect -100 -44445 100 -44398
rect -100 -44479 -84 -44445
rect 84 -44479 100 -44445
rect -100 -44495 100 -44479
rect -100 -44553 100 -44537
rect -100 -44587 -84 -44553
rect 84 -44587 100 -44553
rect -100 -44634 100 -44587
rect -100 -45881 100 -45834
rect -100 -45915 -84 -45881
rect 84 -45915 100 -45881
rect -100 -45931 100 -45915
rect -100 -45989 100 -45973
rect -100 -46023 -84 -45989
rect 84 -46023 100 -45989
rect -100 -46070 100 -46023
rect -100 -47317 100 -47270
rect -100 -47351 -84 -47317
rect 84 -47351 100 -47317
rect -100 -47367 100 -47351
rect -100 -47425 100 -47409
rect -100 -47459 -84 -47425
rect 84 -47459 100 -47425
rect -100 -47506 100 -47459
rect -100 -48753 100 -48706
rect -100 -48787 -84 -48753
rect 84 -48787 100 -48753
rect -100 -48803 100 -48787
rect -100 -48861 100 -48845
rect -100 -48895 -84 -48861
rect 84 -48895 100 -48861
rect -100 -48942 100 -48895
rect -100 -50189 100 -50142
rect -100 -50223 -84 -50189
rect 84 -50223 100 -50189
rect -100 -50239 100 -50223
rect -100 -50297 100 -50281
rect -100 -50331 -84 -50297
rect 84 -50331 100 -50297
rect -100 -50378 100 -50331
rect -100 -51625 100 -51578
rect -100 -51659 -84 -51625
rect 84 -51659 100 -51625
rect -100 -51675 100 -51659
rect -100 -51733 100 -51717
rect -100 -51767 -84 -51733
rect 84 -51767 100 -51733
rect -100 -51814 100 -51767
rect -100 -53061 100 -53014
rect -100 -53095 -84 -53061
rect 84 -53095 100 -53061
rect -100 -53111 100 -53095
rect -100 -53169 100 -53153
rect -100 -53203 -84 -53169
rect 84 -53203 100 -53169
rect -100 -53250 100 -53203
rect -100 -54497 100 -54450
rect -100 -54531 -84 -54497
rect 84 -54531 100 -54497
rect -100 -54547 100 -54531
rect -100 -54605 100 -54589
rect -100 -54639 -84 -54605
rect 84 -54639 100 -54605
rect -100 -54686 100 -54639
rect -100 -55933 100 -55886
rect -100 -55967 -84 -55933
rect 84 -55967 100 -55933
rect -100 -55983 100 -55967
rect -100 -56041 100 -56025
rect -100 -56075 -84 -56041
rect 84 -56075 100 -56041
rect -100 -56122 100 -56075
rect -100 -57369 100 -57322
rect -100 -57403 -84 -57369
rect 84 -57403 100 -57369
rect -100 -57419 100 -57403
rect -100 -57477 100 -57461
rect -100 -57511 -84 -57477
rect 84 -57511 100 -57477
rect -100 -57558 100 -57511
rect -100 -58805 100 -58758
rect -100 -58839 -84 -58805
rect 84 -58839 100 -58805
rect -100 -58855 100 -58839
rect -100 -58913 100 -58897
rect -100 -58947 -84 -58913
rect 84 -58947 100 -58913
rect -100 -58994 100 -58947
rect -100 -60241 100 -60194
rect -100 -60275 -84 -60241
rect 84 -60275 100 -60241
rect -100 -60291 100 -60275
rect -100 -60349 100 -60333
rect -100 -60383 -84 -60349
rect 84 -60383 100 -60349
rect -100 -60430 100 -60383
rect -100 -61677 100 -61630
rect -100 -61711 -84 -61677
rect 84 -61711 100 -61677
rect -100 -61727 100 -61711
rect -100 -61785 100 -61769
rect -100 -61819 -84 -61785
rect 84 -61819 100 -61785
rect -100 -61866 100 -61819
rect -100 -63113 100 -63066
rect -100 -63147 -84 -63113
rect 84 -63147 100 -63113
rect -100 -63163 100 -63147
rect -100 -63221 100 -63205
rect -100 -63255 -84 -63221
rect 84 -63255 100 -63221
rect -100 -63302 100 -63255
rect -100 -64549 100 -64502
rect -100 -64583 -84 -64549
rect 84 -64583 100 -64549
rect -100 -64599 100 -64583
rect -100 -64657 100 -64641
rect -100 -64691 -84 -64657
rect 84 -64691 100 -64657
rect -100 -64738 100 -64691
rect -100 -65985 100 -65938
rect -100 -66019 -84 -65985
rect 84 -66019 100 -65985
rect -100 -66035 100 -66019
rect -100 -66093 100 -66077
rect -100 -66127 -84 -66093
rect 84 -66127 100 -66093
rect -100 -66174 100 -66127
rect -100 -67421 100 -67374
rect -100 -67455 -84 -67421
rect 84 -67455 100 -67421
rect -100 -67471 100 -67455
rect -100 -67529 100 -67513
rect -100 -67563 -84 -67529
rect 84 -67563 100 -67529
rect -100 -67610 100 -67563
rect -100 -68857 100 -68810
rect -100 -68891 -84 -68857
rect 84 -68891 100 -68857
rect -100 -68907 100 -68891
rect -100 -68965 100 -68949
rect -100 -68999 -84 -68965
rect 84 -68999 100 -68965
rect -100 -69046 100 -68999
rect -100 -70293 100 -70246
rect -100 -70327 -84 -70293
rect 84 -70327 100 -70293
rect -100 -70343 100 -70327
rect -100 -70401 100 -70385
rect -100 -70435 -84 -70401
rect 84 -70435 100 -70401
rect -100 -70482 100 -70435
rect -100 -71729 100 -71682
rect -100 -71763 -84 -71729
rect 84 -71763 100 -71729
rect -100 -71779 100 -71763
rect -100 -71837 100 -71821
rect -100 -71871 -84 -71837
rect 84 -71871 100 -71837
rect -100 -71918 100 -71871
rect -100 -73165 100 -73118
rect -100 -73199 -84 -73165
rect 84 -73199 100 -73165
rect -100 -73215 100 -73199
rect -100 -73273 100 -73257
rect -100 -73307 -84 -73273
rect 84 -73307 100 -73273
rect -100 -73354 100 -73307
rect -100 -74601 100 -74554
rect -100 -74635 -84 -74601
rect 84 -74635 100 -74601
rect -100 -74651 100 -74635
rect -100 -74709 100 -74693
rect -100 -74743 -84 -74709
rect 84 -74743 100 -74709
rect -100 -74790 100 -74743
rect -100 -76037 100 -75990
rect -100 -76071 -84 -76037
rect 84 -76071 100 -76037
rect -100 -76087 100 -76071
rect -100 -76145 100 -76129
rect -100 -76179 -84 -76145
rect 84 -76179 100 -76145
rect -100 -76226 100 -76179
rect -100 -77473 100 -77426
rect -100 -77507 -84 -77473
rect 84 -77507 100 -77473
rect -100 -77523 100 -77507
rect -100 -77581 100 -77565
rect -100 -77615 -84 -77581
rect 84 -77615 100 -77581
rect -100 -77662 100 -77615
rect -100 -78909 100 -78862
rect -100 -78943 -84 -78909
rect 84 -78943 100 -78909
rect -100 -78959 100 -78943
rect -100 -79017 100 -79001
rect -100 -79051 -84 -79017
rect 84 -79051 100 -79017
rect -100 -79098 100 -79051
rect -100 -80345 100 -80298
rect -100 -80379 -84 -80345
rect 84 -80379 100 -80345
rect -100 -80395 100 -80379
rect -100 -80453 100 -80437
rect -100 -80487 -84 -80453
rect 84 -80487 100 -80453
rect -100 -80534 100 -80487
rect -100 -81781 100 -81734
rect -100 -81815 -84 -81781
rect 84 -81815 100 -81781
rect -100 -81831 100 -81815
rect -100 -81889 100 -81873
rect -100 -81923 -84 -81889
rect 84 -81923 100 -81889
rect -100 -81970 100 -81923
rect -100 -83217 100 -83170
rect -100 -83251 -84 -83217
rect 84 -83251 100 -83217
rect -100 -83267 100 -83251
rect -100 -83325 100 -83309
rect -100 -83359 -84 -83325
rect 84 -83359 100 -83325
rect -100 -83406 100 -83359
rect -100 -84653 100 -84606
rect -100 -84687 -84 -84653
rect 84 -84687 100 -84653
rect -100 -84703 100 -84687
rect -100 -84761 100 -84745
rect -100 -84795 -84 -84761
rect 84 -84795 100 -84761
rect -100 -84842 100 -84795
rect -100 -86089 100 -86042
rect -100 -86123 -84 -86089
rect 84 -86123 100 -86089
rect -100 -86139 100 -86123
rect -100 -86197 100 -86181
rect -100 -86231 -84 -86197
rect 84 -86231 100 -86197
rect -100 -86278 100 -86231
rect -100 -87525 100 -87478
rect -100 -87559 -84 -87525
rect 84 -87559 100 -87525
rect -100 -87575 100 -87559
rect -100 -87633 100 -87617
rect -100 -87667 -84 -87633
rect 84 -87667 100 -87633
rect -100 -87714 100 -87667
rect -100 -88961 100 -88914
rect -100 -88995 -84 -88961
rect 84 -88995 100 -88961
rect -100 -89011 100 -88995
rect -100 -89069 100 -89053
rect -100 -89103 -84 -89069
rect 84 -89103 100 -89069
rect -100 -89150 100 -89103
rect -100 -90397 100 -90350
rect -100 -90431 -84 -90397
rect 84 -90431 100 -90397
rect -100 -90447 100 -90431
rect -100 -90505 100 -90489
rect -100 -90539 -84 -90505
rect 84 -90539 100 -90505
rect -100 -90586 100 -90539
rect -100 -91833 100 -91786
rect -100 -91867 -84 -91833
rect 84 -91867 100 -91833
rect -100 -91883 100 -91867
rect -100 -91941 100 -91925
rect -100 -91975 -84 -91941
rect 84 -91975 100 -91941
rect -100 -92022 100 -91975
rect -100 -93269 100 -93222
rect -100 -93303 -84 -93269
rect 84 -93303 100 -93269
rect -100 -93319 100 -93303
rect -100 -93377 100 -93361
rect -100 -93411 -84 -93377
rect 84 -93411 100 -93377
rect -100 -93458 100 -93411
rect -100 -94705 100 -94658
rect -100 -94739 -84 -94705
rect 84 -94739 100 -94705
rect -100 -94755 100 -94739
rect -100 -94813 100 -94797
rect -100 -94847 -84 -94813
rect 84 -94847 100 -94813
rect -100 -94894 100 -94847
rect -100 -96141 100 -96094
rect -100 -96175 -84 -96141
rect 84 -96175 100 -96141
rect -100 -96191 100 -96175
rect -100 -96249 100 -96233
rect -100 -96283 -84 -96249
rect 84 -96283 100 -96249
rect -100 -96330 100 -96283
rect -100 -97577 100 -97530
rect -100 -97611 -84 -97577
rect 84 -97611 100 -97577
rect -100 -97627 100 -97611
rect -100 -97685 100 -97669
rect -100 -97719 -84 -97685
rect 84 -97719 100 -97685
rect -100 -97766 100 -97719
rect -100 -99013 100 -98966
rect -100 -99047 -84 -99013
rect 84 -99047 100 -99013
rect -100 -99063 100 -99047
rect -100 -99121 100 -99105
rect -100 -99155 -84 -99121
rect 84 -99155 100 -99121
rect -100 -99202 100 -99155
rect -100 -100449 100 -100402
rect -100 -100483 -84 -100449
rect 84 -100483 100 -100449
rect -100 -100499 100 -100483
rect -100 -100557 100 -100541
rect -100 -100591 -84 -100557
rect 84 -100591 100 -100557
rect -100 -100638 100 -100591
rect -100 -101885 100 -101838
rect -100 -101919 -84 -101885
rect 84 -101919 100 -101885
rect -100 -101935 100 -101919
rect -100 -101993 100 -101977
rect -100 -102027 -84 -101993
rect 84 -102027 100 -101993
rect -100 -102074 100 -102027
rect -100 -103321 100 -103274
rect -100 -103355 -84 -103321
rect 84 -103355 100 -103321
rect -100 -103371 100 -103355
rect -100 -103429 100 -103413
rect -100 -103463 -84 -103429
rect 84 -103463 100 -103429
rect -100 -103510 100 -103463
rect -100 -104757 100 -104710
rect -100 -104791 -84 -104757
rect 84 -104791 100 -104757
rect -100 -104807 100 -104791
rect -100 -104865 100 -104849
rect -100 -104899 -84 -104865
rect 84 -104899 100 -104865
rect -100 -104946 100 -104899
rect -100 -106193 100 -106146
rect -100 -106227 -84 -106193
rect 84 -106227 100 -106193
rect -100 -106243 100 -106227
rect -100 -106301 100 -106285
rect -100 -106335 -84 -106301
rect 84 -106335 100 -106301
rect -100 -106382 100 -106335
rect -100 -107629 100 -107582
rect -100 -107663 -84 -107629
rect 84 -107663 100 -107629
rect -100 -107679 100 -107663
rect -100 -107737 100 -107721
rect -100 -107771 -84 -107737
rect 84 -107771 100 -107737
rect -100 -107818 100 -107771
rect -100 -109065 100 -109018
rect -100 -109099 -84 -109065
rect 84 -109099 100 -109065
rect -100 -109115 100 -109099
rect -100 -109173 100 -109157
rect -100 -109207 -84 -109173
rect 84 -109207 100 -109173
rect -100 -109254 100 -109207
rect -100 -110501 100 -110454
rect -100 -110535 -84 -110501
rect 84 -110535 100 -110501
rect -100 -110551 100 -110535
rect -100 -110609 100 -110593
rect -100 -110643 -84 -110609
rect 84 -110643 100 -110609
rect -100 -110690 100 -110643
rect -100 -111937 100 -111890
rect -100 -111971 -84 -111937
rect 84 -111971 100 -111937
rect -100 -111987 100 -111971
rect -100 -112045 100 -112029
rect -100 -112079 -84 -112045
rect 84 -112079 100 -112045
rect -100 -112126 100 -112079
rect -100 -113373 100 -113326
rect -100 -113407 -84 -113373
rect 84 -113407 100 -113373
rect -100 -113423 100 -113407
rect -100 -113481 100 -113465
rect -100 -113515 -84 -113481
rect 84 -113515 100 -113481
rect -100 -113562 100 -113515
rect -100 -114809 100 -114762
rect -100 -114843 -84 -114809
rect 84 -114843 100 -114809
rect -100 -114859 100 -114843
rect -100 -114917 100 -114901
rect -100 -114951 -84 -114917
rect 84 -114951 100 -114917
rect -100 -114998 100 -114951
rect -100 -116245 100 -116198
rect -100 -116279 -84 -116245
rect 84 -116279 100 -116245
rect -100 -116295 100 -116279
rect -100 -116353 100 -116337
rect -100 -116387 -84 -116353
rect 84 -116387 100 -116353
rect -100 -116434 100 -116387
rect -100 -117681 100 -117634
rect -100 -117715 -84 -117681
rect 84 -117715 100 -117681
rect -100 -117731 100 -117715
rect -100 -117789 100 -117773
rect -100 -117823 -84 -117789
rect 84 -117823 100 -117789
rect -100 -117870 100 -117823
rect -100 -119117 100 -119070
rect -100 -119151 -84 -119117
rect 84 -119151 100 -119117
rect -100 -119167 100 -119151
rect -100 -119225 100 -119209
rect -100 -119259 -84 -119225
rect 84 -119259 100 -119225
rect -100 -119306 100 -119259
rect -100 -120553 100 -120506
rect -100 -120587 -84 -120553
rect 84 -120587 100 -120553
rect -100 -120603 100 -120587
rect -100 -120661 100 -120645
rect -100 -120695 -84 -120661
rect 84 -120695 100 -120661
rect -100 -120742 100 -120695
rect -100 -121989 100 -121942
rect -100 -122023 -84 -121989
rect 84 -122023 100 -121989
rect -100 -122039 100 -122023
rect -100 -122097 100 -122081
rect -100 -122131 -84 -122097
rect 84 -122131 100 -122097
rect -100 -122178 100 -122131
rect -100 -123425 100 -123378
rect -100 -123459 -84 -123425
rect 84 -123459 100 -123425
rect -100 -123475 100 -123459
rect -100 -123533 100 -123517
rect -100 -123567 -84 -123533
rect 84 -123567 100 -123533
rect -100 -123614 100 -123567
rect -100 -124861 100 -124814
rect -100 -124895 -84 -124861
rect 84 -124895 100 -124861
rect -100 -124911 100 -124895
rect -100 -124969 100 -124953
rect -100 -125003 -84 -124969
rect 84 -125003 100 -124969
rect -100 -125050 100 -125003
rect -100 -126297 100 -126250
rect -100 -126331 -84 -126297
rect 84 -126331 100 -126297
rect -100 -126347 100 -126331
rect -100 -126405 100 -126389
rect -100 -126439 -84 -126405
rect 84 -126439 100 -126405
rect -100 -126486 100 -126439
rect -100 -127733 100 -127686
rect -100 -127767 -84 -127733
rect 84 -127767 100 -127733
rect -100 -127783 100 -127767
rect -100 -127841 100 -127825
rect -100 -127875 -84 -127841
rect 84 -127875 100 -127841
rect -100 -127922 100 -127875
rect -100 -129169 100 -129122
rect -100 -129203 -84 -129169
rect 84 -129203 100 -129169
rect -100 -129219 100 -129203
rect -100 -129277 100 -129261
rect -100 -129311 -84 -129277
rect 84 -129311 100 -129277
rect -100 -129358 100 -129311
rect -100 -130605 100 -130558
rect -100 -130639 -84 -130605
rect 84 -130639 100 -130605
rect -100 -130655 100 -130639
rect -100 -130713 100 -130697
rect -100 -130747 -84 -130713
rect 84 -130747 100 -130713
rect -100 -130794 100 -130747
rect -100 -132041 100 -131994
rect -100 -132075 -84 -132041
rect 84 -132075 100 -132041
rect -100 -132091 100 -132075
rect -100 -132149 100 -132133
rect -100 -132183 -84 -132149
rect 84 -132183 100 -132149
rect -100 -132230 100 -132183
rect -100 -133477 100 -133430
rect -100 -133511 -84 -133477
rect 84 -133511 100 -133477
rect -100 -133527 100 -133511
rect -100 -133585 100 -133569
rect -100 -133619 -84 -133585
rect 84 -133619 100 -133585
rect -100 -133666 100 -133619
rect -100 -134913 100 -134866
rect -100 -134947 -84 -134913
rect 84 -134947 100 -134913
rect -100 -134963 100 -134947
rect -100 -135021 100 -135005
rect -100 -135055 -84 -135021
rect 84 -135055 100 -135021
rect -100 -135102 100 -135055
rect -100 -136349 100 -136302
rect -100 -136383 -84 -136349
rect 84 -136383 100 -136349
rect -100 -136399 100 -136383
rect -100 -136457 100 -136441
rect -100 -136491 -84 -136457
rect 84 -136491 100 -136457
rect -100 -136538 100 -136491
rect -100 -137785 100 -137738
rect -100 -137819 -84 -137785
rect 84 -137819 100 -137785
rect -100 -137835 100 -137819
rect -100 -137893 100 -137877
rect -100 -137927 -84 -137893
rect 84 -137927 100 -137893
rect -100 -137974 100 -137927
rect -100 -139221 100 -139174
rect -100 -139255 -84 -139221
rect 84 -139255 100 -139221
rect -100 -139271 100 -139255
rect -100 -139329 100 -139313
rect -100 -139363 -84 -139329
rect 84 -139363 100 -139329
rect -100 -139410 100 -139363
rect -100 -140657 100 -140610
rect -100 -140691 -84 -140657
rect 84 -140691 100 -140657
rect -100 -140707 100 -140691
rect -100 -140765 100 -140749
rect -100 -140799 -84 -140765
rect 84 -140799 100 -140765
rect -100 -140846 100 -140799
rect -100 -142093 100 -142046
rect -100 -142127 -84 -142093
rect 84 -142127 100 -142093
rect -100 -142143 100 -142127
rect -100 -142201 100 -142185
rect -100 -142235 -84 -142201
rect 84 -142235 100 -142201
rect -100 -142282 100 -142235
rect -100 -143529 100 -143482
rect -100 -143563 -84 -143529
rect 84 -143563 100 -143529
rect -100 -143579 100 -143563
rect -100 -143637 100 -143621
rect -100 -143671 -84 -143637
rect 84 -143671 100 -143637
rect -100 -143718 100 -143671
rect -100 -144965 100 -144918
rect -100 -144999 -84 -144965
rect 84 -144999 100 -144965
rect -100 -145015 100 -144999
rect -100 -145073 100 -145057
rect -100 -145107 -84 -145073
rect 84 -145107 100 -145073
rect -100 -145154 100 -145107
rect -100 -146401 100 -146354
rect -100 -146435 -84 -146401
rect 84 -146435 100 -146401
rect -100 -146451 100 -146435
rect -100 -146509 100 -146493
rect -100 -146543 -84 -146509
rect 84 -146543 100 -146509
rect -100 -146590 100 -146543
rect -100 -147837 100 -147790
rect -100 -147871 -84 -147837
rect 84 -147871 100 -147837
rect -100 -147887 100 -147871
rect -100 -147945 100 -147929
rect -100 -147979 -84 -147945
rect 84 -147979 100 -147945
rect -100 -148026 100 -147979
rect -100 -149273 100 -149226
rect -100 -149307 -84 -149273
rect 84 -149307 100 -149273
rect -100 -149323 100 -149307
rect -100 -149381 100 -149365
rect -100 -149415 -84 -149381
rect 84 -149415 100 -149381
rect -100 -149462 100 -149415
rect -100 -150709 100 -150662
rect -100 -150743 -84 -150709
rect 84 -150743 100 -150709
rect -100 -150759 100 -150743
rect -100 -150817 100 -150801
rect -100 -150851 -84 -150817
rect 84 -150851 100 -150817
rect -100 -150898 100 -150851
rect -100 -152145 100 -152098
rect -100 -152179 -84 -152145
rect 84 -152179 100 -152145
rect -100 -152195 100 -152179
rect -100 -152253 100 -152237
rect -100 -152287 -84 -152253
rect 84 -152287 100 -152253
rect -100 -152334 100 -152287
rect -100 -153581 100 -153534
rect -100 -153615 -84 -153581
rect 84 -153615 100 -153581
rect -100 -153631 100 -153615
rect -100 -153689 100 -153673
rect -100 -153723 -84 -153689
rect 84 -153723 100 -153689
rect -100 -153770 100 -153723
rect -100 -155017 100 -154970
rect -100 -155051 -84 -155017
rect 84 -155051 100 -155017
rect -100 -155067 100 -155051
rect -100 -155125 100 -155109
rect -100 -155159 -84 -155125
rect 84 -155159 100 -155125
rect -100 -155206 100 -155159
rect -100 -156453 100 -156406
rect -100 -156487 -84 -156453
rect 84 -156487 100 -156453
rect -100 -156503 100 -156487
rect -100 -156561 100 -156545
rect -100 -156595 -84 -156561
rect 84 -156595 100 -156561
rect -100 -156642 100 -156595
rect -100 -157889 100 -157842
rect -100 -157923 -84 -157889
rect 84 -157923 100 -157889
rect -100 -157939 100 -157923
rect -100 -157997 100 -157981
rect -100 -158031 -84 -157997
rect 84 -158031 100 -157997
rect -100 -158078 100 -158031
rect -100 -159325 100 -159278
rect -100 -159359 -84 -159325
rect 84 -159359 100 -159325
rect -100 -159375 100 -159359
rect -100 -159433 100 -159417
rect -100 -159467 -84 -159433
rect 84 -159467 100 -159433
rect -100 -159514 100 -159467
rect -100 -160761 100 -160714
rect -100 -160795 -84 -160761
rect 84 -160795 100 -160761
rect -100 -160811 100 -160795
rect -100 -160869 100 -160853
rect -100 -160903 -84 -160869
rect 84 -160903 100 -160869
rect -100 -160950 100 -160903
rect -100 -162197 100 -162150
rect -100 -162231 -84 -162197
rect 84 -162231 100 -162197
rect -100 -162247 100 -162231
rect -100 -162305 100 -162289
rect -100 -162339 -84 -162305
rect 84 -162339 100 -162305
rect -100 -162386 100 -162339
rect -100 -163633 100 -163586
rect -100 -163667 -84 -163633
rect 84 -163667 100 -163633
rect -100 -163683 100 -163667
rect -100 -163741 100 -163725
rect -100 -163775 -84 -163741
rect 84 -163775 100 -163741
rect -100 -163822 100 -163775
rect -100 -165069 100 -165022
rect -100 -165103 -84 -165069
rect 84 -165103 100 -165069
rect -100 -165119 100 -165103
rect -100 -165177 100 -165161
rect -100 -165211 -84 -165177
rect 84 -165211 100 -165177
rect -100 -165258 100 -165211
rect -100 -166505 100 -166458
rect -100 -166539 -84 -166505
rect 84 -166539 100 -166505
rect -100 -166555 100 -166539
rect -100 -166613 100 -166597
rect -100 -166647 -84 -166613
rect 84 -166647 100 -166613
rect -100 -166694 100 -166647
rect -100 -167941 100 -167894
rect -100 -167975 -84 -167941
rect 84 -167975 100 -167941
rect -100 -167991 100 -167975
rect -100 -168049 100 -168033
rect -100 -168083 -84 -168049
rect 84 -168083 100 -168049
rect -100 -168130 100 -168083
rect -100 -169377 100 -169330
rect -100 -169411 -84 -169377
rect 84 -169411 100 -169377
rect -100 -169427 100 -169411
rect -100 -169485 100 -169469
rect -100 -169519 -84 -169485
rect 84 -169519 100 -169485
rect -100 -169566 100 -169519
rect -100 -170813 100 -170766
rect -100 -170847 -84 -170813
rect 84 -170847 100 -170813
rect -100 -170863 100 -170847
rect -100 -170921 100 -170905
rect -100 -170955 -84 -170921
rect 84 -170955 100 -170921
rect -100 -171002 100 -170955
rect -100 -172249 100 -172202
rect -100 -172283 -84 -172249
rect 84 -172283 100 -172249
rect -100 -172299 100 -172283
rect -100 -172357 100 -172341
rect -100 -172391 -84 -172357
rect 84 -172391 100 -172357
rect -100 -172438 100 -172391
rect -100 -173685 100 -173638
rect -100 -173719 -84 -173685
rect 84 -173719 100 -173685
rect -100 -173735 100 -173719
rect -100 -173793 100 -173777
rect -100 -173827 -84 -173793
rect 84 -173827 100 -173793
rect -100 -173874 100 -173827
rect -100 -175121 100 -175074
rect -100 -175155 -84 -175121
rect 84 -175155 100 -175121
rect -100 -175171 100 -175155
rect -100 -175229 100 -175213
rect -100 -175263 -84 -175229
rect 84 -175263 100 -175229
rect -100 -175310 100 -175263
rect -100 -176557 100 -176510
rect -100 -176591 -84 -176557
rect 84 -176591 100 -176557
rect -100 -176607 100 -176591
rect -100 -176665 100 -176649
rect -100 -176699 -84 -176665
rect 84 -176699 100 -176665
rect -100 -176746 100 -176699
rect -100 -177993 100 -177946
rect -100 -178027 -84 -177993
rect 84 -178027 100 -177993
rect -100 -178043 100 -178027
rect -100 -178101 100 -178085
rect -100 -178135 -84 -178101
rect 84 -178135 100 -178101
rect -100 -178182 100 -178135
rect -100 -179429 100 -179382
rect -100 -179463 -84 -179429
rect 84 -179463 100 -179429
rect -100 -179479 100 -179463
rect -100 -179537 100 -179521
rect -100 -179571 -84 -179537
rect 84 -179571 100 -179537
rect -100 -179618 100 -179571
rect -100 -180865 100 -180818
rect -100 -180899 -84 -180865
rect 84 -180899 100 -180865
rect -100 -180915 100 -180899
rect -100 -180973 100 -180957
rect -100 -181007 -84 -180973
rect 84 -181007 100 -180973
rect -100 -181054 100 -181007
rect -100 -182301 100 -182254
rect -100 -182335 -84 -182301
rect 84 -182335 100 -182301
rect -100 -182351 100 -182335
rect -100 -182409 100 -182393
rect -100 -182443 -84 -182409
rect 84 -182443 100 -182409
rect -100 -182490 100 -182443
rect -100 -183737 100 -183690
rect -100 -183771 -84 -183737
rect 84 -183771 100 -183737
rect -100 -183787 100 -183771
<< polycont >>
rect -84 183737 84 183771
rect -84 182409 84 182443
rect -84 182301 84 182335
rect -84 180973 84 181007
rect -84 180865 84 180899
rect -84 179537 84 179571
rect -84 179429 84 179463
rect -84 178101 84 178135
rect -84 177993 84 178027
rect -84 176665 84 176699
rect -84 176557 84 176591
rect -84 175229 84 175263
rect -84 175121 84 175155
rect -84 173793 84 173827
rect -84 173685 84 173719
rect -84 172357 84 172391
rect -84 172249 84 172283
rect -84 170921 84 170955
rect -84 170813 84 170847
rect -84 169485 84 169519
rect -84 169377 84 169411
rect -84 168049 84 168083
rect -84 167941 84 167975
rect -84 166613 84 166647
rect -84 166505 84 166539
rect -84 165177 84 165211
rect -84 165069 84 165103
rect -84 163741 84 163775
rect -84 163633 84 163667
rect -84 162305 84 162339
rect -84 162197 84 162231
rect -84 160869 84 160903
rect -84 160761 84 160795
rect -84 159433 84 159467
rect -84 159325 84 159359
rect -84 157997 84 158031
rect -84 157889 84 157923
rect -84 156561 84 156595
rect -84 156453 84 156487
rect -84 155125 84 155159
rect -84 155017 84 155051
rect -84 153689 84 153723
rect -84 153581 84 153615
rect -84 152253 84 152287
rect -84 152145 84 152179
rect -84 150817 84 150851
rect -84 150709 84 150743
rect -84 149381 84 149415
rect -84 149273 84 149307
rect -84 147945 84 147979
rect -84 147837 84 147871
rect -84 146509 84 146543
rect -84 146401 84 146435
rect -84 145073 84 145107
rect -84 144965 84 144999
rect -84 143637 84 143671
rect -84 143529 84 143563
rect -84 142201 84 142235
rect -84 142093 84 142127
rect -84 140765 84 140799
rect -84 140657 84 140691
rect -84 139329 84 139363
rect -84 139221 84 139255
rect -84 137893 84 137927
rect -84 137785 84 137819
rect -84 136457 84 136491
rect -84 136349 84 136383
rect -84 135021 84 135055
rect -84 134913 84 134947
rect -84 133585 84 133619
rect -84 133477 84 133511
rect -84 132149 84 132183
rect -84 132041 84 132075
rect -84 130713 84 130747
rect -84 130605 84 130639
rect -84 129277 84 129311
rect -84 129169 84 129203
rect -84 127841 84 127875
rect -84 127733 84 127767
rect -84 126405 84 126439
rect -84 126297 84 126331
rect -84 124969 84 125003
rect -84 124861 84 124895
rect -84 123533 84 123567
rect -84 123425 84 123459
rect -84 122097 84 122131
rect -84 121989 84 122023
rect -84 120661 84 120695
rect -84 120553 84 120587
rect -84 119225 84 119259
rect -84 119117 84 119151
rect -84 117789 84 117823
rect -84 117681 84 117715
rect -84 116353 84 116387
rect -84 116245 84 116279
rect -84 114917 84 114951
rect -84 114809 84 114843
rect -84 113481 84 113515
rect -84 113373 84 113407
rect -84 112045 84 112079
rect -84 111937 84 111971
rect -84 110609 84 110643
rect -84 110501 84 110535
rect -84 109173 84 109207
rect -84 109065 84 109099
rect -84 107737 84 107771
rect -84 107629 84 107663
rect -84 106301 84 106335
rect -84 106193 84 106227
rect -84 104865 84 104899
rect -84 104757 84 104791
rect -84 103429 84 103463
rect -84 103321 84 103355
rect -84 101993 84 102027
rect -84 101885 84 101919
rect -84 100557 84 100591
rect -84 100449 84 100483
rect -84 99121 84 99155
rect -84 99013 84 99047
rect -84 97685 84 97719
rect -84 97577 84 97611
rect -84 96249 84 96283
rect -84 96141 84 96175
rect -84 94813 84 94847
rect -84 94705 84 94739
rect -84 93377 84 93411
rect -84 93269 84 93303
rect -84 91941 84 91975
rect -84 91833 84 91867
rect -84 90505 84 90539
rect -84 90397 84 90431
rect -84 89069 84 89103
rect -84 88961 84 88995
rect -84 87633 84 87667
rect -84 87525 84 87559
rect -84 86197 84 86231
rect -84 86089 84 86123
rect -84 84761 84 84795
rect -84 84653 84 84687
rect -84 83325 84 83359
rect -84 83217 84 83251
rect -84 81889 84 81923
rect -84 81781 84 81815
rect -84 80453 84 80487
rect -84 80345 84 80379
rect -84 79017 84 79051
rect -84 78909 84 78943
rect -84 77581 84 77615
rect -84 77473 84 77507
rect -84 76145 84 76179
rect -84 76037 84 76071
rect -84 74709 84 74743
rect -84 74601 84 74635
rect -84 73273 84 73307
rect -84 73165 84 73199
rect -84 71837 84 71871
rect -84 71729 84 71763
rect -84 70401 84 70435
rect -84 70293 84 70327
rect -84 68965 84 68999
rect -84 68857 84 68891
rect -84 67529 84 67563
rect -84 67421 84 67455
rect -84 66093 84 66127
rect -84 65985 84 66019
rect -84 64657 84 64691
rect -84 64549 84 64583
rect -84 63221 84 63255
rect -84 63113 84 63147
rect -84 61785 84 61819
rect -84 61677 84 61711
rect -84 60349 84 60383
rect -84 60241 84 60275
rect -84 58913 84 58947
rect -84 58805 84 58839
rect -84 57477 84 57511
rect -84 57369 84 57403
rect -84 56041 84 56075
rect -84 55933 84 55967
rect -84 54605 84 54639
rect -84 54497 84 54531
rect -84 53169 84 53203
rect -84 53061 84 53095
rect -84 51733 84 51767
rect -84 51625 84 51659
rect -84 50297 84 50331
rect -84 50189 84 50223
rect -84 48861 84 48895
rect -84 48753 84 48787
rect -84 47425 84 47459
rect -84 47317 84 47351
rect -84 45989 84 46023
rect -84 45881 84 45915
rect -84 44553 84 44587
rect -84 44445 84 44479
rect -84 43117 84 43151
rect -84 43009 84 43043
rect -84 41681 84 41715
rect -84 41573 84 41607
rect -84 40245 84 40279
rect -84 40137 84 40171
rect -84 38809 84 38843
rect -84 38701 84 38735
rect -84 37373 84 37407
rect -84 37265 84 37299
rect -84 35937 84 35971
rect -84 35829 84 35863
rect -84 34501 84 34535
rect -84 34393 84 34427
rect -84 33065 84 33099
rect -84 32957 84 32991
rect -84 31629 84 31663
rect -84 31521 84 31555
rect -84 30193 84 30227
rect -84 30085 84 30119
rect -84 28757 84 28791
rect -84 28649 84 28683
rect -84 27321 84 27355
rect -84 27213 84 27247
rect -84 25885 84 25919
rect -84 25777 84 25811
rect -84 24449 84 24483
rect -84 24341 84 24375
rect -84 23013 84 23047
rect -84 22905 84 22939
rect -84 21577 84 21611
rect -84 21469 84 21503
rect -84 20141 84 20175
rect -84 20033 84 20067
rect -84 18705 84 18739
rect -84 18597 84 18631
rect -84 17269 84 17303
rect -84 17161 84 17195
rect -84 15833 84 15867
rect -84 15725 84 15759
rect -84 14397 84 14431
rect -84 14289 84 14323
rect -84 12961 84 12995
rect -84 12853 84 12887
rect -84 11525 84 11559
rect -84 11417 84 11451
rect -84 10089 84 10123
rect -84 9981 84 10015
rect -84 8653 84 8687
rect -84 8545 84 8579
rect -84 7217 84 7251
rect -84 7109 84 7143
rect -84 5781 84 5815
rect -84 5673 84 5707
rect -84 4345 84 4379
rect -84 4237 84 4271
rect -84 2909 84 2943
rect -84 2801 84 2835
rect -84 1473 84 1507
rect -84 1365 84 1399
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1399 84 -1365
rect -84 -1507 84 -1473
rect -84 -2835 84 -2801
rect -84 -2943 84 -2909
rect -84 -4271 84 -4237
rect -84 -4379 84 -4345
rect -84 -5707 84 -5673
rect -84 -5815 84 -5781
rect -84 -7143 84 -7109
rect -84 -7251 84 -7217
rect -84 -8579 84 -8545
rect -84 -8687 84 -8653
rect -84 -10015 84 -9981
rect -84 -10123 84 -10089
rect -84 -11451 84 -11417
rect -84 -11559 84 -11525
rect -84 -12887 84 -12853
rect -84 -12995 84 -12961
rect -84 -14323 84 -14289
rect -84 -14431 84 -14397
rect -84 -15759 84 -15725
rect -84 -15867 84 -15833
rect -84 -17195 84 -17161
rect -84 -17303 84 -17269
rect -84 -18631 84 -18597
rect -84 -18739 84 -18705
rect -84 -20067 84 -20033
rect -84 -20175 84 -20141
rect -84 -21503 84 -21469
rect -84 -21611 84 -21577
rect -84 -22939 84 -22905
rect -84 -23047 84 -23013
rect -84 -24375 84 -24341
rect -84 -24483 84 -24449
rect -84 -25811 84 -25777
rect -84 -25919 84 -25885
rect -84 -27247 84 -27213
rect -84 -27355 84 -27321
rect -84 -28683 84 -28649
rect -84 -28791 84 -28757
rect -84 -30119 84 -30085
rect -84 -30227 84 -30193
rect -84 -31555 84 -31521
rect -84 -31663 84 -31629
rect -84 -32991 84 -32957
rect -84 -33099 84 -33065
rect -84 -34427 84 -34393
rect -84 -34535 84 -34501
rect -84 -35863 84 -35829
rect -84 -35971 84 -35937
rect -84 -37299 84 -37265
rect -84 -37407 84 -37373
rect -84 -38735 84 -38701
rect -84 -38843 84 -38809
rect -84 -40171 84 -40137
rect -84 -40279 84 -40245
rect -84 -41607 84 -41573
rect -84 -41715 84 -41681
rect -84 -43043 84 -43009
rect -84 -43151 84 -43117
rect -84 -44479 84 -44445
rect -84 -44587 84 -44553
rect -84 -45915 84 -45881
rect -84 -46023 84 -45989
rect -84 -47351 84 -47317
rect -84 -47459 84 -47425
rect -84 -48787 84 -48753
rect -84 -48895 84 -48861
rect -84 -50223 84 -50189
rect -84 -50331 84 -50297
rect -84 -51659 84 -51625
rect -84 -51767 84 -51733
rect -84 -53095 84 -53061
rect -84 -53203 84 -53169
rect -84 -54531 84 -54497
rect -84 -54639 84 -54605
rect -84 -55967 84 -55933
rect -84 -56075 84 -56041
rect -84 -57403 84 -57369
rect -84 -57511 84 -57477
rect -84 -58839 84 -58805
rect -84 -58947 84 -58913
rect -84 -60275 84 -60241
rect -84 -60383 84 -60349
rect -84 -61711 84 -61677
rect -84 -61819 84 -61785
rect -84 -63147 84 -63113
rect -84 -63255 84 -63221
rect -84 -64583 84 -64549
rect -84 -64691 84 -64657
rect -84 -66019 84 -65985
rect -84 -66127 84 -66093
rect -84 -67455 84 -67421
rect -84 -67563 84 -67529
rect -84 -68891 84 -68857
rect -84 -68999 84 -68965
rect -84 -70327 84 -70293
rect -84 -70435 84 -70401
rect -84 -71763 84 -71729
rect -84 -71871 84 -71837
rect -84 -73199 84 -73165
rect -84 -73307 84 -73273
rect -84 -74635 84 -74601
rect -84 -74743 84 -74709
rect -84 -76071 84 -76037
rect -84 -76179 84 -76145
rect -84 -77507 84 -77473
rect -84 -77615 84 -77581
rect -84 -78943 84 -78909
rect -84 -79051 84 -79017
rect -84 -80379 84 -80345
rect -84 -80487 84 -80453
rect -84 -81815 84 -81781
rect -84 -81923 84 -81889
rect -84 -83251 84 -83217
rect -84 -83359 84 -83325
rect -84 -84687 84 -84653
rect -84 -84795 84 -84761
rect -84 -86123 84 -86089
rect -84 -86231 84 -86197
rect -84 -87559 84 -87525
rect -84 -87667 84 -87633
rect -84 -88995 84 -88961
rect -84 -89103 84 -89069
rect -84 -90431 84 -90397
rect -84 -90539 84 -90505
rect -84 -91867 84 -91833
rect -84 -91975 84 -91941
rect -84 -93303 84 -93269
rect -84 -93411 84 -93377
rect -84 -94739 84 -94705
rect -84 -94847 84 -94813
rect -84 -96175 84 -96141
rect -84 -96283 84 -96249
rect -84 -97611 84 -97577
rect -84 -97719 84 -97685
rect -84 -99047 84 -99013
rect -84 -99155 84 -99121
rect -84 -100483 84 -100449
rect -84 -100591 84 -100557
rect -84 -101919 84 -101885
rect -84 -102027 84 -101993
rect -84 -103355 84 -103321
rect -84 -103463 84 -103429
rect -84 -104791 84 -104757
rect -84 -104899 84 -104865
rect -84 -106227 84 -106193
rect -84 -106335 84 -106301
rect -84 -107663 84 -107629
rect -84 -107771 84 -107737
rect -84 -109099 84 -109065
rect -84 -109207 84 -109173
rect -84 -110535 84 -110501
rect -84 -110643 84 -110609
rect -84 -111971 84 -111937
rect -84 -112079 84 -112045
rect -84 -113407 84 -113373
rect -84 -113515 84 -113481
rect -84 -114843 84 -114809
rect -84 -114951 84 -114917
rect -84 -116279 84 -116245
rect -84 -116387 84 -116353
rect -84 -117715 84 -117681
rect -84 -117823 84 -117789
rect -84 -119151 84 -119117
rect -84 -119259 84 -119225
rect -84 -120587 84 -120553
rect -84 -120695 84 -120661
rect -84 -122023 84 -121989
rect -84 -122131 84 -122097
rect -84 -123459 84 -123425
rect -84 -123567 84 -123533
rect -84 -124895 84 -124861
rect -84 -125003 84 -124969
rect -84 -126331 84 -126297
rect -84 -126439 84 -126405
rect -84 -127767 84 -127733
rect -84 -127875 84 -127841
rect -84 -129203 84 -129169
rect -84 -129311 84 -129277
rect -84 -130639 84 -130605
rect -84 -130747 84 -130713
rect -84 -132075 84 -132041
rect -84 -132183 84 -132149
rect -84 -133511 84 -133477
rect -84 -133619 84 -133585
rect -84 -134947 84 -134913
rect -84 -135055 84 -135021
rect -84 -136383 84 -136349
rect -84 -136491 84 -136457
rect -84 -137819 84 -137785
rect -84 -137927 84 -137893
rect -84 -139255 84 -139221
rect -84 -139363 84 -139329
rect -84 -140691 84 -140657
rect -84 -140799 84 -140765
rect -84 -142127 84 -142093
rect -84 -142235 84 -142201
rect -84 -143563 84 -143529
rect -84 -143671 84 -143637
rect -84 -144999 84 -144965
rect -84 -145107 84 -145073
rect -84 -146435 84 -146401
rect -84 -146543 84 -146509
rect -84 -147871 84 -147837
rect -84 -147979 84 -147945
rect -84 -149307 84 -149273
rect -84 -149415 84 -149381
rect -84 -150743 84 -150709
rect -84 -150851 84 -150817
rect -84 -152179 84 -152145
rect -84 -152287 84 -152253
rect -84 -153615 84 -153581
rect -84 -153723 84 -153689
rect -84 -155051 84 -155017
rect -84 -155159 84 -155125
rect -84 -156487 84 -156453
rect -84 -156595 84 -156561
rect -84 -157923 84 -157889
rect -84 -158031 84 -157997
rect -84 -159359 84 -159325
rect -84 -159467 84 -159433
rect -84 -160795 84 -160761
rect -84 -160903 84 -160869
rect -84 -162231 84 -162197
rect -84 -162339 84 -162305
rect -84 -163667 84 -163633
rect -84 -163775 84 -163741
rect -84 -165103 84 -165069
rect -84 -165211 84 -165177
rect -84 -166539 84 -166505
rect -84 -166647 84 -166613
rect -84 -167975 84 -167941
rect -84 -168083 84 -168049
rect -84 -169411 84 -169377
rect -84 -169519 84 -169485
rect -84 -170847 84 -170813
rect -84 -170955 84 -170921
rect -84 -172283 84 -172249
rect -84 -172391 84 -172357
rect -84 -173719 84 -173685
rect -84 -173827 84 -173793
rect -84 -175155 84 -175121
rect -84 -175263 84 -175229
rect -84 -176591 84 -176557
rect -84 -176699 84 -176665
rect -84 -178027 84 -177993
rect -84 -178135 84 -178101
rect -84 -179463 84 -179429
rect -84 -179571 84 -179537
rect -84 -180899 84 -180865
rect -84 -181007 84 -180973
rect -84 -182335 84 -182301
rect -84 -182443 84 -182409
rect -84 -183771 84 -183737
<< locali >>
rect -280 183875 -184 183909
rect 184 183875 280 183909
rect -280 183813 -246 183875
rect 246 183813 280 183875
rect -100 183737 -84 183771
rect 84 183737 100 183771
rect -146 183678 -112 183694
rect -146 182486 -112 182502
rect 112 183678 146 183694
rect 112 182486 146 182502
rect -100 182409 -84 182443
rect 84 182409 100 182443
rect -100 182301 -84 182335
rect 84 182301 100 182335
rect -146 182242 -112 182258
rect -146 181050 -112 181066
rect 112 182242 146 182258
rect 112 181050 146 181066
rect -100 180973 -84 181007
rect 84 180973 100 181007
rect -100 180865 -84 180899
rect 84 180865 100 180899
rect -146 180806 -112 180822
rect -146 179614 -112 179630
rect 112 180806 146 180822
rect 112 179614 146 179630
rect -100 179537 -84 179571
rect 84 179537 100 179571
rect -100 179429 -84 179463
rect 84 179429 100 179463
rect -146 179370 -112 179386
rect -146 178178 -112 178194
rect 112 179370 146 179386
rect 112 178178 146 178194
rect -100 178101 -84 178135
rect 84 178101 100 178135
rect -100 177993 -84 178027
rect 84 177993 100 178027
rect -146 177934 -112 177950
rect -146 176742 -112 176758
rect 112 177934 146 177950
rect 112 176742 146 176758
rect -100 176665 -84 176699
rect 84 176665 100 176699
rect -100 176557 -84 176591
rect 84 176557 100 176591
rect -146 176498 -112 176514
rect -146 175306 -112 175322
rect 112 176498 146 176514
rect 112 175306 146 175322
rect -100 175229 -84 175263
rect 84 175229 100 175263
rect -100 175121 -84 175155
rect 84 175121 100 175155
rect -146 175062 -112 175078
rect -146 173870 -112 173886
rect 112 175062 146 175078
rect 112 173870 146 173886
rect -100 173793 -84 173827
rect 84 173793 100 173827
rect -100 173685 -84 173719
rect 84 173685 100 173719
rect -146 173626 -112 173642
rect -146 172434 -112 172450
rect 112 173626 146 173642
rect 112 172434 146 172450
rect -100 172357 -84 172391
rect 84 172357 100 172391
rect -100 172249 -84 172283
rect 84 172249 100 172283
rect -146 172190 -112 172206
rect -146 170998 -112 171014
rect 112 172190 146 172206
rect 112 170998 146 171014
rect -100 170921 -84 170955
rect 84 170921 100 170955
rect -100 170813 -84 170847
rect 84 170813 100 170847
rect -146 170754 -112 170770
rect -146 169562 -112 169578
rect 112 170754 146 170770
rect 112 169562 146 169578
rect -100 169485 -84 169519
rect 84 169485 100 169519
rect -100 169377 -84 169411
rect 84 169377 100 169411
rect -146 169318 -112 169334
rect -146 168126 -112 168142
rect 112 169318 146 169334
rect 112 168126 146 168142
rect -100 168049 -84 168083
rect 84 168049 100 168083
rect -100 167941 -84 167975
rect 84 167941 100 167975
rect -146 167882 -112 167898
rect -146 166690 -112 166706
rect 112 167882 146 167898
rect 112 166690 146 166706
rect -100 166613 -84 166647
rect 84 166613 100 166647
rect -100 166505 -84 166539
rect 84 166505 100 166539
rect -146 166446 -112 166462
rect -146 165254 -112 165270
rect 112 166446 146 166462
rect 112 165254 146 165270
rect -100 165177 -84 165211
rect 84 165177 100 165211
rect -100 165069 -84 165103
rect 84 165069 100 165103
rect -146 165010 -112 165026
rect -146 163818 -112 163834
rect 112 165010 146 165026
rect 112 163818 146 163834
rect -100 163741 -84 163775
rect 84 163741 100 163775
rect -100 163633 -84 163667
rect 84 163633 100 163667
rect -146 163574 -112 163590
rect -146 162382 -112 162398
rect 112 163574 146 163590
rect 112 162382 146 162398
rect -100 162305 -84 162339
rect 84 162305 100 162339
rect -100 162197 -84 162231
rect 84 162197 100 162231
rect -146 162138 -112 162154
rect -146 160946 -112 160962
rect 112 162138 146 162154
rect 112 160946 146 160962
rect -100 160869 -84 160903
rect 84 160869 100 160903
rect -100 160761 -84 160795
rect 84 160761 100 160795
rect -146 160702 -112 160718
rect -146 159510 -112 159526
rect 112 160702 146 160718
rect 112 159510 146 159526
rect -100 159433 -84 159467
rect 84 159433 100 159467
rect -100 159325 -84 159359
rect 84 159325 100 159359
rect -146 159266 -112 159282
rect -146 158074 -112 158090
rect 112 159266 146 159282
rect 112 158074 146 158090
rect -100 157997 -84 158031
rect 84 157997 100 158031
rect -100 157889 -84 157923
rect 84 157889 100 157923
rect -146 157830 -112 157846
rect -146 156638 -112 156654
rect 112 157830 146 157846
rect 112 156638 146 156654
rect -100 156561 -84 156595
rect 84 156561 100 156595
rect -100 156453 -84 156487
rect 84 156453 100 156487
rect -146 156394 -112 156410
rect -146 155202 -112 155218
rect 112 156394 146 156410
rect 112 155202 146 155218
rect -100 155125 -84 155159
rect 84 155125 100 155159
rect -100 155017 -84 155051
rect 84 155017 100 155051
rect -146 154958 -112 154974
rect -146 153766 -112 153782
rect 112 154958 146 154974
rect 112 153766 146 153782
rect -100 153689 -84 153723
rect 84 153689 100 153723
rect -100 153581 -84 153615
rect 84 153581 100 153615
rect -146 153522 -112 153538
rect -146 152330 -112 152346
rect 112 153522 146 153538
rect 112 152330 146 152346
rect -100 152253 -84 152287
rect 84 152253 100 152287
rect -100 152145 -84 152179
rect 84 152145 100 152179
rect -146 152086 -112 152102
rect -146 150894 -112 150910
rect 112 152086 146 152102
rect 112 150894 146 150910
rect -100 150817 -84 150851
rect 84 150817 100 150851
rect -100 150709 -84 150743
rect 84 150709 100 150743
rect -146 150650 -112 150666
rect -146 149458 -112 149474
rect 112 150650 146 150666
rect 112 149458 146 149474
rect -100 149381 -84 149415
rect 84 149381 100 149415
rect -100 149273 -84 149307
rect 84 149273 100 149307
rect -146 149214 -112 149230
rect -146 148022 -112 148038
rect 112 149214 146 149230
rect 112 148022 146 148038
rect -100 147945 -84 147979
rect 84 147945 100 147979
rect -100 147837 -84 147871
rect 84 147837 100 147871
rect -146 147778 -112 147794
rect -146 146586 -112 146602
rect 112 147778 146 147794
rect 112 146586 146 146602
rect -100 146509 -84 146543
rect 84 146509 100 146543
rect -100 146401 -84 146435
rect 84 146401 100 146435
rect -146 146342 -112 146358
rect -146 145150 -112 145166
rect 112 146342 146 146358
rect 112 145150 146 145166
rect -100 145073 -84 145107
rect 84 145073 100 145107
rect -100 144965 -84 144999
rect 84 144965 100 144999
rect -146 144906 -112 144922
rect -146 143714 -112 143730
rect 112 144906 146 144922
rect 112 143714 146 143730
rect -100 143637 -84 143671
rect 84 143637 100 143671
rect -100 143529 -84 143563
rect 84 143529 100 143563
rect -146 143470 -112 143486
rect -146 142278 -112 142294
rect 112 143470 146 143486
rect 112 142278 146 142294
rect -100 142201 -84 142235
rect 84 142201 100 142235
rect -100 142093 -84 142127
rect 84 142093 100 142127
rect -146 142034 -112 142050
rect -146 140842 -112 140858
rect 112 142034 146 142050
rect 112 140842 146 140858
rect -100 140765 -84 140799
rect 84 140765 100 140799
rect -100 140657 -84 140691
rect 84 140657 100 140691
rect -146 140598 -112 140614
rect -146 139406 -112 139422
rect 112 140598 146 140614
rect 112 139406 146 139422
rect -100 139329 -84 139363
rect 84 139329 100 139363
rect -100 139221 -84 139255
rect 84 139221 100 139255
rect -146 139162 -112 139178
rect -146 137970 -112 137986
rect 112 139162 146 139178
rect 112 137970 146 137986
rect -100 137893 -84 137927
rect 84 137893 100 137927
rect -100 137785 -84 137819
rect 84 137785 100 137819
rect -146 137726 -112 137742
rect -146 136534 -112 136550
rect 112 137726 146 137742
rect 112 136534 146 136550
rect -100 136457 -84 136491
rect 84 136457 100 136491
rect -100 136349 -84 136383
rect 84 136349 100 136383
rect -146 136290 -112 136306
rect -146 135098 -112 135114
rect 112 136290 146 136306
rect 112 135098 146 135114
rect -100 135021 -84 135055
rect 84 135021 100 135055
rect -100 134913 -84 134947
rect 84 134913 100 134947
rect -146 134854 -112 134870
rect -146 133662 -112 133678
rect 112 134854 146 134870
rect 112 133662 146 133678
rect -100 133585 -84 133619
rect 84 133585 100 133619
rect -100 133477 -84 133511
rect 84 133477 100 133511
rect -146 133418 -112 133434
rect -146 132226 -112 132242
rect 112 133418 146 133434
rect 112 132226 146 132242
rect -100 132149 -84 132183
rect 84 132149 100 132183
rect -100 132041 -84 132075
rect 84 132041 100 132075
rect -146 131982 -112 131998
rect -146 130790 -112 130806
rect 112 131982 146 131998
rect 112 130790 146 130806
rect -100 130713 -84 130747
rect 84 130713 100 130747
rect -100 130605 -84 130639
rect 84 130605 100 130639
rect -146 130546 -112 130562
rect -146 129354 -112 129370
rect 112 130546 146 130562
rect 112 129354 146 129370
rect -100 129277 -84 129311
rect 84 129277 100 129311
rect -100 129169 -84 129203
rect 84 129169 100 129203
rect -146 129110 -112 129126
rect -146 127918 -112 127934
rect 112 129110 146 129126
rect 112 127918 146 127934
rect -100 127841 -84 127875
rect 84 127841 100 127875
rect -100 127733 -84 127767
rect 84 127733 100 127767
rect -146 127674 -112 127690
rect -146 126482 -112 126498
rect 112 127674 146 127690
rect 112 126482 146 126498
rect -100 126405 -84 126439
rect 84 126405 100 126439
rect -100 126297 -84 126331
rect 84 126297 100 126331
rect -146 126238 -112 126254
rect -146 125046 -112 125062
rect 112 126238 146 126254
rect 112 125046 146 125062
rect -100 124969 -84 125003
rect 84 124969 100 125003
rect -100 124861 -84 124895
rect 84 124861 100 124895
rect -146 124802 -112 124818
rect -146 123610 -112 123626
rect 112 124802 146 124818
rect 112 123610 146 123626
rect -100 123533 -84 123567
rect 84 123533 100 123567
rect -100 123425 -84 123459
rect 84 123425 100 123459
rect -146 123366 -112 123382
rect -146 122174 -112 122190
rect 112 123366 146 123382
rect 112 122174 146 122190
rect -100 122097 -84 122131
rect 84 122097 100 122131
rect -100 121989 -84 122023
rect 84 121989 100 122023
rect -146 121930 -112 121946
rect -146 120738 -112 120754
rect 112 121930 146 121946
rect 112 120738 146 120754
rect -100 120661 -84 120695
rect 84 120661 100 120695
rect -100 120553 -84 120587
rect 84 120553 100 120587
rect -146 120494 -112 120510
rect -146 119302 -112 119318
rect 112 120494 146 120510
rect 112 119302 146 119318
rect -100 119225 -84 119259
rect 84 119225 100 119259
rect -100 119117 -84 119151
rect 84 119117 100 119151
rect -146 119058 -112 119074
rect -146 117866 -112 117882
rect 112 119058 146 119074
rect 112 117866 146 117882
rect -100 117789 -84 117823
rect 84 117789 100 117823
rect -100 117681 -84 117715
rect 84 117681 100 117715
rect -146 117622 -112 117638
rect -146 116430 -112 116446
rect 112 117622 146 117638
rect 112 116430 146 116446
rect -100 116353 -84 116387
rect 84 116353 100 116387
rect -100 116245 -84 116279
rect 84 116245 100 116279
rect -146 116186 -112 116202
rect -146 114994 -112 115010
rect 112 116186 146 116202
rect 112 114994 146 115010
rect -100 114917 -84 114951
rect 84 114917 100 114951
rect -100 114809 -84 114843
rect 84 114809 100 114843
rect -146 114750 -112 114766
rect -146 113558 -112 113574
rect 112 114750 146 114766
rect 112 113558 146 113574
rect -100 113481 -84 113515
rect 84 113481 100 113515
rect -100 113373 -84 113407
rect 84 113373 100 113407
rect -146 113314 -112 113330
rect -146 112122 -112 112138
rect 112 113314 146 113330
rect 112 112122 146 112138
rect -100 112045 -84 112079
rect 84 112045 100 112079
rect -100 111937 -84 111971
rect 84 111937 100 111971
rect -146 111878 -112 111894
rect -146 110686 -112 110702
rect 112 111878 146 111894
rect 112 110686 146 110702
rect -100 110609 -84 110643
rect 84 110609 100 110643
rect -100 110501 -84 110535
rect 84 110501 100 110535
rect -146 110442 -112 110458
rect -146 109250 -112 109266
rect 112 110442 146 110458
rect 112 109250 146 109266
rect -100 109173 -84 109207
rect 84 109173 100 109207
rect -100 109065 -84 109099
rect 84 109065 100 109099
rect -146 109006 -112 109022
rect -146 107814 -112 107830
rect 112 109006 146 109022
rect 112 107814 146 107830
rect -100 107737 -84 107771
rect 84 107737 100 107771
rect -100 107629 -84 107663
rect 84 107629 100 107663
rect -146 107570 -112 107586
rect -146 106378 -112 106394
rect 112 107570 146 107586
rect 112 106378 146 106394
rect -100 106301 -84 106335
rect 84 106301 100 106335
rect -100 106193 -84 106227
rect 84 106193 100 106227
rect -146 106134 -112 106150
rect -146 104942 -112 104958
rect 112 106134 146 106150
rect 112 104942 146 104958
rect -100 104865 -84 104899
rect 84 104865 100 104899
rect -100 104757 -84 104791
rect 84 104757 100 104791
rect -146 104698 -112 104714
rect -146 103506 -112 103522
rect 112 104698 146 104714
rect 112 103506 146 103522
rect -100 103429 -84 103463
rect 84 103429 100 103463
rect -100 103321 -84 103355
rect 84 103321 100 103355
rect -146 103262 -112 103278
rect -146 102070 -112 102086
rect 112 103262 146 103278
rect 112 102070 146 102086
rect -100 101993 -84 102027
rect 84 101993 100 102027
rect -100 101885 -84 101919
rect 84 101885 100 101919
rect -146 101826 -112 101842
rect -146 100634 -112 100650
rect 112 101826 146 101842
rect 112 100634 146 100650
rect -100 100557 -84 100591
rect 84 100557 100 100591
rect -100 100449 -84 100483
rect 84 100449 100 100483
rect -146 100390 -112 100406
rect -146 99198 -112 99214
rect 112 100390 146 100406
rect 112 99198 146 99214
rect -100 99121 -84 99155
rect 84 99121 100 99155
rect -100 99013 -84 99047
rect 84 99013 100 99047
rect -146 98954 -112 98970
rect -146 97762 -112 97778
rect 112 98954 146 98970
rect 112 97762 146 97778
rect -100 97685 -84 97719
rect 84 97685 100 97719
rect -100 97577 -84 97611
rect 84 97577 100 97611
rect -146 97518 -112 97534
rect -146 96326 -112 96342
rect 112 97518 146 97534
rect 112 96326 146 96342
rect -100 96249 -84 96283
rect 84 96249 100 96283
rect -100 96141 -84 96175
rect 84 96141 100 96175
rect -146 96082 -112 96098
rect -146 94890 -112 94906
rect 112 96082 146 96098
rect 112 94890 146 94906
rect -100 94813 -84 94847
rect 84 94813 100 94847
rect -100 94705 -84 94739
rect 84 94705 100 94739
rect -146 94646 -112 94662
rect -146 93454 -112 93470
rect 112 94646 146 94662
rect 112 93454 146 93470
rect -100 93377 -84 93411
rect 84 93377 100 93411
rect -100 93269 -84 93303
rect 84 93269 100 93303
rect -146 93210 -112 93226
rect -146 92018 -112 92034
rect 112 93210 146 93226
rect 112 92018 146 92034
rect -100 91941 -84 91975
rect 84 91941 100 91975
rect -100 91833 -84 91867
rect 84 91833 100 91867
rect -146 91774 -112 91790
rect -146 90582 -112 90598
rect 112 91774 146 91790
rect 112 90582 146 90598
rect -100 90505 -84 90539
rect 84 90505 100 90539
rect -100 90397 -84 90431
rect 84 90397 100 90431
rect -146 90338 -112 90354
rect -146 89146 -112 89162
rect 112 90338 146 90354
rect 112 89146 146 89162
rect -100 89069 -84 89103
rect 84 89069 100 89103
rect -100 88961 -84 88995
rect 84 88961 100 88995
rect -146 88902 -112 88918
rect -146 87710 -112 87726
rect 112 88902 146 88918
rect 112 87710 146 87726
rect -100 87633 -84 87667
rect 84 87633 100 87667
rect -100 87525 -84 87559
rect 84 87525 100 87559
rect -146 87466 -112 87482
rect -146 86274 -112 86290
rect 112 87466 146 87482
rect 112 86274 146 86290
rect -100 86197 -84 86231
rect 84 86197 100 86231
rect -100 86089 -84 86123
rect 84 86089 100 86123
rect -146 86030 -112 86046
rect -146 84838 -112 84854
rect 112 86030 146 86046
rect 112 84838 146 84854
rect -100 84761 -84 84795
rect 84 84761 100 84795
rect -100 84653 -84 84687
rect 84 84653 100 84687
rect -146 84594 -112 84610
rect -146 83402 -112 83418
rect 112 84594 146 84610
rect 112 83402 146 83418
rect -100 83325 -84 83359
rect 84 83325 100 83359
rect -100 83217 -84 83251
rect 84 83217 100 83251
rect -146 83158 -112 83174
rect -146 81966 -112 81982
rect 112 83158 146 83174
rect 112 81966 146 81982
rect -100 81889 -84 81923
rect 84 81889 100 81923
rect -100 81781 -84 81815
rect 84 81781 100 81815
rect -146 81722 -112 81738
rect -146 80530 -112 80546
rect 112 81722 146 81738
rect 112 80530 146 80546
rect -100 80453 -84 80487
rect 84 80453 100 80487
rect -100 80345 -84 80379
rect 84 80345 100 80379
rect -146 80286 -112 80302
rect -146 79094 -112 79110
rect 112 80286 146 80302
rect 112 79094 146 79110
rect -100 79017 -84 79051
rect 84 79017 100 79051
rect -100 78909 -84 78943
rect 84 78909 100 78943
rect -146 78850 -112 78866
rect -146 77658 -112 77674
rect 112 78850 146 78866
rect 112 77658 146 77674
rect -100 77581 -84 77615
rect 84 77581 100 77615
rect -100 77473 -84 77507
rect 84 77473 100 77507
rect -146 77414 -112 77430
rect -146 76222 -112 76238
rect 112 77414 146 77430
rect 112 76222 146 76238
rect -100 76145 -84 76179
rect 84 76145 100 76179
rect -100 76037 -84 76071
rect 84 76037 100 76071
rect -146 75978 -112 75994
rect -146 74786 -112 74802
rect 112 75978 146 75994
rect 112 74786 146 74802
rect -100 74709 -84 74743
rect 84 74709 100 74743
rect -100 74601 -84 74635
rect 84 74601 100 74635
rect -146 74542 -112 74558
rect -146 73350 -112 73366
rect 112 74542 146 74558
rect 112 73350 146 73366
rect -100 73273 -84 73307
rect 84 73273 100 73307
rect -100 73165 -84 73199
rect 84 73165 100 73199
rect -146 73106 -112 73122
rect -146 71914 -112 71930
rect 112 73106 146 73122
rect 112 71914 146 71930
rect -100 71837 -84 71871
rect 84 71837 100 71871
rect -100 71729 -84 71763
rect 84 71729 100 71763
rect -146 71670 -112 71686
rect -146 70478 -112 70494
rect 112 71670 146 71686
rect 112 70478 146 70494
rect -100 70401 -84 70435
rect 84 70401 100 70435
rect -100 70293 -84 70327
rect 84 70293 100 70327
rect -146 70234 -112 70250
rect -146 69042 -112 69058
rect 112 70234 146 70250
rect 112 69042 146 69058
rect -100 68965 -84 68999
rect 84 68965 100 68999
rect -100 68857 -84 68891
rect 84 68857 100 68891
rect -146 68798 -112 68814
rect -146 67606 -112 67622
rect 112 68798 146 68814
rect 112 67606 146 67622
rect -100 67529 -84 67563
rect 84 67529 100 67563
rect -100 67421 -84 67455
rect 84 67421 100 67455
rect -146 67362 -112 67378
rect -146 66170 -112 66186
rect 112 67362 146 67378
rect 112 66170 146 66186
rect -100 66093 -84 66127
rect 84 66093 100 66127
rect -100 65985 -84 66019
rect 84 65985 100 66019
rect -146 65926 -112 65942
rect -146 64734 -112 64750
rect 112 65926 146 65942
rect 112 64734 146 64750
rect -100 64657 -84 64691
rect 84 64657 100 64691
rect -100 64549 -84 64583
rect 84 64549 100 64583
rect -146 64490 -112 64506
rect -146 63298 -112 63314
rect 112 64490 146 64506
rect 112 63298 146 63314
rect -100 63221 -84 63255
rect 84 63221 100 63255
rect -100 63113 -84 63147
rect 84 63113 100 63147
rect -146 63054 -112 63070
rect -146 61862 -112 61878
rect 112 63054 146 63070
rect 112 61862 146 61878
rect -100 61785 -84 61819
rect 84 61785 100 61819
rect -100 61677 -84 61711
rect 84 61677 100 61711
rect -146 61618 -112 61634
rect -146 60426 -112 60442
rect 112 61618 146 61634
rect 112 60426 146 60442
rect -100 60349 -84 60383
rect 84 60349 100 60383
rect -100 60241 -84 60275
rect 84 60241 100 60275
rect -146 60182 -112 60198
rect -146 58990 -112 59006
rect 112 60182 146 60198
rect 112 58990 146 59006
rect -100 58913 -84 58947
rect 84 58913 100 58947
rect -100 58805 -84 58839
rect 84 58805 100 58839
rect -146 58746 -112 58762
rect -146 57554 -112 57570
rect 112 58746 146 58762
rect 112 57554 146 57570
rect -100 57477 -84 57511
rect 84 57477 100 57511
rect -100 57369 -84 57403
rect 84 57369 100 57403
rect -146 57310 -112 57326
rect -146 56118 -112 56134
rect 112 57310 146 57326
rect 112 56118 146 56134
rect -100 56041 -84 56075
rect 84 56041 100 56075
rect -100 55933 -84 55967
rect 84 55933 100 55967
rect -146 55874 -112 55890
rect -146 54682 -112 54698
rect 112 55874 146 55890
rect 112 54682 146 54698
rect -100 54605 -84 54639
rect 84 54605 100 54639
rect -100 54497 -84 54531
rect 84 54497 100 54531
rect -146 54438 -112 54454
rect -146 53246 -112 53262
rect 112 54438 146 54454
rect 112 53246 146 53262
rect -100 53169 -84 53203
rect 84 53169 100 53203
rect -100 53061 -84 53095
rect 84 53061 100 53095
rect -146 53002 -112 53018
rect -146 51810 -112 51826
rect 112 53002 146 53018
rect 112 51810 146 51826
rect -100 51733 -84 51767
rect 84 51733 100 51767
rect -100 51625 -84 51659
rect 84 51625 100 51659
rect -146 51566 -112 51582
rect -146 50374 -112 50390
rect 112 51566 146 51582
rect 112 50374 146 50390
rect -100 50297 -84 50331
rect 84 50297 100 50331
rect -100 50189 -84 50223
rect 84 50189 100 50223
rect -146 50130 -112 50146
rect -146 48938 -112 48954
rect 112 50130 146 50146
rect 112 48938 146 48954
rect -100 48861 -84 48895
rect 84 48861 100 48895
rect -100 48753 -84 48787
rect 84 48753 100 48787
rect -146 48694 -112 48710
rect -146 47502 -112 47518
rect 112 48694 146 48710
rect 112 47502 146 47518
rect -100 47425 -84 47459
rect 84 47425 100 47459
rect -100 47317 -84 47351
rect 84 47317 100 47351
rect -146 47258 -112 47274
rect -146 46066 -112 46082
rect 112 47258 146 47274
rect 112 46066 146 46082
rect -100 45989 -84 46023
rect 84 45989 100 46023
rect -100 45881 -84 45915
rect 84 45881 100 45915
rect -146 45822 -112 45838
rect -146 44630 -112 44646
rect 112 45822 146 45838
rect 112 44630 146 44646
rect -100 44553 -84 44587
rect 84 44553 100 44587
rect -100 44445 -84 44479
rect 84 44445 100 44479
rect -146 44386 -112 44402
rect -146 43194 -112 43210
rect 112 44386 146 44402
rect 112 43194 146 43210
rect -100 43117 -84 43151
rect 84 43117 100 43151
rect -100 43009 -84 43043
rect 84 43009 100 43043
rect -146 42950 -112 42966
rect -146 41758 -112 41774
rect 112 42950 146 42966
rect 112 41758 146 41774
rect -100 41681 -84 41715
rect 84 41681 100 41715
rect -100 41573 -84 41607
rect 84 41573 100 41607
rect -146 41514 -112 41530
rect -146 40322 -112 40338
rect 112 41514 146 41530
rect 112 40322 146 40338
rect -100 40245 -84 40279
rect 84 40245 100 40279
rect -100 40137 -84 40171
rect 84 40137 100 40171
rect -146 40078 -112 40094
rect -146 38886 -112 38902
rect 112 40078 146 40094
rect 112 38886 146 38902
rect -100 38809 -84 38843
rect 84 38809 100 38843
rect -100 38701 -84 38735
rect 84 38701 100 38735
rect -146 38642 -112 38658
rect -146 37450 -112 37466
rect 112 38642 146 38658
rect 112 37450 146 37466
rect -100 37373 -84 37407
rect 84 37373 100 37407
rect -100 37265 -84 37299
rect 84 37265 100 37299
rect -146 37206 -112 37222
rect -146 36014 -112 36030
rect 112 37206 146 37222
rect 112 36014 146 36030
rect -100 35937 -84 35971
rect 84 35937 100 35971
rect -100 35829 -84 35863
rect 84 35829 100 35863
rect -146 35770 -112 35786
rect -146 34578 -112 34594
rect 112 35770 146 35786
rect 112 34578 146 34594
rect -100 34501 -84 34535
rect 84 34501 100 34535
rect -100 34393 -84 34427
rect 84 34393 100 34427
rect -146 34334 -112 34350
rect -146 33142 -112 33158
rect 112 34334 146 34350
rect 112 33142 146 33158
rect -100 33065 -84 33099
rect 84 33065 100 33099
rect -100 32957 -84 32991
rect 84 32957 100 32991
rect -146 32898 -112 32914
rect -146 31706 -112 31722
rect 112 32898 146 32914
rect 112 31706 146 31722
rect -100 31629 -84 31663
rect 84 31629 100 31663
rect -100 31521 -84 31555
rect 84 31521 100 31555
rect -146 31462 -112 31478
rect -146 30270 -112 30286
rect 112 31462 146 31478
rect 112 30270 146 30286
rect -100 30193 -84 30227
rect 84 30193 100 30227
rect -100 30085 -84 30119
rect 84 30085 100 30119
rect -146 30026 -112 30042
rect -146 28834 -112 28850
rect 112 30026 146 30042
rect 112 28834 146 28850
rect -100 28757 -84 28791
rect 84 28757 100 28791
rect -100 28649 -84 28683
rect 84 28649 100 28683
rect -146 28590 -112 28606
rect -146 27398 -112 27414
rect 112 28590 146 28606
rect 112 27398 146 27414
rect -100 27321 -84 27355
rect 84 27321 100 27355
rect -100 27213 -84 27247
rect 84 27213 100 27247
rect -146 27154 -112 27170
rect -146 25962 -112 25978
rect 112 27154 146 27170
rect 112 25962 146 25978
rect -100 25885 -84 25919
rect 84 25885 100 25919
rect -100 25777 -84 25811
rect 84 25777 100 25811
rect -146 25718 -112 25734
rect -146 24526 -112 24542
rect 112 25718 146 25734
rect 112 24526 146 24542
rect -100 24449 -84 24483
rect 84 24449 100 24483
rect -100 24341 -84 24375
rect 84 24341 100 24375
rect -146 24282 -112 24298
rect -146 23090 -112 23106
rect 112 24282 146 24298
rect 112 23090 146 23106
rect -100 23013 -84 23047
rect 84 23013 100 23047
rect -100 22905 -84 22939
rect 84 22905 100 22939
rect -146 22846 -112 22862
rect -146 21654 -112 21670
rect 112 22846 146 22862
rect 112 21654 146 21670
rect -100 21577 -84 21611
rect 84 21577 100 21611
rect -100 21469 -84 21503
rect 84 21469 100 21503
rect -146 21410 -112 21426
rect -146 20218 -112 20234
rect 112 21410 146 21426
rect 112 20218 146 20234
rect -100 20141 -84 20175
rect 84 20141 100 20175
rect -100 20033 -84 20067
rect 84 20033 100 20067
rect -146 19974 -112 19990
rect -146 18782 -112 18798
rect 112 19974 146 19990
rect 112 18782 146 18798
rect -100 18705 -84 18739
rect 84 18705 100 18739
rect -100 18597 -84 18631
rect 84 18597 100 18631
rect -146 18538 -112 18554
rect -146 17346 -112 17362
rect 112 18538 146 18554
rect 112 17346 146 17362
rect -100 17269 -84 17303
rect 84 17269 100 17303
rect -100 17161 -84 17195
rect 84 17161 100 17195
rect -146 17102 -112 17118
rect -146 15910 -112 15926
rect 112 17102 146 17118
rect 112 15910 146 15926
rect -100 15833 -84 15867
rect 84 15833 100 15867
rect -100 15725 -84 15759
rect 84 15725 100 15759
rect -146 15666 -112 15682
rect -146 14474 -112 14490
rect 112 15666 146 15682
rect 112 14474 146 14490
rect -100 14397 -84 14431
rect 84 14397 100 14431
rect -100 14289 -84 14323
rect 84 14289 100 14323
rect -146 14230 -112 14246
rect -146 13038 -112 13054
rect 112 14230 146 14246
rect 112 13038 146 13054
rect -100 12961 -84 12995
rect 84 12961 100 12995
rect -100 12853 -84 12887
rect 84 12853 100 12887
rect -146 12794 -112 12810
rect -146 11602 -112 11618
rect 112 12794 146 12810
rect 112 11602 146 11618
rect -100 11525 -84 11559
rect 84 11525 100 11559
rect -100 11417 -84 11451
rect 84 11417 100 11451
rect -146 11358 -112 11374
rect -146 10166 -112 10182
rect 112 11358 146 11374
rect 112 10166 146 10182
rect -100 10089 -84 10123
rect 84 10089 100 10123
rect -100 9981 -84 10015
rect 84 9981 100 10015
rect -146 9922 -112 9938
rect -146 8730 -112 8746
rect 112 9922 146 9938
rect 112 8730 146 8746
rect -100 8653 -84 8687
rect 84 8653 100 8687
rect -100 8545 -84 8579
rect 84 8545 100 8579
rect -146 8486 -112 8502
rect -146 7294 -112 7310
rect 112 8486 146 8502
rect 112 7294 146 7310
rect -100 7217 -84 7251
rect 84 7217 100 7251
rect -100 7109 -84 7143
rect 84 7109 100 7143
rect -146 7050 -112 7066
rect -146 5858 -112 5874
rect 112 7050 146 7066
rect 112 5858 146 5874
rect -100 5781 -84 5815
rect 84 5781 100 5815
rect -100 5673 -84 5707
rect 84 5673 100 5707
rect -146 5614 -112 5630
rect -146 4422 -112 4438
rect 112 5614 146 5630
rect 112 4422 146 4438
rect -100 4345 -84 4379
rect 84 4345 100 4379
rect -100 4237 -84 4271
rect 84 4237 100 4271
rect -146 4178 -112 4194
rect -146 2986 -112 3002
rect 112 4178 146 4194
rect 112 2986 146 3002
rect -100 2909 -84 2943
rect 84 2909 100 2943
rect -100 2801 -84 2835
rect 84 2801 100 2835
rect -146 2742 -112 2758
rect -146 1550 -112 1566
rect 112 2742 146 2758
rect 112 1550 146 1566
rect -100 1473 -84 1507
rect 84 1473 100 1507
rect -100 1365 -84 1399
rect 84 1365 100 1399
rect -146 1306 -112 1322
rect -146 114 -112 130
rect 112 1306 146 1322
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -1322 -112 -1306
rect 112 -130 146 -114
rect 112 -1322 146 -1306
rect -100 -1399 -84 -1365
rect 84 -1399 100 -1365
rect -100 -1507 -84 -1473
rect 84 -1507 100 -1473
rect -146 -1566 -112 -1550
rect -146 -2758 -112 -2742
rect 112 -1566 146 -1550
rect 112 -2758 146 -2742
rect -100 -2835 -84 -2801
rect 84 -2835 100 -2801
rect -100 -2943 -84 -2909
rect 84 -2943 100 -2909
rect -146 -3002 -112 -2986
rect -146 -4194 -112 -4178
rect 112 -3002 146 -2986
rect 112 -4194 146 -4178
rect -100 -4271 -84 -4237
rect 84 -4271 100 -4237
rect -100 -4379 -84 -4345
rect 84 -4379 100 -4345
rect -146 -4438 -112 -4422
rect -146 -5630 -112 -5614
rect 112 -4438 146 -4422
rect 112 -5630 146 -5614
rect -100 -5707 -84 -5673
rect 84 -5707 100 -5673
rect -100 -5815 -84 -5781
rect 84 -5815 100 -5781
rect -146 -5874 -112 -5858
rect -146 -7066 -112 -7050
rect 112 -5874 146 -5858
rect 112 -7066 146 -7050
rect -100 -7143 -84 -7109
rect 84 -7143 100 -7109
rect -100 -7251 -84 -7217
rect 84 -7251 100 -7217
rect -146 -7310 -112 -7294
rect -146 -8502 -112 -8486
rect 112 -7310 146 -7294
rect 112 -8502 146 -8486
rect -100 -8579 -84 -8545
rect 84 -8579 100 -8545
rect -100 -8687 -84 -8653
rect 84 -8687 100 -8653
rect -146 -8746 -112 -8730
rect -146 -9938 -112 -9922
rect 112 -8746 146 -8730
rect 112 -9938 146 -9922
rect -100 -10015 -84 -9981
rect 84 -10015 100 -9981
rect -100 -10123 -84 -10089
rect 84 -10123 100 -10089
rect -146 -10182 -112 -10166
rect -146 -11374 -112 -11358
rect 112 -10182 146 -10166
rect 112 -11374 146 -11358
rect -100 -11451 -84 -11417
rect 84 -11451 100 -11417
rect -100 -11559 -84 -11525
rect 84 -11559 100 -11525
rect -146 -11618 -112 -11602
rect -146 -12810 -112 -12794
rect 112 -11618 146 -11602
rect 112 -12810 146 -12794
rect -100 -12887 -84 -12853
rect 84 -12887 100 -12853
rect -100 -12995 -84 -12961
rect 84 -12995 100 -12961
rect -146 -13054 -112 -13038
rect -146 -14246 -112 -14230
rect 112 -13054 146 -13038
rect 112 -14246 146 -14230
rect -100 -14323 -84 -14289
rect 84 -14323 100 -14289
rect -100 -14431 -84 -14397
rect 84 -14431 100 -14397
rect -146 -14490 -112 -14474
rect -146 -15682 -112 -15666
rect 112 -14490 146 -14474
rect 112 -15682 146 -15666
rect -100 -15759 -84 -15725
rect 84 -15759 100 -15725
rect -100 -15867 -84 -15833
rect 84 -15867 100 -15833
rect -146 -15926 -112 -15910
rect -146 -17118 -112 -17102
rect 112 -15926 146 -15910
rect 112 -17118 146 -17102
rect -100 -17195 -84 -17161
rect 84 -17195 100 -17161
rect -100 -17303 -84 -17269
rect 84 -17303 100 -17269
rect -146 -17362 -112 -17346
rect -146 -18554 -112 -18538
rect 112 -17362 146 -17346
rect 112 -18554 146 -18538
rect -100 -18631 -84 -18597
rect 84 -18631 100 -18597
rect -100 -18739 -84 -18705
rect 84 -18739 100 -18705
rect -146 -18798 -112 -18782
rect -146 -19990 -112 -19974
rect 112 -18798 146 -18782
rect 112 -19990 146 -19974
rect -100 -20067 -84 -20033
rect 84 -20067 100 -20033
rect -100 -20175 -84 -20141
rect 84 -20175 100 -20141
rect -146 -20234 -112 -20218
rect -146 -21426 -112 -21410
rect 112 -20234 146 -20218
rect 112 -21426 146 -21410
rect -100 -21503 -84 -21469
rect 84 -21503 100 -21469
rect -100 -21611 -84 -21577
rect 84 -21611 100 -21577
rect -146 -21670 -112 -21654
rect -146 -22862 -112 -22846
rect 112 -21670 146 -21654
rect 112 -22862 146 -22846
rect -100 -22939 -84 -22905
rect 84 -22939 100 -22905
rect -100 -23047 -84 -23013
rect 84 -23047 100 -23013
rect -146 -23106 -112 -23090
rect -146 -24298 -112 -24282
rect 112 -23106 146 -23090
rect 112 -24298 146 -24282
rect -100 -24375 -84 -24341
rect 84 -24375 100 -24341
rect -100 -24483 -84 -24449
rect 84 -24483 100 -24449
rect -146 -24542 -112 -24526
rect -146 -25734 -112 -25718
rect 112 -24542 146 -24526
rect 112 -25734 146 -25718
rect -100 -25811 -84 -25777
rect 84 -25811 100 -25777
rect -100 -25919 -84 -25885
rect 84 -25919 100 -25885
rect -146 -25978 -112 -25962
rect -146 -27170 -112 -27154
rect 112 -25978 146 -25962
rect 112 -27170 146 -27154
rect -100 -27247 -84 -27213
rect 84 -27247 100 -27213
rect -100 -27355 -84 -27321
rect 84 -27355 100 -27321
rect -146 -27414 -112 -27398
rect -146 -28606 -112 -28590
rect 112 -27414 146 -27398
rect 112 -28606 146 -28590
rect -100 -28683 -84 -28649
rect 84 -28683 100 -28649
rect -100 -28791 -84 -28757
rect 84 -28791 100 -28757
rect -146 -28850 -112 -28834
rect -146 -30042 -112 -30026
rect 112 -28850 146 -28834
rect 112 -30042 146 -30026
rect -100 -30119 -84 -30085
rect 84 -30119 100 -30085
rect -100 -30227 -84 -30193
rect 84 -30227 100 -30193
rect -146 -30286 -112 -30270
rect -146 -31478 -112 -31462
rect 112 -30286 146 -30270
rect 112 -31478 146 -31462
rect -100 -31555 -84 -31521
rect 84 -31555 100 -31521
rect -100 -31663 -84 -31629
rect 84 -31663 100 -31629
rect -146 -31722 -112 -31706
rect -146 -32914 -112 -32898
rect 112 -31722 146 -31706
rect 112 -32914 146 -32898
rect -100 -32991 -84 -32957
rect 84 -32991 100 -32957
rect -100 -33099 -84 -33065
rect 84 -33099 100 -33065
rect -146 -33158 -112 -33142
rect -146 -34350 -112 -34334
rect 112 -33158 146 -33142
rect 112 -34350 146 -34334
rect -100 -34427 -84 -34393
rect 84 -34427 100 -34393
rect -100 -34535 -84 -34501
rect 84 -34535 100 -34501
rect -146 -34594 -112 -34578
rect -146 -35786 -112 -35770
rect 112 -34594 146 -34578
rect 112 -35786 146 -35770
rect -100 -35863 -84 -35829
rect 84 -35863 100 -35829
rect -100 -35971 -84 -35937
rect 84 -35971 100 -35937
rect -146 -36030 -112 -36014
rect -146 -37222 -112 -37206
rect 112 -36030 146 -36014
rect 112 -37222 146 -37206
rect -100 -37299 -84 -37265
rect 84 -37299 100 -37265
rect -100 -37407 -84 -37373
rect 84 -37407 100 -37373
rect -146 -37466 -112 -37450
rect -146 -38658 -112 -38642
rect 112 -37466 146 -37450
rect 112 -38658 146 -38642
rect -100 -38735 -84 -38701
rect 84 -38735 100 -38701
rect -100 -38843 -84 -38809
rect 84 -38843 100 -38809
rect -146 -38902 -112 -38886
rect -146 -40094 -112 -40078
rect 112 -38902 146 -38886
rect 112 -40094 146 -40078
rect -100 -40171 -84 -40137
rect 84 -40171 100 -40137
rect -100 -40279 -84 -40245
rect 84 -40279 100 -40245
rect -146 -40338 -112 -40322
rect -146 -41530 -112 -41514
rect 112 -40338 146 -40322
rect 112 -41530 146 -41514
rect -100 -41607 -84 -41573
rect 84 -41607 100 -41573
rect -100 -41715 -84 -41681
rect 84 -41715 100 -41681
rect -146 -41774 -112 -41758
rect -146 -42966 -112 -42950
rect 112 -41774 146 -41758
rect 112 -42966 146 -42950
rect -100 -43043 -84 -43009
rect 84 -43043 100 -43009
rect -100 -43151 -84 -43117
rect 84 -43151 100 -43117
rect -146 -43210 -112 -43194
rect -146 -44402 -112 -44386
rect 112 -43210 146 -43194
rect 112 -44402 146 -44386
rect -100 -44479 -84 -44445
rect 84 -44479 100 -44445
rect -100 -44587 -84 -44553
rect 84 -44587 100 -44553
rect -146 -44646 -112 -44630
rect -146 -45838 -112 -45822
rect 112 -44646 146 -44630
rect 112 -45838 146 -45822
rect -100 -45915 -84 -45881
rect 84 -45915 100 -45881
rect -100 -46023 -84 -45989
rect 84 -46023 100 -45989
rect -146 -46082 -112 -46066
rect -146 -47274 -112 -47258
rect 112 -46082 146 -46066
rect 112 -47274 146 -47258
rect -100 -47351 -84 -47317
rect 84 -47351 100 -47317
rect -100 -47459 -84 -47425
rect 84 -47459 100 -47425
rect -146 -47518 -112 -47502
rect -146 -48710 -112 -48694
rect 112 -47518 146 -47502
rect 112 -48710 146 -48694
rect -100 -48787 -84 -48753
rect 84 -48787 100 -48753
rect -100 -48895 -84 -48861
rect 84 -48895 100 -48861
rect -146 -48954 -112 -48938
rect -146 -50146 -112 -50130
rect 112 -48954 146 -48938
rect 112 -50146 146 -50130
rect -100 -50223 -84 -50189
rect 84 -50223 100 -50189
rect -100 -50331 -84 -50297
rect 84 -50331 100 -50297
rect -146 -50390 -112 -50374
rect -146 -51582 -112 -51566
rect 112 -50390 146 -50374
rect 112 -51582 146 -51566
rect -100 -51659 -84 -51625
rect 84 -51659 100 -51625
rect -100 -51767 -84 -51733
rect 84 -51767 100 -51733
rect -146 -51826 -112 -51810
rect -146 -53018 -112 -53002
rect 112 -51826 146 -51810
rect 112 -53018 146 -53002
rect -100 -53095 -84 -53061
rect 84 -53095 100 -53061
rect -100 -53203 -84 -53169
rect 84 -53203 100 -53169
rect -146 -53262 -112 -53246
rect -146 -54454 -112 -54438
rect 112 -53262 146 -53246
rect 112 -54454 146 -54438
rect -100 -54531 -84 -54497
rect 84 -54531 100 -54497
rect -100 -54639 -84 -54605
rect 84 -54639 100 -54605
rect -146 -54698 -112 -54682
rect -146 -55890 -112 -55874
rect 112 -54698 146 -54682
rect 112 -55890 146 -55874
rect -100 -55967 -84 -55933
rect 84 -55967 100 -55933
rect -100 -56075 -84 -56041
rect 84 -56075 100 -56041
rect -146 -56134 -112 -56118
rect -146 -57326 -112 -57310
rect 112 -56134 146 -56118
rect 112 -57326 146 -57310
rect -100 -57403 -84 -57369
rect 84 -57403 100 -57369
rect -100 -57511 -84 -57477
rect 84 -57511 100 -57477
rect -146 -57570 -112 -57554
rect -146 -58762 -112 -58746
rect 112 -57570 146 -57554
rect 112 -58762 146 -58746
rect -100 -58839 -84 -58805
rect 84 -58839 100 -58805
rect -100 -58947 -84 -58913
rect 84 -58947 100 -58913
rect -146 -59006 -112 -58990
rect -146 -60198 -112 -60182
rect 112 -59006 146 -58990
rect 112 -60198 146 -60182
rect -100 -60275 -84 -60241
rect 84 -60275 100 -60241
rect -100 -60383 -84 -60349
rect 84 -60383 100 -60349
rect -146 -60442 -112 -60426
rect -146 -61634 -112 -61618
rect 112 -60442 146 -60426
rect 112 -61634 146 -61618
rect -100 -61711 -84 -61677
rect 84 -61711 100 -61677
rect -100 -61819 -84 -61785
rect 84 -61819 100 -61785
rect -146 -61878 -112 -61862
rect -146 -63070 -112 -63054
rect 112 -61878 146 -61862
rect 112 -63070 146 -63054
rect -100 -63147 -84 -63113
rect 84 -63147 100 -63113
rect -100 -63255 -84 -63221
rect 84 -63255 100 -63221
rect -146 -63314 -112 -63298
rect -146 -64506 -112 -64490
rect 112 -63314 146 -63298
rect 112 -64506 146 -64490
rect -100 -64583 -84 -64549
rect 84 -64583 100 -64549
rect -100 -64691 -84 -64657
rect 84 -64691 100 -64657
rect -146 -64750 -112 -64734
rect -146 -65942 -112 -65926
rect 112 -64750 146 -64734
rect 112 -65942 146 -65926
rect -100 -66019 -84 -65985
rect 84 -66019 100 -65985
rect -100 -66127 -84 -66093
rect 84 -66127 100 -66093
rect -146 -66186 -112 -66170
rect -146 -67378 -112 -67362
rect 112 -66186 146 -66170
rect 112 -67378 146 -67362
rect -100 -67455 -84 -67421
rect 84 -67455 100 -67421
rect -100 -67563 -84 -67529
rect 84 -67563 100 -67529
rect -146 -67622 -112 -67606
rect -146 -68814 -112 -68798
rect 112 -67622 146 -67606
rect 112 -68814 146 -68798
rect -100 -68891 -84 -68857
rect 84 -68891 100 -68857
rect -100 -68999 -84 -68965
rect 84 -68999 100 -68965
rect -146 -69058 -112 -69042
rect -146 -70250 -112 -70234
rect 112 -69058 146 -69042
rect 112 -70250 146 -70234
rect -100 -70327 -84 -70293
rect 84 -70327 100 -70293
rect -100 -70435 -84 -70401
rect 84 -70435 100 -70401
rect -146 -70494 -112 -70478
rect -146 -71686 -112 -71670
rect 112 -70494 146 -70478
rect 112 -71686 146 -71670
rect -100 -71763 -84 -71729
rect 84 -71763 100 -71729
rect -100 -71871 -84 -71837
rect 84 -71871 100 -71837
rect -146 -71930 -112 -71914
rect -146 -73122 -112 -73106
rect 112 -71930 146 -71914
rect 112 -73122 146 -73106
rect -100 -73199 -84 -73165
rect 84 -73199 100 -73165
rect -100 -73307 -84 -73273
rect 84 -73307 100 -73273
rect -146 -73366 -112 -73350
rect -146 -74558 -112 -74542
rect 112 -73366 146 -73350
rect 112 -74558 146 -74542
rect -100 -74635 -84 -74601
rect 84 -74635 100 -74601
rect -100 -74743 -84 -74709
rect 84 -74743 100 -74709
rect -146 -74802 -112 -74786
rect -146 -75994 -112 -75978
rect 112 -74802 146 -74786
rect 112 -75994 146 -75978
rect -100 -76071 -84 -76037
rect 84 -76071 100 -76037
rect -100 -76179 -84 -76145
rect 84 -76179 100 -76145
rect -146 -76238 -112 -76222
rect -146 -77430 -112 -77414
rect 112 -76238 146 -76222
rect 112 -77430 146 -77414
rect -100 -77507 -84 -77473
rect 84 -77507 100 -77473
rect -100 -77615 -84 -77581
rect 84 -77615 100 -77581
rect -146 -77674 -112 -77658
rect -146 -78866 -112 -78850
rect 112 -77674 146 -77658
rect 112 -78866 146 -78850
rect -100 -78943 -84 -78909
rect 84 -78943 100 -78909
rect -100 -79051 -84 -79017
rect 84 -79051 100 -79017
rect -146 -79110 -112 -79094
rect -146 -80302 -112 -80286
rect 112 -79110 146 -79094
rect 112 -80302 146 -80286
rect -100 -80379 -84 -80345
rect 84 -80379 100 -80345
rect -100 -80487 -84 -80453
rect 84 -80487 100 -80453
rect -146 -80546 -112 -80530
rect -146 -81738 -112 -81722
rect 112 -80546 146 -80530
rect 112 -81738 146 -81722
rect -100 -81815 -84 -81781
rect 84 -81815 100 -81781
rect -100 -81923 -84 -81889
rect 84 -81923 100 -81889
rect -146 -81982 -112 -81966
rect -146 -83174 -112 -83158
rect 112 -81982 146 -81966
rect 112 -83174 146 -83158
rect -100 -83251 -84 -83217
rect 84 -83251 100 -83217
rect -100 -83359 -84 -83325
rect 84 -83359 100 -83325
rect -146 -83418 -112 -83402
rect -146 -84610 -112 -84594
rect 112 -83418 146 -83402
rect 112 -84610 146 -84594
rect -100 -84687 -84 -84653
rect 84 -84687 100 -84653
rect -100 -84795 -84 -84761
rect 84 -84795 100 -84761
rect -146 -84854 -112 -84838
rect -146 -86046 -112 -86030
rect 112 -84854 146 -84838
rect 112 -86046 146 -86030
rect -100 -86123 -84 -86089
rect 84 -86123 100 -86089
rect -100 -86231 -84 -86197
rect 84 -86231 100 -86197
rect -146 -86290 -112 -86274
rect -146 -87482 -112 -87466
rect 112 -86290 146 -86274
rect 112 -87482 146 -87466
rect -100 -87559 -84 -87525
rect 84 -87559 100 -87525
rect -100 -87667 -84 -87633
rect 84 -87667 100 -87633
rect -146 -87726 -112 -87710
rect -146 -88918 -112 -88902
rect 112 -87726 146 -87710
rect 112 -88918 146 -88902
rect -100 -88995 -84 -88961
rect 84 -88995 100 -88961
rect -100 -89103 -84 -89069
rect 84 -89103 100 -89069
rect -146 -89162 -112 -89146
rect -146 -90354 -112 -90338
rect 112 -89162 146 -89146
rect 112 -90354 146 -90338
rect -100 -90431 -84 -90397
rect 84 -90431 100 -90397
rect -100 -90539 -84 -90505
rect 84 -90539 100 -90505
rect -146 -90598 -112 -90582
rect -146 -91790 -112 -91774
rect 112 -90598 146 -90582
rect 112 -91790 146 -91774
rect -100 -91867 -84 -91833
rect 84 -91867 100 -91833
rect -100 -91975 -84 -91941
rect 84 -91975 100 -91941
rect -146 -92034 -112 -92018
rect -146 -93226 -112 -93210
rect 112 -92034 146 -92018
rect 112 -93226 146 -93210
rect -100 -93303 -84 -93269
rect 84 -93303 100 -93269
rect -100 -93411 -84 -93377
rect 84 -93411 100 -93377
rect -146 -93470 -112 -93454
rect -146 -94662 -112 -94646
rect 112 -93470 146 -93454
rect 112 -94662 146 -94646
rect -100 -94739 -84 -94705
rect 84 -94739 100 -94705
rect -100 -94847 -84 -94813
rect 84 -94847 100 -94813
rect -146 -94906 -112 -94890
rect -146 -96098 -112 -96082
rect 112 -94906 146 -94890
rect 112 -96098 146 -96082
rect -100 -96175 -84 -96141
rect 84 -96175 100 -96141
rect -100 -96283 -84 -96249
rect 84 -96283 100 -96249
rect -146 -96342 -112 -96326
rect -146 -97534 -112 -97518
rect 112 -96342 146 -96326
rect 112 -97534 146 -97518
rect -100 -97611 -84 -97577
rect 84 -97611 100 -97577
rect -100 -97719 -84 -97685
rect 84 -97719 100 -97685
rect -146 -97778 -112 -97762
rect -146 -98970 -112 -98954
rect 112 -97778 146 -97762
rect 112 -98970 146 -98954
rect -100 -99047 -84 -99013
rect 84 -99047 100 -99013
rect -100 -99155 -84 -99121
rect 84 -99155 100 -99121
rect -146 -99214 -112 -99198
rect -146 -100406 -112 -100390
rect 112 -99214 146 -99198
rect 112 -100406 146 -100390
rect -100 -100483 -84 -100449
rect 84 -100483 100 -100449
rect -100 -100591 -84 -100557
rect 84 -100591 100 -100557
rect -146 -100650 -112 -100634
rect -146 -101842 -112 -101826
rect 112 -100650 146 -100634
rect 112 -101842 146 -101826
rect -100 -101919 -84 -101885
rect 84 -101919 100 -101885
rect -100 -102027 -84 -101993
rect 84 -102027 100 -101993
rect -146 -102086 -112 -102070
rect -146 -103278 -112 -103262
rect 112 -102086 146 -102070
rect 112 -103278 146 -103262
rect -100 -103355 -84 -103321
rect 84 -103355 100 -103321
rect -100 -103463 -84 -103429
rect 84 -103463 100 -103429
rect -146 -103522 -112 -103506
rect -146 -104714 -112 -104698
rect 112 -103522 146 -103506
rect 112 -104714 146 -104698
rect -100 -104791 -84 -104757
rect 84 -104791 100 -104757
rect -100 -104899 -84 -104865
rect 84 -104899 100 -104865
rect -146 -104958 -112 -104942
rect -146 -106150 -112 -106134
rect 112 -104958 146 -104942
rect 112 -106150 146 -106134
rect -100 -106227 -84 -106193
rect 84 -106227 100 -106193
rect -100 -106335 -84 -106301
rect 84 -106335 100 -106301
rect -146 -106394 -112 -106378
rect -146 -107586 -112 -107570
rect 112 -106394 146 -106378
rect 112 -107586 146 -107570
rect -100 -107663 -84 -107629
rect 84 -107663 100 -107629
rect -100 -107771 -84 -107737
rect 84 -107771 100 -107737
rect -146 -107830 -112 -107814
rect -146 -109022 -112 -109006
rect 112 -107830 146 -107814
rect 112 -109022 146 -109006
rect -100 -109099 -84 -109065
rect 84 -109099 100 -109065
rect -100 -109207 -84 -109173
rect 84 -109207 100 -109173
rect -146 -109266 -112 -109250
rect -146 -110458 -112 -110442
rect 112 -109266 146 -109250
rect 112 -110458 146 -110442
rect -100 -110535 -84 -110501
rect 84 -110535 100 -110501
rect -100 -110643 -84 -110609
rect 84 -110643 100 -110609
rect -146 -110702 -112 -110686
rect -146 -111894 -112 -111878
rect 112 -110702 146 -110686
rect 112 -111894 146 -111878
rect -100 -111971 -84 -111937
rect 84 -111971 100 -111937
rect -100 -112079 -84 -112045
rect 84 -112079 100 -112045
rect -146 -112138 -112 -112122
rect -146 -113330 -112 -113314
rect 112 -112138 146 -112122
rect 112 -113330 146 -113314
rect -100 -113407 -84 -113373
rect 84 -113407 100 -113373
rect -100 -113515 -84 -113481
rect 84 -113515 100 -113481
rect -146 -113574 -112 -113558
rect -146 -114766 -112 -114750
rect 112 -113574 146 -113558
rect 112 -114766 146 -114750
rect -100 -114843 -84 -114809
rect 84 -114843 100 -114809
rect -100 -114951 -84 -114917
rect 84 -114951 100 -114917
rect -146 -115010 -112 -114994
rect -146 -116202 -112 -116186
rect 112 -115010 146 -114994
rect 112 -116202 146 -116186
rect -100 -116279 -84 -116245
rect 84 -116279 100 -116245
rect -100 -116387 -84 -116353
rect 84 -116387 100 -116353
rect -146 -116446 -112 -116430
rect -146 -117638 -112 -117622
rect 112 -116446 146 -116430
rect 112 -117638 146 -117622
rect -100 -117715 -84 -117681
rect 84 -117715 100 -117681
rect -100 -117823 -84 -117789
rect 84 -117823 100 -117789
rect -146 -117882 -112 -117866
rect -146 -119074 -112 -119058
rect 112 -117882 146 -117866
rect 112 -119074 146 -119058
rect -100 -119151 -84 -119117
rect 84 -119151 100 -119117
rect -100 -119259 -84 -119225
rect 84 -119259 100 -119225
rect -146 -119318 -112 -119302
rect -146 -120510 -112 -120494
rect 112 -119318 146 -119302
rect 112 -120510 146 -120494
rect -100 -120587 -84 -120553
rect 84 -120587 100 -120553
rect -100 -120695 -84 -120661
rect 84 -120695 100 -120661
rect -146 -120754 -112 -120738
rect -146 -121946 -112 -121930
rect 112 -120754 146 -120738
rect 112 -121946 146 -121930
rect -100 -122023 -84 -121989
rect 84 -122023 100 -121989
rect -100 -122131 -84 -122097
rect 84 -122131 100 -122097
rect -146 -122190 -112 -122174
rect -146 -123382 -112 -123366
rect 112 -122190 146 -122174
rect 112 -123382 146 -123366
rect -100 -123459 -84 -123425
rect 84 -123459 100 -123425
rect -100 -123567 -84 -123533
rect 84 -123567 100 -123533
rect -146 -123626 -112 -123610
rect -146 -124818 -112 -124802
rect 112 -123626 146 -123610
rect 112 -124818 146 -124802
rect -100 -124895 -84 -124861
rect 84 -124895 100 -124861
rect -100 -125003 -84 -124969
rect 84 -125003 100 -124969
rect -146 -125062 -112 -125046
rect -146 -126254 -112 -126238
rect 112 -125062 146 -125046
rect 112 -126254 146 -126238
rect -100 -126331 -84 -126297
rect 84 -126331 100 -126297
rect -100 -126439 -84 -126405
rect 84 -126439 100 -126405
rect -146 -126498 -112 -126482
rect -146 -127690 -112 -127674
rect 112 -126498 146 -126482
rect 112 -127690 146 -127674
rect -100 -127767 -84 -127733
rect 84 -127767 100 -127733
rect -100 -127875 -84 -127841
rect 84 -127875 100 -127841
rect -146 -127934 -112 -127918
rect -146 -129126 -112 -129110
rect 112 -127934 146 -127918
rect 112 -129126 146 -129110
rect -100 -129203 -84 -129169
rect 84 -129203 100 -129169
rect -100 -129311 -84 -129277
rect 84 -129311 100 -129277
rect -146 -129370 -112 -129354
rect -146 -130562 -112 -130546
rect 112 -129370 146 -129354
rect 112 -130562 146 -130546
rect -100 -130639 -84 -130605
rect 84 -130639 100 -130605
rect -100 -130747 -84 -130713
rect 84 -130747 100 -130713
rect -146 -130806 -112 -130790
rect -146 -131998 -112 -131982
rect 112 -130806 146 -130790
rect 112 -131998 146 -131982
rect -100 -132075 -84 -132041
rect 84 -132075 100 -132041
rect -100 -132183 -84 -132149
rect 84 -132183 100 -132149
rect -146 -132242 -112 -132226
rect -146 -133434 -112 -133418
rect 112 -132242 146 -132226
rect 112 -133434 146 -133418
rect -100 -133511 -84 -133477
rect 84 -133511 100 -133477
rect -100 -133619 -84 -133585
rect 84 -133619 100 -133585
rect -146 -133678 -112 -133662
rect -146 -134870 -112 -134854
rect 112 -133678 146 -133662
rect 112 -134870 146 -134854
rect -100 -134947 -84 -134913
rect 84 -134947 100 -134913
rect -100 -135055 -84 -135021
rect 84 -135055 100 -135021
rect -146 -135114 -112 -135098
rect -146 -136306 -112 -136290
rect 112 -135114 146 -135098
rect 112 -136306 146 -136290
rect -100 -136383 -84 -136349
rect 84 -136383 100 -136349
rect -100 -136491 -84 -136457
rect 84 -136491 100 -136457
rect -146 -136550 -112 -136534
rect -146 -137742 -112 -137726
rect 112 -136550 146 -136534
rect 112 -137742 146 -137726
rect -100 -137819 -84 -137785
rect 84 -137819 100 -137785
rect -100 -137927 -84 -137893
rect 84 -137927 100 -137893
rect -146 -137986 -112 -137970
rect -146 -139178 -112 -139162
rect 112 -137986 146 -137970
rect 112 -139178 146 -139162
rect -100 -139255 -84 -139221
rect 84 -139255 100 -139221
rect -100 -139363 -84 -139329
rect 84 -139363 100 -139329
rect -146 -139422 -112 -139406
rect -146 -140614 -112 -140598
rect 112 -139422 146 -139406
rect 112 -140614 146 -140598
rect -100 -140691 -84 -140657
rect 84 -140691 100 -140657
rect -100 -140799 -84 -140765
rect 84 -140799 100 -140765
rect -146 -140858 -112 -140842
rect -146 -142050 -112 -142034
rect 112 -140858 146 -140842
rect 112 -142050 146 -142034
rect -100 -142127 -84 -142093
rect 84 -142127 100 -142093
rect -100 -142235 -84 -142201
rect 84 -142235 100 -142201
rect -146 -142294 -112 -142278
rect -146 -143486 -112 -143470
rect 112 -142294 146 -142278
rect 112 -143486 146 -143470
rect -100 -143563 -84 -143529
rect 84 -143563 100 -143529
rect -100 -143671 -84 -143637
rect 84 -143671 100 -143637
rect -146 -143730 -112 -143714
rect -146 -144922 -112 -144906
rect 112 -143730 146 -143714
rect 112 -144922 146 -144906
rect -100 -144999 -84 -144965
rect 84 -144999 100 -144965
rect -100 -145107 -84 -145073
rect 84 -145107 100 -145073
rect -146 -145166 -112 -145150
rect -146 -146358 -112 -146342
rect 112 -145166 146 -145150
rect 112 -146358 146 -146342
rect -100 -146435 -84 -146401
rect 84 -146435 100 -146401
rect -100 -146543 -84 -146509
rect 84 -146543 100 -146509
rect -146 -146602 -112 -146586
rect -146 -147794 -112 -147778
rect 112 -146602 146 -146586
rect 112 -147794 146 -147778
rect -100 -147871 -84 -147837
rect 84 -147871 100 -147837
rect -100 -147979 -84 -147945
rect 84 -147979 100 -147945
rect -146 -148038 -112 -148022
rect -146 -149230 -112 -149214
rect 112 -148038 146 -148022
rect 112 -149230 146 -149214
rect -100 -149307 -84 -149273
rect 84 -149307 100 -149273
rect -100 -149415 -84 -149381
rect 84 -149415 100 -149381
rect -146 -149474 -112 -149458
rect -146 -150666 -112 -150650
rect 112 -149474 146 -149458
rect 112 -150666 146 -150650
rect -100 -150743 -84 -150709
rect 84 -150743 100 -150709
rect -100 -150851 -84 -150817
rect 84 -150851 100 -150817
rect -146 -150910 -112 -150894
rect -146 -152102 -112 -152086
rect 112 -150910 146 -150894
rect 112 -152102 146 -152086
rect -100 -152179 -84 -152145
rect 84 -152179 100 -152145
rect -100 -152287 -84 -152253
rect 84 -152287 100 -152253
rect -146 -152346 -112 -152330
rect -146 -153538 -112 -153522
rect 112 -152346 146 -152330
rect 112 -153538 146 -153522
rect -100 -153615 -84 -153581
rect 84 -153615 100 -153581
rect -100 -153723 -84 -153689
rect 84 -153723 100 -153689
rect -146 -153782 -112 -153766
rect -146 -154974 -112 -154958
rect 112 -153782 146 -153766
rect 112 -154974 146 -154958
rect -100 -155051 -84 -155017
rect 84 -155051 100 -155017
rect -100 -155159 -84 -155125
rect 84 -155159 100 -155125
rect -146 -155218 -112 -155202
rect -146 -156410 -112 -156394
rect 112 -155218 146 -155202
rect 112 -156410 146 -156394
rect -100 -156487 -84 -156453
rect 84 -156487 100 -156453
rect -100 -156595 -84 -156561
rect 84 -156595 100 -156561
rect -146 -156654 -112 -156638
rect -146 -157846 -112 -157830
rect 112 -156654 146 -156638
rect 112 -157846 146 -157830
rect -100 -157923 -84 -157889
rect 84 -157923 100 -157889
rect -100 -158031 -84 -157997
rect 84 -158031 100 -157997
rect -146 -158090 -112 -158074
rect -146 -159282 -112 -159266
rect 112 -158090 146 -158074
rect 112 -159282 146 -159266
rect -100 -159359 -84 -159325
rect 84 -159359 100 -159325
rect -100 -159467 -84 -159433
rect 84 -159467 100 -159433
rect -146 -159526 -112 -159510
rect -146 -160718 -112 -160702
rect 112 -159526 146 -159510
rect 112 -160718 146 -160702
rect -100 -160795 -84 -160761
rect 84 -160795 100 -160761
rect -100 -160903 -84 -160869
rect 84 -160903 100 -160869
rect -146 -160962 -112 -160946
rect -146 -162154 -112 -162138
rect 112 -160962 146 -160946
rect 112 -162154 146 -162138
rect -100 -162231 -84 -162197
rect 84 -162231 100 -162197
rect -100 -162339 -84 -162305
rect 84 -162339 100 -162305
rect -146 -162398 -112 -162382
rect -146 -163590 -112 -163574
rect 112 -162398 146 -162382
rect 112 -163590 146 -163574
rect -100 -163667 -84 -163633
rect 84 -163667 100 -163633
rect -100 -163775 -84 -163741
rect 84 -163775 100 -163741
rect -146 -163834 -112 -163818
rect -146 -165026 -112 -165010
rect 112 -163834 146 -163818
rect 112 -165026 146 -165010
rect -100 -165103 -84 -165069
rect 84 -165103 100 -165069
rect -100 -165211 -84 -165177
rect 84 -165211 100 -165177
rect -146 -165270 -112 -165254
rect -146 -166462 -112 -166446
rect 112 -165270 146 -165254
rect 112 -166462 146 -166446
rect -100 -166539 -84 -166505
rect 84 -166539 100 -166505
rect -100 -166647 -84 -166613
rect 84 -166647 100 -166613
rect -146 -166706 -112 -166690
rect -146 -167898 -112 -167882
rect 112 -166706 146 -166690
rect 112 -167898 146 -167882
rect -100 -167975 -84 -167941
rect 84 -167975 100 -167941
rect -100 -168083 -84 -168049
rect 84 -168083 100 -168049
rect -146 -168142 -112 -168126
rect -146 -169334 -112 -169318
rect 112 -168142 146 -168126
rect 112 -169334 146 -169318
rect -100 -169411 -84 -169377
rect 84 -169411 100 -169377
rect -100 -169519 -84 -169485
rect 84 -169519 100 -169485
rect -146 -169578 -112 -169562
rect -146 -170770 -112 -170754
rect 112 -169578 146 -169562
rect 112 -170770 146 -170754
rect -100 -170847 -84 -170813
rect 84 -170847 100 -170813
rect -100 -170955 -84 -170921
rect 84 -170955 100 -170921
rect -146 -171014 -112 -170998
rect -146 -172206 -112 -172190
rect 112 -171014 146 -170998
rect 112 -172206 146 -172190
rect -100 -172283 -84 -172249
rect 84 -172283 100 -172249
rect -100 -172391 -84 -172357
rect 84 -172391 100 -172357
rect -146 -172450 -112 -172434
rect -146 -173642 -112 -173626
rect 112 -172450 146 -172434
rect 112 -173642 146 -173626
rect -100 -173719 -84 -173685
rect 84 -173719 100 -173685
rect -100 -173827 -84 -173793
rect 84 -173827 100 -173793
rect -146 -173886 -112 -173870
rect -146 -175078 -112 -175062
rect 112 -173886 146 -173870
rect 112 -175078 146 -175062
rect -100 -175155 -84 -175121
rect 84 -175155 100 -175121
rect -100 -175263 -84 -175229
rect 84 -175263 100 -175229
rect -146 -175322 -112 -175306
rect -146 -176514 -112 -176498
rect 112 -175322 146 -175306
rect 112 -176514 146 -176498
rect -100 -176591 -84 -176557
rect 84 -176591 100 -176557
rect -100 -176699 -84 -176665
rect 84 -176699 100 -176665
rect -146 -176758 -112 -176742
rect -146 -177950 -112 -177934
rect 112 -176758 146 -176742
rect 112 -177950 146 -177934
rect -100 -178027 -84 -177993
rect 84 -178027 100 -177993
rect -100 -178135 -84 -178101
rect 84 -178135 100 -178101
rect -146 -178194 -112 -178178
rect -146 -179386 -112 -179370
rect 112 -178194 146 -178178
rect 112 -179386 146 -179370
rect -100 -179463 -84 -179429
rect 84 -179463 100 -179429
rect -100 -179571 -84 -179537
rect 84 -179571 100 -179537
rect -146 -179630 -112 -179614
rect -146 -180822 -112 -180806
rect 112 -179630 146 -179614
rect 112 -180822 146 -180806
rect -100 -180899 -84 -180865
rect 84 -180899 100 -180865
rect -100 -181007 -84 -180973
rect 84 -181007 100 -180973
rect -146 -181066 -112 -181050
rect -146 -182258 -112 -182242
rect 112 -181066 146 -181050
rect 112 -182258 146 -182242
rect -100 -182335 -84 -182301
rect 84 -182335 100 -182301
rect -100 -182443 -84 -182409
rect 84 -182443 100 -182409
rect -146 -182502 -112 -182486
rect -146 -183694 -112 -183678
rect 112 -182502 146 -182486
rect 112 -183694 146 -183678
rect -100 -183771 -84 -183737
rect 84 -183771 100 -183737
rect -280 -183875 -246 -183813
rect 246 -183875 280 -183813
rect -280 -183909 -184 -183875
rect 184 -183909 280 -183875
<< viali >>
rect -84 183737 84 183771
rect -146 182502 -112 183678
rect 112 182502 146 183678
rect -84 182409 84 182443
rect -84 182301 84 182335
rect -146 181066 -112 182242
rect 112 181066 146 182242
rect -84 180973 84 181007
rect -84 180865 84 180899
rect -146 179630 -112 180806
rect 112 179630 146 180806
rect -84 179537 84 179571
rect -84 179429 84 179463
rect -146 178194 -112 179370
rect 112 178194 146 179370
rect -84 178101 84 178135
rect -84 177993 84 178027
rect -146 176758 -112 177934
rect 112 176758 146 177934
rect -84 176665 84 176699
rect -84 176557 84 176591
rect -146 175322 -112 176498
rect 112 175322 146 176498
rect -84 175229 84 175263
rect -84 175121 84 175155
rect -146 173886 -112 175062
rect 112 173886 146 175062
rect -84 173793 84 173827
rect -84 173685 84 173719
rect -146 172450 -112 173626
rect 112 172450 146 173626
rect -84 172357 84 172391
rect -84 172249 84 172283
rect -146 171014 -112 172190
rect 112 171014 146 172190
rect -84 170921 84 170955
rect -84 170813 84 170847
rect -146 169578 -112 170754
rect 112 169578 146 170754
rect -84 169485 84 169519
rect -84 169377 84 169411
rect -146 168142 -112 169318
rect 112 168142 146 169318
rect -84 168049 84 168083
rect -84 167941 84 167975
rect -146 166706 -112 167882
rect 112 166706 146 167882
rect -84 166613 84 166647
rect -84 166505 84 166539
rect -146 165270 -112 166446
rect 112 165270 146 166446
rect -84 165177 84 165211
rect -84 165069 84 165103
rect -146 163834 -112 165010
rect 112 163834 146 165010
rect -84 163741 84 163775
rect -84 163633 84 163667
rect -146 162398 -112 163574
rect 112 162398 146 163574
rect -84 162305 84 162339
rect -84 162197 84 162231
rect -146 160962 -112 162138
rect 112 160962 146 162138
rect -84 160869 84 160903
rect -84 160761 84 160795
rect -146 159526 -112 160702
rect 112 159526 146 160702
rect -84 159433 84 159467
rect -84 159325 84 159359
rect -146 158090 -112 159266
rect 112 158090 146 159266
rect -84 157997 84 158031
rect -84 157889 84 157923
rect -146 156654 -112 157830
rect 112 156654 146 157830
rect -84 156561 84 156595
rect -84 156453 84 156487
rect -146 155218 -112 156394
rect 112 155218 146 156394
rect -84 155125 84 155159
rect -84 155017 84 155051
rect -146 153782 -112 154958
rect 112 153782 146 154958
rect -84 153689 84 153723
rect -84 153581 84 153615
rect -146 152346 -112 153522
rect 112 152346 146 153522
rect -84 152253 84 152287
rect -84 152145 84 152179
rect -146 150910 -112 152086
rect 112 150910 146 152086
rect -84 150817 84 150851
rect -84 150709 84 150743
rect -146 149474 -112 150650
rect 112 149474 146 150650
rect -84 149381 84 149415
rect -84 149273 84 149307
rect -146 148038 -112 149214
rect 112 148038 146 149214
rect -84 147945 84 147979
rect -84 147837 84 147871
rect -146 146602 -112 147778
rect 112 146602 146 147778
rect -84 146509 84 146543
rect -84 146401 84 146435
rect -146 145166 -112 146342
rect 112 145166 146 146342
rect -84 145073 84 145107
rect -84 144965 84 144999
rect -146 143730 -112 144906
rect 112 143730 146 144906
rect -84 143637 84 143671
rect -84 143529 84 143563
rect -146 142294 -112 143470
rect 112 142294 146 143470
rect -84 142201 84 142235
rect -84 142093 84 142127
rect -146 140858 -112 142034
rect 112 140858 146 142034
rect -84 140765 84 140799
rect -84 140657 84 140691
rect -146 139422 -112 140598
rect 112 139422 146 140598
rect -84 139329 84 139363
rect -84 139221 84 139255
rect -146 137986 -112 139162
rect 112 137986 146 139162
rect -84 137893 84 137927
rect -84 137785 84 137819
rect -146 136550 -112 137726
rect 112 136550 146 137726
rect -84 136457 84 136491
rect -84 136349 84 136383
rect -146 135114 -112 136290
rect 112 135114 146 136290
rect -84 135021 84 135055
rect -84 134913 84 134947
rect -146 133678 -112 134854
rect 112 133678 146 134854
rect -84 133585 84 133619
rect -84 133477 84 133511
rect -146 132242 -112 133418
rect 112 132242 146 133418
rect -84 132149 84 132183
rect -84 132041 84 132075
rect -146 130806 -112 131982
rect 112 130806 146 131982
rect -84 130713 84 130747
rect -84 130605 84 130639
rect -146 129370 -112 130546
rect 112 129370 146 130546
rect -84 129277 84 129311
rect -84 129169 84 129203
rect -146 127934 -112 129110
rect 112 127934 146 129110
rect -84 127841 84 127875
rect -84 127733 84 127767
rect -146 126498 -112 127674
rect 112 126498 146 127674
rect -84 126405 84 126439
rect -84 126297 84 126331
rect -146 125062 -112 126238
rect 112 125062 146 126238
rect -84 124969 84 125003
rect -84 124861 84 124895
rect -146 123626 -112 124802
rect 112 123626 146 124802
rect -84 123533 84 123567
rect -84 123425 84 123459
rect -146 122190 -112 123366
rect 112 122190 146 123366
rect -84 122097 84 122131
rect -84 121989 84 122023
rect -146 120754 -112 121930
rect 112 120754 146 121930
rect -84 120661 84 120695
rect -84 120553 84 120587
rect -146 119318 -112 120494
rect 112 119318 146 120494
rect -84 119225 84 119259
rect -84 119117 84 119151
rect -146 117882 -112 119058
rect 112 117882 146 119058
rect -84 117789 84 117823
rect -84 117681 84 117715
rect -146 116446 -112 117622
rect 112 116446 146 117622
rect -84 116353 84 116387
rect -84 116245 84 116279
rect -146 115010 -112 116186
rect 112 115010 146 116186
rect -84 114917 84 114951
rect -84 114809 84 114843
rect -146 113574 -112 114750
rect 112 113574 146 114750
rect -84 113481 84 113515
rect -84 113373 84 113407
rect -146 112138 -112 113314
rect 112 112138 146 113314
rect -84 112045 84 112079
rect -84 111937 84 111971
rect -146 110702 -112 111878
rect 112 110702 146 111878
rect -84 110609 84 110643
rect -84 110501 84 110535
rect -146 109266 -112 110442
rect 112 109266 146 110442
rect -84 109173 84 109207
rect -84 109065 84 109099
rect -146 107830 -112 109006
rect 112 107830 146 109006
rect -84 107737 84 107771
rect -84 107629 84 107663
rect -146 106394 -112 107570
rect 112 106394 146 107570
rect -84 106301 84 106335
rect -84 106193 84 106227
rect -146 104958 -112 106134
rect 112 104958 146 106134
rect -84 104865 84 104899
rect -84 104757 84 104791
rect -146 103522 -112 104698
rect 112 103522 146 104698
rect -84 103429 84 103463
rect -84 103321 84 103355
rect -146 102086 -112 103262
rect 112 102086 146 103262
rect -84 101993 84 102027
rect -84 101885 84 101919
rect -146 100650 -112 101826
rect 112 100650 146 101826
rect -84 100557 84 100591
rect -84 100449 84 100483
rect -146 99214 -112 100390
rect 112 99214 146 100390
rect -84 99121 84 99155
rect -84 99013 84 99047
rect -146 97778 -112 98954
rect 112 97778 146 98954
rect -84 97685 84 97719
rect -84 97577 84 97611
rect -146 96342 -112 97518
rect 112 96342 146 97518
rect -84 96249 84 96283
rect -84 96141 84 96175
rect -146 94906 -112 96082
rect 112 94906 146 96082
rect -84 94813 84 94847
rect -84 94705 84 94739
rect -146 93470 -112 94646
rect 112 93470 146 94646
rect -84 93377 84 93411
rect -84 93269 84 93303
rect -146 92034 -112 93210
rect 112 92034 146 93210
rect -84 91941 84 91975
rect -84 91833 84 91867
rect -146 90598 -112 91774
rect 112 90598 146 91774
rect -84 90505 84 90539
rect -84 90397 84 90431
rect -146 89162 -112 90338
rect 112 89162 146 90338
rect -84 89069 84 89103
rect -84 88961 84 88995
rect -146 87726 -112 88902
rect 112 87726 146 88902
rect -84 87633 84 87667
rect -84 87525 84 87559
rect -146 86290 -112 87466
rect 112 86290 146 87466
rect -84 86197 84 86231
rect -84 86089 84 86123
rect -146 84854 -112 86030
rect 112 84854 146 86030
rect -84 84761 84 84795
rect -84 84653 84 84687
rect -146 83418 -112 84594
rect 112 83418 146 84594
rect -84 83325 84 83359
rect -84 83217 84 83251
rect -146 81982 -112 83158
rect 112 81982 146 83158
rect -84 81889 84 81923
rect -84 81781 84 81815
rect -146 80546 -112 81722
rect 112 80546 146 81722
rect -84 80453 84 80487
rect -84 80345 84 80379
rect -146 79110 -112 80286
rect 112 79110 146 80286
rect -84 79017 84 79051
rect -84 78909 84 78943
rect -146 77674 -112 78850
rect 112 77674 146 78850
rect -84 77581 84 77615
rect -84 77473 84 77507
rect -146 76238 -112 77414
rect 112 76238 146 77414
rect -84 76145 84 76179
rect -84 76037 84 76071
rect -146 74802 -112 75978
rect 112 74802 146 75978
rect -84 74709 84 74743
rect -84 74601 84 74635
rect -146 73366 -112 74542
rect 112 73366 146 74542
rect -84 73273 84 73307
rect -84 73165 84 73199
rect -146 71930 -112 73106
rect 112 71930 146 73106
rect -84 71837 84 71871
rect -84 71729 84 71763
rect -146 70494 -112 71670
rect 112 70494 146 71670
rect -84 70401 84 70435
rect -84 70293 84 70327
rect -146 69058 -112 70234
rect 112 69058 146 70234
rect -84 68965 84 68999
rect -84 68857 84 68891
rect -146 67622 -112 68798
rect 112 67622 146 68798
rect -84 67529 84 67563
rect -84 67421 84 67455
rect -146 66186 -112 67362
rect 112 66186 146 67362
rect -84 66093 84 66127
rect -84 65985 84 66019
rect -146 64750 -112 65926
rect 112 64750 146 65926
rect -84 64657 84 64691
rect -84 64549 84 64583
rect -146 63314 -112 64490
rect 112 63314 146 64490
rect -84 63221 84 63255
rect -84 63113 84 63147
rect -146 61878 -112 63054
rect 112 61878 146 63054
rect -84 61785 84 61819
rect -84 61677 84 61711
rect -146 60442 -112 61618
rect 112 60442 146 61618
rect -84 60349 84 60383
rect -84 60241 84 60275
rect -146 59006 -112 60182
rect 112 59006 146 60182
rect -84 58913 84 58947
rect -84 58805 84 58839
rect -146 57570 -112 58746
rect 112 57570 146 58746
rect -84 57477 84 57511
rect -84 57369 84 57403
rect -146 56134 -112 57310
rect 112 56134 146 57310
rect -84 56041 84 56075
rect -84 55933 84 55967
rect -146 54698 -112 55874
rect 112 54698 146 55874
rect -84 54605 84 54639
rect -84 54497 84 54531
rect -146 53262 -112 54438
rect 112 53262 146 54438
rect -84 53169 84 53203
rect -84 53061 84 53095
rect -146 51826 -112 53002
rect 112 51826 146 53002
rect -84 51733 84 51767
rect -84 51625 84 51659
rect -146 50390 -112 51566
rect 112 50390 146 51566
rect -84 50297 84 50331
rect -84 50189 84 50223
rect -146 48954 -112 50130
rect 112 48954 146 50130
rect -84 48861 84 48895
rect -84 48753 84 48787
rect -146 47518 -112 48694
rect 112 47518 146 48694
rect -84 47425 84 47459
rect -84 47317 84 47351
rect -146 46082 -112 47258
rect 112 46082 146 47258
rect -84 45989 84 46023
rect -84 45881 84 45915
rect -146 44646 -112 45822
rect 112 44646 146 45822
rect -84 44553 84 44587
rect -84 44445 84 44479
rect -146 43210 -112 44386
rect 112 43210 146 44386
rect -84 43117 84 43151
rect -84 43009 84 43043
rect -146 41774 -112 42950
rect 112 41774 146 42950
rect -84 41681 84 41715
rect -84 41573 84 41607
rect -146 40338 -112 41514
rect 112 40338 146 41514
rect -84 40245 84 40279
rect -84 40137 84 40171
rect -146 38902 -112 40078
rect 112 38902 146 40078
rect -84 38809 84 38843
rect -84 38701 84 38735
rect -146 37466 -112 38642
rect 112 37466 146 38642
rect -84 37373 84 37407
rect -84 37265 84 37299
rect -146 36030 -112 37206
rect 112 36030 146 37206
rect -84 35937 84 35971
rect -84 35829 84 35863
rect -146 34594 -112 35770
rect 112 34594 146 35770
rect -84 34501 84 34535
rect -84 34393 84 34427
rect -146 33158 -112 34334
rect 112 33158 146 34334
rect -84 33065 84 33099
rect -84 32957 84 32991
rect -146 31722 -112 32898
rect 112 31722 146 32898
rect -84 31629 84 31663
rect -84 31521 84 31555
rect -146 30286 -112 31462
rect 112 30286 146 31462
rect -84 30193 84 30227
rect -84 30085 84 30119
rect -146 28850 -112 30026
rect 112 28850 146 30026
rect -84 28757 84 28791
rect -84 28649 84 28683
rect -146 27414 -112 28590
rect 112 27414 146 28590
rect -84 27321 84 27355
rect -84 27213 84 27247
rect -146 25978 -112 27154
rect 112 25978 146 27154
rect -84 25885 84 25919
rect -84 25777 84 25811
rect -146 24542 -112 25718
rect 112 24542 146 25718
rect -84 24449 84 24483
rect -84 24341 84 24375
rect -146 23106 -112 24282
rect 112 23106 146 24282
rect -84 23013 84 23047
rect -84 22905 84 22939
rect -146 21670 -112 22846
rect 112 21670 146 22846
rect -84 21577 84 21611
rect -84 21469 84 21503
rect -146 20234 -112 21410
rect 112 20234 146 21410
rect -84 20141 84 20175
rect -84 20033 84 20067
rect -146 18798 -112 19974
rect 112 18798 146 19974
rect -84 18705 84 18739
rect -84 18597 84 18631
rect -146 17362 -112 18538
rect 112 17362 146 18538
rect -84 17269 84 17303
rect -84 17161 84 17195
rect -146 15926 -112 17102
rect 112 15926 146 17102
rect -84 15833 84 15867
rect -84 15725 84 15759
rect -146 14490 -112 15666
rect 112 14490 146 15666
rect -84 14397 84 14431
rect -84 14289 84 14323
rect -146 13054 -112 14230
rect 112 13054 146 14230
rect -84 12961 84 12995
rect -84 12853 84 12887
rect -146 11618 -112 12794
rect 112 11618 146 12794
rect -84 11525 84 11559
rect -84 11417 84 11451
rect -146 10182 -112 11358
rect 112 10182 146 11358
rect -84 10089 84 10123
rect -84 9981 84 10015
rect -146 8746 -112 9922
rect 112 8746 146 9922
rect -84 8653 84 8687
rect -84 8545 84 8579
rect -146 7310 -112 8486
rect 112 7310 146 8486
rect -84 7217 84 7251
rect -84 7109 84 7143
rect -146 5874 -112 7050
rect 112 5874 146 7050
rect -84 5781 84 5815
rect -84 5673 84 5707
rect -146 4438 -112 5614
rect 112 4438 146 5614
rect -84 4345 84 4379
rect -84 4237 84 4271
rect -146 3002 -112 4178
rect 112 3002 146 4178
rect -84 2909 84 2943
rect -84 2801 84 2835
rect -146 1566 -112 2742
rect 112 1566 146 2742
rect -84 1473 84 1507
rect -84 1365 84 1399
rect -146 130 -112 1306
rect 112 130 146 1306
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1306 -112 -130
rect 112 -1306 146 -130
rect -84 -1399 84 -1365
rect -84 -1507 84 -1473
rect -146 -2742 -112 -1566
rect 112 -2742 146 -1566
rect -84 -2835 84 -2801
rect -84 -2943 84 -2909
rect -146 -4178 -112 -3002
rect 112 -4178 146 -3002
rect -84 -4271 84 -4237
rect -84 -4379 84 -4345
rect -146 -5614 -112 -4438
rect 112 -5614 146 -4438
rect -84 -5707 84 -5673
rect -84 -5815 84 -5781
rect -146 -7050 -112 -5874
rect 112 -7050 146 -5874
rect -84 -7143 84 -7109
rect -84 -7251 84 -7217
rect -146 -8486 -112 -7310
rect 112 -8486 146 -7310
rect -84 -8579 84 -8545
rect -84 -8687 84 -8653
rect -146 -9922 -112 -8746
rect 112 -9922 146 -8746
rect -84 -10015 84 -9981
rect -84 -10123 84 -10089
rect -146 -11358 -112 -10182
rect 112 -11358 146 -10182
rect -84 -11451 84 -11417
rect -84 -11559 84 -11525
rect -146 -12794 -112 -11618
rect 112 -12794 146 -11618
rect -84 -12887 84 -12853
rect -84 -12995 84 -12961
rect -146 -14230 -112 -13054
rect 112 -14230 146 -13054
rect -84 -14323 84 -14289
rect -84 -14431 84 -14397
rect -146 -15666 -112 -14490
rect 112 -15666 146 -14490
rect -84 -15759 84 -15725
rect -84 -15867 84 -15833
rect -146 -17102 -112 -15926
rect 112 -17102 146 -15926
rect -84 -17195 84 -17161
rect -84 -17303 84 -17269
rect -146 -18538 -112 -17362
rect 112 -18538 146 -17362
rect -84 -18631 84 -18597
rect -84 -18739 84 -18705
rect -146 -19974 -112 -18798
rect 112 -19974 146 -18798
rect -84 -20067 84 -20033
rect -84 -20175 84 -20141
rect -146 -21410 -112 -20234
rect 112 -21410 146 -20234
rect -84 -21503 84 -21469
rect -84 -21611 84 -21577
rect -146 -22846 -112 -21670
rect 112 -22846 146 -21670
rect -84 -22939 84 -22905
rect -84 -23047 84 -23013
rect -146 -24282 -112 -23106
rect 112 -24282 146 -23106
rect -84 -24375 84 -24341
rect -84 -24483 84 -24449
rect -146 -25718 -112 -24542
rect 112 -25718 146 -24542
rect -84 -25811 84 -25777
rect -84 -25919 84 -25885
rect -146 -27154 -112 -25978
rect 112 -27154 146 -25978
rect -84 -27247 84 -27213
rect -84 -27355 84 -27321
rect -146 -28590 -112 -27414
rect 112 -28590 146 -27414
rect -84 -28683 84 -28649
rect -84 -28791 84 -28757
rect -146 -30026 -112 -28850
rect 112 -30026 146 -28850
rect -84 -30119 84 -30085
rect -84 -30227 84 -30193
rect -146 -31462 -112 -30286
rect 112 -31462 146 -30286
rect -84 -31555 84 -31521
rect -84 -31663 84 -31629
rect -146 -32898 -112 -31722
rect 112 -32898 146 -31722
rect -84 -32991 84 -32957
rect -84 -33099 84 -33065
rect -146 -34334 -112 -33158
rect 112 -34334 146 -33158
rect -84 -34427 84 -34393
rect -84 -34535 84 -34501
rect -146 -35770 -112 -34594
rect 112 -35770 146 -34594
rect -84 -35863 84 -35829
rect -84 -35971 84 -35937
rect -146 -37206 -112 -36030
rect 112 -37206 146 -36030
rect -84 -37299 84 -37265
rect -84 -37407 84 -37373
rect -146 -38642 -112 -37466
rect 112 -38642 146 -37466
rect -84 -38735 84 -38701
rect -84 -38843 84 -38809
rect -146 -40078 -112 -38902
rect 112 -40078 146 -38902
rect -84 -40171 84 -40137
rect -84 -40279 84 -40245
rect -146 -41514 -112 -40338
rect 112 -41514 146 -40338
rect -84 -41607 84 -41573
rect -84 -41715 84 -41681
rect -146 -42950 -112 -41774
rect 112 -42950 146 -41774
rect -84 -43043 84 -43009
rect -84 -43151 84 -43117
rect -146 -44386 -112 -43210
rect 112 -44386 146 -43210
rect -84 -44479 84 -44445
rect -84 -44587 84 -44553
rect -146 -45822 -112 -44646
rect 112 -45822 146 -44646
rect -84 -45915 84 -45881
rect -84 -46023 84 -45989
rect -146 -47258 -112 -46082
rect 112 -47258 146 -46082
rect -84 -47351 84 -47317
rect -84 -47459 84 -47425
rect -146 -48694 -112 -47518
rect 112 -48694 146 -47518
rect -84 -48787 84 -48753
rect -84 -48895 84 -48861
rect -146 -50130 -112 -48954
rect 112 -50130 146 -48954
rect -84 -50223 84 -50189
rect -84 -50331 84 -50297
rect -146 -51566 -112 -50390
rect 112 -51566 146 -50390
rect -84 -51659 84 -51625
rect -84 -51767 84 -51733
rect -146 -53002 -112 -51826
rect 112 -53002 146 -51826
rect -84 -53095 84 -53061
rect -84 -53203 84 -53169
rect -146 -54438 -112 -53262
rect 112 -54438 146 -53262
rect -84 -54531 84 -54497
rect -84 -54639 84 -54605
rect -146 -55874 -112 -54698
rect 112 -55874 146 -54698
rect -84 -55967 84 -55933
rect -84 -56075 84 -56041
rect -146 -57310 -112 -56134
rect 112 -57310 146 -56134
rect -84 -57403 84 -57369
rect -84 -57511 84 -57477
rect -146 -58746 -112 -57570
rect 112 -58746 146 -57570
rect -84 -58839 84 -58805
rect -84 -58947 84 -58913
rect -146 -60182 -112 -59006
rect 112 -60182 146 -59006
rect -84 -60275 84 -60241
rect -84 -60383 84 -60349
rect -146 -61618 -112 -60442
rect 112 -61618 146 -60442
rect -84 -61711 84 -61677
rect -84 -61819 84 -61785
rect -146 -63054 -112 -61878
rect 112 -63054 146 -61878
rect -84 -63147 84 -63113
rect -84 -63255 84 -63221
rect -146 -64490 -112 -63314
rect 112 -64490 146 -63314
rect -84 -64583 84 -64549
rect -84 -64691 84 -64657
rect -146 -65926 -112 -64750
rect 112 -65926 146 -64750
rect -84 -66019 84 -65985
rect -84 -66127 84 -66093
rect -146 -67362 -112 -66186
rect 112 -67362 146 -66186
rect -84 -67455 84 -67421
rect -84 -67563 84 -67529
rect -146 -68798 -112 -67622
rect 112 -68798 146 -67622
rect -84 -68891 84 -68857
rect -84 -68999 84 -68965
rect -146 -70234 -112 -69058
rect 112 -70234 146 -69058
rect -84 -70327 84 -70293
rect -84 -70435 84 -70401
rect -146 -71670 -112 -70494
rect 112 -71670 146 -70494
rect -84 -71763 84 -71729
rect -84 -71871 84 -71837
rect -146 -73106 -112 -71930
rect 112 -73106 146 -71930
rect -84 -73199 84 -73165
rect -84 -73307 84 -73273
rect -146 -74542 -112 -73366
rect 112 -74542 146 -73366
rect -84 -74635 84 -74601
rect -84 -74743 84 -74709
rect -146 -75978 -112 -74802
rect 112 -75978 146 -74802
rect -84 -76071 84 -76037
rect -84 -76179 84 -76145
rect -146 -77414 -112 -76238
rect 112 -77414 146 -76238
rect -84 -77507 84 -77473
rect -84 -77615 84 -77581
rect -146 -78850 -112 -77674
rect 112 -78850 146 -77674
rect -84 -78943 84 -78909
rect -84 -79051 84 -79017
rect -146 -80286 -112 -79110
rect 112 -80286 146 -79110
rect -84 -80379 84 -80345
rect -84 -80487 84 -80453
rect -146 -81722 -112 -80546
rect 112 -81722 146 -80546
rect -84 -81815 84 -81781
rect -84 -81923 84 -81889
rect -146 -83158 -112 -81982
rect 112 -83158 146 -81982
rect -84 -83251 84 -83217
rect -84 -83359 84 -83325
rect -146 -84594 -112 -83418
rect 112 -84594 146 -83418
rect -84 -84687 84 -84653
rect -84 -84795 84 -84761
rect -146 -86030 -112 -84854
rect 112 -86030 146 -84854
rect -84 -86123 84 -86089
rect -84 -86231 84 -86197
rect -146 -87466 -112 -86290
rect 112 -87466 146 -86290
rect -84 -87559 84 -87525
rect -84 -87667 84 -87633
rect -146 -88902 -112 -87726
rect 112 -88902 146 -87726
rect -84 -88995 84 -88961
rect -84 -89103 84 -89069
rect -146 -90338 -112 -89162
rect 112 -90338 146 -89162
rect -84 -90431 84 -90397
rect -84 -90539 84 -90505
rect -146 -91774 -112 -90598
rect 112 -91774 146 -90598
rect -84 -91867 84 -91833
rect -84 -91975 84 -91941
rect -146 -93210 -112 -92034
rect 112 -93210 146 -92034
rect -84 -93303 84 -93269
rect -84 -93411 84 -93377
rect -146 -94646 -112 -93470
rect 112 -94646 146 -93470
rect -84 -94739 84 -94705
rect -84 -94847 84 -94813
rect -146 -96082 -112 -94906
rect 112 -96082 146 -94906
rect -84 -96175 84 -96141
rect -84 -96283 84 -96249
rect -146 -97518 -112 -96342
rect 112 -97518 146 -96342
rect -84 -97611 84 -97577
rect -84 -97719 84 -97685
rect -146 -98954 -112 -97778
rect 112 -98954 146 -97778
rect -84 -99047 84 -99013
rect -84 -99155 84 -99121
rect -146 -100390 -112 -99214
rect 112 -100390 146 -99214
rect -84 -100483 84 -100449
rect -84 -100591 84 -100557
rect -146 -101826 -112 -100650
rect 112 -101826 146 -100650
rect -84 -101919 84 -101885
rect -84 -102027 84 -101993
rect -146 -103262 -112 -102086
rect 112 -103262 146 -102086
rect -84 -103355 84 -103321
rect -84 -103463 84 -103429
rect -146 -104698 -112 -103522
rect 112 -104698 146 -103522
rect -84 -104791 84 -104757
rect -84 -104899 84 -104865
rect -146 -106134 -112 -104958
rect 112 -106134 146 -104958
rect -84 -106227 84 -106193
rect -84 -106335 84 -106301
rect -146 -107570 -112 -106394
rect 112 -107570 146 -106394
rect -84 -107663 84 -107629
rect -84 -107771 84 -107737
rect -146 -109006 -112 -107830
rect 112 -109006 146 -107830
rect -84 -109099 84 -109065
rect -84 -109207 84 -109173
rect -146 -110442 -112 -109266
rect 112 -110442 146 -109266
rect -84 -110535 84 -110501
rect -84 -110643 84 -110609
rect -146 -111878 -112 -110702
rect 112 -111878 146 -110702
rect -84 -111971 84 -111937
rect -84 -112079 84 -112045
rect -146 -113314 -112 -112138
rect 112 -113314 146 -112138
rect -84 -113407 84 -113373
rect -84 -113515 84 -113481
rect -146 -114750 -112 -113574
rect 112 -114750 146 -113574
rect -84 -114843 84 -114809
rect -84 -114951 84 -114917
rect -146 -116186 -112 -115010
rect 112 -116186 146 -115010
rect -84 -116279 84 -116245
rect -84 -116387 84 -116353
rect -146 -117622 -112 -116446
rect 112 -117622 146 -116446
rect -84 -117715 84 -117681
rect -84 -117823 84 -117789
rect -146 -119058 -112 -117882
rect 112 -119058 146 -117882
rect -84 -119151 84 -119117
rect -84 -119259 84 -119225
rect -146 -120494 -112 -119318
rect 112 -120494 146 -119318
rect -84 -120587 84 -120553
rect -84 -120695 84 -120661
rect -146 -121930 -112 -120754
rect 112 -121930 146 -120754
rect -84 -122023 84 -121989
rect -84 -122131 84 -122097
rect -146 -123366 -112 -122190
rect 112 -123366 146 -122190
rect -84 -123459 84 -123425
rect -84 -123567 84 -123533
rect -146 -124802 -112 -123626
rect 112 -124802 146 -123626
rect -84 -124895 84 -124861
rect -84 -125003 84 -124969
rect -146 -126238 -112 -125062
rect 112 -126238 146 -125062
rect -84 -126331 84 -126297
rect -84 -126439 84 -126405
rect -146 -127674 -112 -126498
rect 112 -127674 146 -126498
rect -84 -127767 84 -127733
rect -84 -127875 84 -127841
rect -146 -129110 -112 -127934
rect 112 -129110 146 -127934
rect -84 -129203 84 -129169
rect -84 -129311 84 -129277
rect -146 -130546 -112 -129370
rect 112 -130546 146 -129370
rect -84 -130639 84 -130605
rect -84 -130747 84 -130713
rect -146 -131982 -112 -130806
rect 112 -131982 146 -130806
rect -84 -132075 84 -132041
rect -84 -132183 84 -132149
rect -146 -133418 -112 -132242
rect 112 -133418 146 -132242
rect -84 -133511 84 -133477
rect -84 -133619 84 -133585
rect -146 -134854 -112 -133678
rect 112 -134854 146 -133678
rect -84 -134947 84 -134913
rect -84 -135055 84 -135021
rect -146 -136290 -112 -135114
rect 112 -136290 146 -135114
rect -84 -136383 84 -136349
rect -84 -136491 84 -136457
rect -146 -137726 -112 -136550
rect 112 -137726 146 -136550
rect -84 -137819 84 -137785
rect -84 -137927 84 -137893
rect -146 -139162 -112 -137986
rect 112 -139162 146 -137986
rect -84 -139255 84 -139221
rect -84 -139363 84 -139329
rect -146 -140598 -112 -139422
rect 112 -140598 146 -139422
rect -84 -140691 84 -140657
rect -84 -140799 84 -140765
rect -146 -142034 -112 -140858
rect 112 -142034 146 -140858
rect -84 -142127 84 -142093
rect -84 -142235 84 -142201
rect -146 -143470 -112 -142294
rect 112 -143470 146 -142294
rect -84 -143563 84 -143529
rect -84 -143671 84 -143637
rect -146 -144906 -112 -143730
rect 112 -144906 146 -143730
rect -84 -144999 84 -144965
rect -84 -145107 84 -145073
rect -146 -146342 -112 -145166
rect 112 -146342 146 -145166
rect -84 -146435 84 -146401
rect -84 -146543 84 -146509
rect -146 -147778 -112 -146602
rect 112 -147778 146 -146602
rect -84 -147871 84 -147837
rect -84 -147979 84 -147945
rect -146 -149214 -112 -148038
rect 112 -149214 146 -148038
rect -84 -149307 84 -149273
rect -84 -149415 84 -149381
rect -146 -150650 -112 -149474
rect 112 -150650 146 -149474
rect -84 -150743 84 -150709
rect -84 -150851 84 -150817
rect -146 -152086 -112 -150910
rect 112 -152086 146 -150910
rect -84 -152179 84 -152145
rect -84 -152287 84 -152253
rect -146 -153522 -112 -152346
rect 112 -153522 146 -152346
rect -84 -153615 84 -153581
rect -84 -153723 84 -153689
rect -146 -154958 -112 -153782
rect 112 -154958 146 -153782
rect -84 -155051 84 -155017
rect -84 -155159 84 -155125
rect -146 -156394 -112 -155218
rect 112 -156394 146 -155218
rect -84 -156487 84 -156453
rect -84 -156595 84 -156561
rect -146 -157830 -112 -156654
rect 112 -157830 146 -156654
rect -84 -157923 84 -157889
rect -84 -158031 84 -157997
rect -146 -159266 -112 -158090
rect 112 -159266 146 -158090
rect -84 -159359 84 -159325
rect -84 -159467 84 -159433
rect -146 -160702 -112 -159526
rect 112 -160702 146 -159526
rect -84 -160795 84 -160761
rect -84 -160903 84 -160869
rect -146 -162138 -112 -160962
rect 112 -162138 146 -160962
rect -84 -162231 84 -162197
rect -84 -162339 84 -162305
rect -146 -163574 -112 -162398
rect 112 -163574 146 -162398
rect -84 -163667 84 -163633
rect -84 -163775 84 -163741
rect -146 -165010 -112 -163834
rect 112 -165010 146 -163834
rect -84 -165103 84 -165069
rect -84 -165211 84 -165177
rect -146 -166446 -112 -165270
rect 112 -166446 146 -165270
rect -84 -166539 84 -166505
rect -84 -166647 84 -166613
rect -146 -167882 -112 -166706
rect 112 -167882 146 -166706
rect -84 -167975 84 -167941
rect -84 -168083 84 -168049
rect -146 -169318 -112 -168142
rect 112 -169318 146 -168142
rect -84 -169411 84 -169377
rect -84 -169519 84 -169485
rect -146 -170754 -112 -169578
rect 112 -170754 146 -169578
rect -84 -170847 84 -170813
rect -84 -170955 84 -170921
rect -146 -172190 -112 -171014
rect 112 -172190 146 -171014
rect -84 -172283 84 -172249
rect -84 -172391 84 -172357
rect -146 -173626 -112 -172450
rect 112 -173626 146 -172450
rect -84 -173719 84 -173685
rect -84 -173827 84 -173793
rect -146 -175062 -112 -173886
rect 112 -175062 146 -173886
rect -84 -175155 84 -175121
rect -84 -175263 84 -175229
rect -146 -176498 -112 -175322
rect 112 -176498 146 -175322
rect -84 -176591 84 -176557
rect -84 -176699 84 -176665
rect -146 -177934 -112 -176758
rect 112 -177934 146 -176758
rect -84 -178027 84 -177993
rect -84 -178135 84 -178101
rect -146 -179370 -112 -178194
rect 112 -179370 146 -178194
rect -84 -179463 84 -179429
rect -84 -179571 84 -179537
rect -146 -180806 -112 -179630
rect 112 -180806 146 -179630
rect -84 -180899 84 -180865
rect -84 -181007 84 -180973
rect -146 -182242 -112 -181066
rect 112 -182242 146 -181066
rect -84 -182335 84 -182301
rect -84 -182443 84 -182409
rect -146 -183678 -112 -182502
rect 112 -183678 146 -182502
rect -84 -183771 84 -183737
<< metal1 >>
rect -96 183771 96 183777
rect -96 183737 -84 183771
rect 84 183737 96 183771
rect -96 183731 96 183737
rect -152 183678 -106 183690
rect -152 182502 -146 183678
rect -112 182502 -106 183678
rect -152 182490 -106 182502
rect 106 183678 152 183690
rect 106 182502 112 183678
rect 146 182502 152 183678
rect 106 182490 152 182502
rect -96 182443 96 182449
rect -96 182409 -84 182443
rect 84 182409 96 182443
rect -96 182403 96 182409
rect -96 182335 96 182341
rect -96 182301 -84 182335
rect 84 182301 96 182335
rect -96 182295 96 182301
rect -152 182242 -106 182254
rect -152 181066 -146 182242
rect -112 181066 -106 182242
rect -152 181054 -106 181066
rect 106 182242 152 182254
rect 106 181066 112 182242
rect 146 181066 152 182242
rect 106 181054 152 181066
rect -96 181007 96 181013
rect -96 180973 -84 181007
rect 84 180973 96 181007
rect -96 180967 96 180973
rect -96 180899 96 180905
rect -96 180865 -84 180899
rect 84 180865 96 180899
rect -96 180859 96 180865
rect -152 180806 -106 180818
rect -152 179630 -146 180806
rect -112 179630 -106 180806
rect -152 179618 -106 179630
rect 106 180806 152 180818
rect 106 179630 112 180806
rect 146 179630 152 180806
rect 106 179618 152 179630
rect -96 179571 96 179577
rect -96 179537 -84 179571
rect 84 179537 96 179571
rect -96 179531 96 179537
rect -96 179463 96 179469
rect -96 179429 -84 179463
rect 84 179429 96 179463
rect -96 179423 96 179429
rect -152 179370 -106 179382
rect -152 178194 -146 179370
rect -112 178194 -106 179370
rect -152 178182 -106 178194
rect 106 179370 152 179382
rect 106 178194 112 179370
rect 146 178194 152 179370
rect 106 178182 152 178194
rect -96 178135 96 178141
rect -96 178101 -84 178135
rect 84 178101 96 178135
rect -96 178095 96 178101
rect -96 178027 96 178033
rect -96 177993 -84 178027
rect 84 177993 96 178027
rect -96 177987 96 177993
rect -152 177934 -106 177946
rect -152 176758 -146 177934
rect -112 176758 -106 177934
rect -152 176746 -106 176758
rect 106 177934 152 177946
rect 106 176758 112 177934
rect 146 176758 152 177934
rect 106 176746 152 176758
rect -96 176699 96 176705
rect -96 176665 -84 176699
rect 84 176665 96 176699
rect -96 176659 96 176665
rect -96 176591 96 176597
rect -96 176557 -84 176591
rect 84 176557 96 176591
rect -96 176551 96 176557
rect -152 176498 -106 176510
rect -152 175322 -146 176498
rect -112 175322 -106 176498
rect -152 175310 -106 175322
rect 106 176498 152 176510
rect 106 175322 112 176498
rect 146 175322 152 176498
rect 106 175310 152 175322
rect -96 175263 96 175269
rect -96 175229 -84 175263
rect 84 175229 96 175263
rect -96 175223 96 175229
rect -96 175155 96 175161
rect -96 175121 -84 175155
rect 84 175121 96 175155
rect -96 175115 96 175121
rect -152 175062 -106 175074
rect -152 173886 -146 175062
rect -112 173886 -106 175062
rect -152 173874 -106 173886
rect 106 175062 152 175074
rect 106 173886 112 175062
rect 146 173886 152 175062
rect 106 173874 152 173886
rect -96 173827 96 173833
rect -96 173793 -84 173827
rect 84 173793 96 173827
rect -96 173787 96 173793
rect -96 173719 96 173725
rect -96 173685 -84 173719
rect 84 173685 96 173719
rect -96 173679 96 173685
rect -152 173626 -106 173638
rect -152 172450 -146 173626
rect -112 172450 -106 173626
rect -152 172438 -106 172450
rect 106 173626 152 173638
rect 106 172450 112 173626
rect 146 172450 152 173626
rect 106 172438 152 172450
rect -96 172391 96 172397
rect -96 172357 -84 172391
rect 84 172357 96 172391
rect -96 172351 96 172357
rect -96 172283 96 172289
rect -96 172249 -84 172283
rect 84 172249 96 172283
rect -96 172243 96 172249
rect -152 172190 -106 172202
rect -152 171014 -146 172190
rect -112 171014 -106 172190
rect -152 171002 -106 171014
rect 106 172190 152 172202
rect 106 171014 112 172190
rect 146 171014 152 172190
rect 106 171002 152 171014
rect -96 170955 96 170961
rect -96 170921 -84 170955
rect 84 170921 96 170955
rect -96 170915 96 170921
rect -96 170847 96 170853
rect -96 170813 -84 170847
rect 84 170813 96 170847
rect -96 170807 96 170813
rect -152 170754 -106 170766
rect -152 169578 -146 170754
rect -112 169578 -106 170754
rect -152 169566 -106 169578
rect 106 170754 152 170766
rect 106 169578 112 170754
rect 146 169578 152 170754
rect 106 169566 152 169578
rect -96 169519 96 169525
rect -96 169485 -84 169519
rect 84 169485 96 169519
rect -96 169479 96 169485
rect -96 169411 96 169417
rect -96 169377 -84 169411
rect 84 169377 96 169411
rect -96 169371 96 169377
rect -152 169318 -106 169330
rect -152 168142 -146 169318
rect -112 168142 -106 169318
rect -152 168130 -106 168142
rect 106 169318 152 169330
rect 106 168142 112 169318
rect 146 168142 152 169318
rect 106 168130 152 168142
rect -96 168083 96 168089
rect -96 168049 -84 168083
rect 84 168049 96 168083
rect -96 168043 96 168049
rect -96 167975 96 167981
rect -96 167941 -84 167975
rect 84 167941 96 167975
rect -96 167935 96 167941
rect -152 167882 -106 167894
rect -152 166706 -146 167882
rect -112 166706 -106 167882
rect -152 166694 -106 166706
rect 106 167882 152 167894
rect 106 166706 112 167882
rect 146 166706 152 167882
rect 106 166694 152 166706
rect -96 166647 96 166653
rect -96 166613 -84 166647
rect 84 166613 96 166647
rect -96 166607 96 166613
rect -96 166539 96 166545
rect -96 166505 -84 166539
rect 84 166505 96 166539
rect -96 166499 96 166505
rect -152 166446 -106 166458
rect -152 165270 -146 166446
rect -112 165270 -106 166446
rect -152 165258 -106 165270
rect 106 166446 152 166458
rect 106 165270 112 166446
rect 146 165270 152 166446
rect 106 165258 152 165270
rect -96 165211 96 165217
rect -96 165177 -84 165211
rect 84 165177 96 165211
rect -96 165171 96 165177
rect -96 165103 96 165109
rect -96 165069 -84 165103
rect 84 165069 96 165103
rect -96 165063 96 165069
rect -152 165010 -106 165022
rect -152 163834 -146 165010
rect -112 163834 -106 165010
rect -152 163822 -106 163834
rect 106 165010 152 165022
rect 106 163834 112 165010
rect 146 163834 152 165010
rect 106 163822 152 163834
rect -96 163775 96 163781
rect -96 163741 -84 163775
rect 84 163741 96 163775
rect -96 163735 96 163741
rect -96 163667 96 163673
rect -96 163633 -84 163667
rect 84 163633 96 163667
rect -96 163627 96 163633
rect -152 163574 -106 163586
rect -152 162398 -146 163574
rect -112 162398 -106 163574
rect -152 162386 -106 162398
rect 106 163574 152 163586
rect 106 162398 112 163574
rect 146 162398 152 163574
rect 106 162386 152 162398
rect -96 162339 96 162345
rect -96 162305 -84 162339
rect 84 162305 96 162339
rect -96 162299 96 162305
rect -96 162231 96 162237
rect -96 162197 -84 162231
rect 84 162197 96 162231
rect -96 162191 96 162197
rect -152 162138 -106 162150
rect -152 160962 -146 162138
rect -112 160962 -106 162138
rect -152 160950 -106 160962
rect 106 162138 152 162150
rect 106 160962 112 162138
rect 146 160962 152 162138
rect 106 160950 152 160962
rect -96 160903 96 160909
rect -96 160869 -84 160903
rect 84 160869 96 160903
rect -96 160863 96 160869
rect -96 160795 96 160801
rect -96 160761 -84 160795
rect 84 160761 96 160795
rect -96 160755 96 160761
rect -152 160702 -106 160714
rect -152 159526 -146 160702
rect -112 159526 -106 160702
rect -152 159514 -106 159526
rect 106 160702 152 160714
rect 106 159526 112 160702
rect 146 159526 152 160702
rect 106 159514 152 159526
rect -96 159467 96 159473
rect -96 159433 -84 159467
rect 84 159433 96 159467
rect -96 159427 96 159433
rect -96 159359 96 159365
rect -96 159325 -84 159359
rect 84 159325 96 159359
rect -96 159319 96 159325
rect -152 159266 -106 159278
rect -152 158090 -146 159266
rect -112 158090 -106 159266
rect -152 158078 -106 158090
rect 106 159266 152 159278
rect 106 158090 112 159266
rect 146 158090 152 159266
rect 106 158078 152 158090
rect -96 158031 96 158037
rect -96 157997 -84 158031
rect 84 157997 96 158031
rect -96 157991 96 157997
rect -96 157923 96 157929
rect -96 157889 -84 157923
rect 84 157889 96 157923
rect -96 157883 96 157889
rect -152 157830 -106 157842
rect -152 156654 -146 157830
rect -112 156654 -106 157830
rect -152 156642 -106 156654
rect 106 157830 152 157842
rect 106 156654 112 157830
rect 146 156654 152 157830
rect 106 156642 152 156654
rect -96 156595 96 156601
rect -96 156561 -84 156595
rect 84 156561 96 156595
rect -96 156555 96 156561
rect -96 156487 96 156493
rect -96 156453 -84 156487
rect 84 156453 96 156487
rect -96 156447 96 156453
rect -152 156394 -106 156406
rect -152 155218 -146 156394
rect -112 155218 -106 156394
rect -152 155206 -106 155218
rect 106 156394 152 156406
rect 106 155218 112 156394
rect 146 155218 152 156394
rect 106 155206 152 155218
rect -96 155159 96 155165
rect -96 155125 -84 155159
rect 84 155125 96 155159
rect -96 155119 96 155125
rect -96 155051 96 155057
rect -96 155017 -84 155051
rect 84 155017 96 155051
rect -96 155011 96 155017
rect -152 154958 -106 154970
rect -152 153782 -146 154958
rect -112 153782 -106 154958
rect -152 153770 -106 153782
rect 106 154958 152 154970
rect 106 153782 112 154958
rect 146 153782 152 154958
rect 106 153770 152 153782
rect -96 153723 96 153729
rect -96 153689 -84 153723
rect 84 153689 96 153723
rect -96 153683 96 153689
rect -96 153615 96 153621
rect -96 153581 -84 153615
rect 84 153581 96 153615
rect -96 153575 96 153581
rect -152 153522 -106 153534
rect -152 152346 -146 153522
rect -112 152346 -106 153522
rect -152 152334 -106 152346
rect 106 153522 152 153534
rect 106 152346 112 153522
rect 146 152346 152 153522
rect 106 152334 152 152346
rect -96 152287 96 152293
rect -96 152253 -84 152287
rect 84 152253 96 152287
rect -96 152247 96 152253
rect -96 152179 96 152185
rect -96 152145 -84 152179
rect 84 152145 96 152179
rect -96 152139 96 152145
rect -152 152086 -106 152098
rect -152 150910 -146 152086
rect -112 150910 -106 152086
rect -152 150898 -106 150910
rect 106 152086 152 152098
rect 106 150910 112 152086
rect 146 150910 152 152086
rect 106 150898 152 150910
rect -96 150851 96 150857
rect -96 150817 -84 150851
rect 84 150817 96 150851
rect -96 150811 96 150817
rect -96 150743 96 150749
rect -96 150709 -84 150743
rect 84 150709 96 150743
rect -96 150703 96 150709
rect -152 150650 -106 150662
rect -152 149474 -146 150650
rect -112 149474 -106 150650
rect -152 149462 -106 149474
rect 106 150650 152 150662
rect 106 149474 112 150650
rect 146 149474 152 150650
rect 106 149462 152 149474
rect -96 149415 96 149421
rect -96 149381 -84 149415
rect 84 149381 96 149415
rect -96 149375 96 149381
rect -96 149307 96 149313
rect -96 149273 -84 149307
rect 84 149273 96 149307
rect -96 149267 96 149273
rect -152 149214 -106 149226
rect -152 148038 -146 149214
rect -112 148038 -106 149214
rect -152 148026 -106 148038
rect 106 149214 152 149226
rect 106 148038 112 149214
rect 146 148038 152 149214
rect 106 148026 152 148038
rect -96 147979 96 147985
rect -96 147945 -84 147979
rect 84 147945 96 147979
rect -96 147939 96 147945
rect -96 147871 96 147877
rect -96 147837 -84 147871
rect 84 147837 96 147871
rect -96 147831 96 147837
rect -152 147778 -106 147790
rect -152 146602 -146 147778
rect -112 146602 -106 147778
rect -152 146590 -106 146602
rect 106 147778 152 147790
rect 106 146602 112 147778
rect 146 146602 152 147778
rect 106 146590 152 146602
rect -96 146543 96 146549
rect -96 146509 -84 146543
rect 84 146509 96 146543
rect -96 146503 96 146509
rect -96 146435 96 146441
rect -96 146401 -84 146435
rect 84 146401 96 146435
rect -96 146395 96 146401
rect -152 146342 -106 146354
rect -152 145166 -146 146342
rect -112 145166 -106 146342
rect -152 145154 -106 145166
rect 106 146342 152 146354
rect 106 145166 112 146342
rect 146 145166 152 146342
rect 106 145154 152 145166
rect -96 145107 96 145113
rect -96 145073 -84 145107
rect 84 145073 96 145107
rect -96 145067 96 145073
rect -96 144999 96 145005
rect -96 144965 -84 144999
rect 84 144965 96 144999
rect -96 144959 96 144965
rect -152 144906 -106 144918
rect -152 143730 -146 144906
rect -112 143730 -106 144906
rect -152 143718 -106 143730
rect 106 144906 152 144918
rect 106 143730 112 144906
rect 146 143730 152 144906
rect 106 143718 152 143730
rect -96 143671 96 143677
rect -96 143637 -84 143671
rect 84 143637 96 143671
rect -96 143631 96 143637
rect -96 143563 96 143569
rect -96 143529 -84 143563
rect 84 143529 96 143563
rect -96 143523 96 143529
rect -152 143470 -106 143482
rect -152 142294 -146 143470
rect -112 142294 -106 143470
rect -152 142282 -106 142294
rect 106 143470 152 143482
rect 106 142294 112 143470
rect 146 142294 152 143470
rect 106 142282 152 142294
rect -96 142235 96 142241
rect -96 142201 -84 142235
rect 84 142201 96 142235
rect -96 142195 96 142201
rect -96 142127 96 142133
rect -96 142093 -84 142127
rect 84 142093 96 142127
rect -96 142087 96 142093
rect -152 142034 -106 142046
rect -152 140858 -146 142034
rect -112 140858 -106 142034
rect -152 140846 -106 140858
rect 106 142034 152 142046
rect 106 140858 112 142034
rect 146 140858 152 142034
rect 106 140846 152 140858
rect -96 140799 96 140805
rect -96 140765 -84 140799
rect 84 140765 96 140799
rect -96 140759 96 140765
rect -96 140691 96 140697
rect -96 140657 -84 140691
rect 84 140657 96 140691
rect -96 140651 96 140657
rect -152 140598 -106 140610
rect -152 139422 -146 140598
rect -112 139422 -106 140598
rect -152 139410 -106 139422
rect 106 140598 152 140610
rect 106 139422 112 140598
rect 146 139422 152 140598
rect 106 139410 152 139422
rect -96 139363 96 139369
rect -96 139329 -84 139363
rect 84 139329 96 139363
rect -96 139323 96 139329
rect -96 139255 96 139261
rect -96 139221 -84 139255
rect 84 139221 96 139255
rect -96 139215 96 139221
rect -152 139162 -106 139174
rect -152 137986 -146 139162
rect -112 137986 -106 139162
rect -152 137974 -106 137986
rect 106 139162 152 139174
rect 106 137986 112 139162
rect 146 137986 152 139162
rect 106 137974 152 137986
rect -96 137927 96 137933
rect -96 137893 -84 137927
rect 84 137893 96 137927
rect -96 137887 96 137893
rect -96 137819 96 137825
rect -96 137785 -84 137819
rect 84 137785 96 137819
rect -96 137779 96 137785
rect -152 137726 -106 137738
rect -152 136550 -146 137726
rect -112 136550 -106 137726
rect -152 136538 -106 136550
rect 106 137726 152 137738
rect 106 136550 112 137726
rect 146 136550 152 137726
rect 106 136538 152 136550
rect -96 136491 96 136497
rect -96 136457 -84 136491
rect 84 136457 96 136491
rect -96 136451 96 136457
rect -96 136383 96 136389
rect -96 136349 -84 136383
rect 84 136349 96 136383
rect -96 136343 96 136349
rect -152 136290 -106 136302
rect -152 135114 -146 136290
rect -112 135114 -106 136290
rect -152 135102 -106 135114
rect 106 136290 152 136302
rect 106 135114 112 136290
rect 146 135114 152 136290
rect 106 135102 152 135114
rect -96 135055 96 135061
rect -96 135021 -84 135055
rect 84 135021 96 135055
rect -96 135015 96 135021
rect -96 134947 96 134953
rect -96 134913 -84 134947
rect 84 134913 96 134947
rect -96 134907 96 134913
rect -152 134854 -106 134866
rect -152 133678 -146 134854
rect -112 133678 -106 134854
rect -152 133666 -106 133678
rect 106 134854 152 134866
rect 106 133678 112 134854
rect 146 133678 152 134854
rect 106 133666 152 133678
rect -96 133619 96 133625
rect -96 133585 -84 133619
rect 84 133585 96 133619
rect -96 133579 96 133585
rect -96 133511 96 133517
rect -96 133477 -84 133511
rect 84 133477 96 133511
rect -96 133471 96 133477
rect -152 133418 -106 133430
rect -152 132242 -146 133418
rect -112 132242 -106 133418
rect -152 132230 -106 132242
rect 106 133418 152 133430
rect 106 132242 112 133418
rect 146 132242 152 133418
rect 106 132230 152 132242
rect -96 132183 96 132189
rect -96 132149 -84 132183
rect 84 132149 96 132183
rect -96 132143 96 132149
rect -96 132075 96 132081
rect -96 132041 -84 132075
rect 84 132041 96 132075
rect -96 132035 96 132041
rect -152 131982 -106 131994
rect -152 130806 -146 131982
rect -112 130806 -106 131982
rect -152 130794 -106 130806
rect 106 131982 152 131994
rect 106 130806 112 131982
rect 146 130806 152 131982
rect 106 130794 152 130806
rect -96 130747 96 130753
rect -96 130713 -84 130747
rect 84 130713 96 130747
rect -96 130707 96 130713
rect -96 130639 96 130645
rect -96 130605 -84 130639
rect 84 130605 96 130639
rect -96 130599 96 130605
rect -152 130546 -106 130558
rect -152 129370 -146 130546
rect -112 129370 -106 130546
rect -152 129358 -106 129370
rect 106 130546 152 130558
rect 106 129370 112 130546
rect 146 129370 152 130546
rect 106 129358 152 129370
rect -96 129311 96 129317
rect -96 129277 -84 129311
rect 84 129277 96 129311
rect -96 129271 96 129277
rect -96 129203 96 129209
rect -96 129169 -84 129203
rect 84 129169 96 129203
rect -96 129163 96 129169
rect -152 129110 -106 129122
rect -152 127934 -146 129110
rect -112 127934 -106 129110
rect -152 127922 -106 127934
rect 106 129110 152 129122
rect 106 127934 112 129110
rect 146 127934 152 129110
rect 106 127922 152 127934
rect -96 127875 96 127881
rect -96 127841 -84 127875
rect 84 127841 96 127875
rect -96 127835 96 127841
rect -96 127767 96 127773
rect -96 127733 -84 127767
rect 84 127733 96 127767
rect -96 127727 96 127733
rect -152 127674 -106 127686
rect -152 126498 -146 127674
rect -112 126498 -106 127674
rect -152 126486 -106 126498
rect 106 127674 152 127686
rect 106 126498 112 127674
rect 146 126498 152 127674
rect 106 126486 152 126498
rect -96 126439 96 126445
rect -96 126405 -84 126439
rect 84 126405 96 126439
rect -96 126399 96 126405
rect -96 126331 96 126337
rect -96 126297 -84 126331
rect 84 126297 96 126331
rect -96 126291 96 126297
rect -152 126238 -106 126250
rect -152 125062 -146 126238
rect -112 125062 -106 126238
rect -152 125050 -106 125062
rect 106 126238 152 126250
rect 106 125062 112 126238
rect 146 125062 152 126238
rect 106 125050 152 125062
rect -96 125003 96 125009
rect -96 124969 -84 125003
rect 84 124969 96 125003
rect -96 124963 96 124969
rect -96 124895 96 124901
rect -96 124861 -84 124895
rect 84 124861 96 124895
rect -96 124855 96 124861
rect -152 124802 -106 124814
rect -152 123626 -146 124802
rect -112 123626 -106 124802
rect -152 123614 -106 123626
rect 106 124802 152 124814
rect 106 123626 112 124802
rect 146 123626 152 124802
rect 106 123614 152 123626
rect -96 123567 96 123573
rect -96 123533 -84 123567
rect 84 123533 96 123567
rect -96 123527 96 123533
rect -96 123459 96 123465
rect -96 123425 -84 123459
rect 84 123425 96 123459
rect -96 123419 96 123425
rect -152 123366 -106 123378
rect -152 122190 -146 123366
rect -112 122190 -106 123366
rect -152 122178 -106 122190
rect 106 123366 152 123378
rect 106 122190 112 123366
rect 146 122190 152 123366
rect 106 122178 152 122190
rect -96 122131 96 122137
rect -96 122097 -84 122131
rect 84 122097 96 122131
rect -96 122091 96 122097
rect -96 122023 96 122029
rect -96 121989 -84 122023
rect 84 121989 96 122023
rect -96 121983 96 121989
rect -152 121930 -106 121942
rect -152 120754 -146 121930
rect -112 120754 -106 121930
rect -152 120742 -106 120754
rect 106 121930 152 121942
rect 106 120754 112 121930
rect 146 120754 152 121930
rect 106 120742 152 120754
rect -96 120695 96 120701
rect -96 120661 -84 120695
rect 84 120661 96 120695
rect -96 120655 96 120661
rect -96 120587 96 120593
rect -96 120553 -84 120587
rect 84 120553 96 120587
rect -96 120547 96 120553
rect -152 120494 -106 120506
rect -152 119318 -146 120494
rect -112 119318 -106 120494
rect -152 119306 -106 119318
rect 106 120494 152 120506
rect 106 119318 112 120494
rect 146 119318 152 120494
rect 106 119306 152 119318
rect -96 119259 96 119265
rect -96 119225 -84 119259
rect 84 119225 96 119259
rect -96 119219 96 119225
rect -96 119151 96 119157
rect -96 119117 -84 119151
rect 84 119117 96 119151
rect -96 119111 96 119117
rect -152 119058 -106 119070
rect -152 117882 -146 119058
rect -112 117882 -106 119058
rect -152 117870 -106 117882
rect 106 119058 152 119070
rect 106 117882 112 119058
rect 146 117882 152 119058
rect 106 117870 152 117882
rect -96 117823 96 117829
rect -96 117789 -84 117823
rect 84 117789 96 117823
rect -96 117783 96 117789
rect -96 117715 96 117721
rect -96 117681 -84 117715
rect 84 117681 96 117715
rect -96 117675 96 117681
rect -152 117622 -106 117634
rect -152 116446 -146 117622
rect -112 116446 -106 117622
rect -152 116434 -106 116446
rect 106 117622 152 117634
rect 106 116446 112 117622
rect 146 116446 152 117622
rect 106 116434 152 116446
rect -96 116387 96 116393
rect -96 116353 -84 116387
rect 84 116353 96 116387
rect -96 116347 96 116353
rect -96 116279 96 116285
rect -96 116245 -84 116279
rect 84 116245 96 116279
rect -96 116239 96 116245
rect -152 116186 -106 116198
rect -152 115010 -146 116186
rect -112 115010 -106 116186
rect -152 114998 -106 115010
rect 106 116186 152 116198
rect 106 115010 112 116186
rect 146 115010 152 116186
rect 106 114998 152 115010
rect -96 114951 96 114957
rect -96 114917 -84 114951
rect 84 114917 96 114951
rect -96 114911 96 114917
rect -96 114843 96 114849
rect -96 114809 -84 114843
rect 84 114809 96 114843
rect -96 114803 96 114809
rect -152 114750 -106 114762
rect -152 113574 -146 114750
rect -112 113574 -106 114750
rect -152 113562 -106 113574
rect 106 114750 152 114762
rect 106 113574 112 114750
rect 146 113574 152 114750
rect 106 113562 152 113574
rect -96 113515 96 113521
rect -96 113481 -84 113515
rect 84 113481 96 113515
rect -96 113475 96 113481
rect -96 113407 96 113413
rect -96 113373 -84 113407
rect 84 113373 96 113407
rect -96 113367 96 113373
rect -152 113314 -106 113326
rect -152 112138 -146 113314
rect -112 112138 -106 113314
rect -152 112126 -106 112138
rect 106 113314 152 113326
rect 106 112138 112 113314
rect 146 112138 152 113314
rect 106 112126 152 112138
rect -96 112079 96 112085
rect -96 112045 -84 112079
rect 84 112045 96 112079
rect -96 112039 96 112045
rect -96 111971 96 111977
rect -96 111937 -84 111971
rect 84 111937 96 111971
rect -96 111931 96 111937
rect -152 111878 -106 111890
rect -152 110702 -146 111878
rect -112 110702 -106 111878
rect -152 110690 -106 110702
rect 106 111878 152 111890
rect 106 110702 112 111878
rect 146 110702 152 111878
rect 106 110690 152 110702
rect -96 110643 96 110649
rect -96 110609 -84 110643
rect 84 110609 96 110643
rect -96 110603 96 110609
rect -96 110535 96 110541
rect -96 110501 -84 110535
rect 84 110501 96 110535
rect -96 110495 96 110501
rect -152 110442 -106 110454
rect -152 109266 -146 110442
rect -112 109266 -106 110442
rect -152 109254 -106 109266
rect 106 110442 152 110454
rect 106 109266 112 110442
rect 146 109266 152 110442
rect 106 109254 152 109266
rect -96 109207 96 109213
rect -96 109173 -84 109207
rect 84 109173 96 109207
rect -96 109167 96 109173
rect -96 109099 96 109105
rect -96 109065 -84 109099
rect 84 109065 96 109099
rect -96 109059 96 109065
rect -152 109006 -106 109018
rect -152 107830 -146 109006
rect -112 107830 -106 109006
rect -152 107818 -106 107830
rect 106 109006 152 109018
rect 106 107830 112 109006
rect 146 107830 152 109006
rect 106 107818 152 107830
rect -96 107771 96 107777
rect -96 107737 -84 107771
rect 84 107737 96 107771
rect -96 107731 96 107737
rect -96 107663 96 107669
rect -96 107629 -84 107663
rect 84 107629 96 107663
rect -96 107623 96 107629
rect -152 107570 -106 107582
rect -152 106394 -146 107570
rect -112 106394 -106 107570
rect -152 106382 -106 106394
rect 106 107570 152 107582
rect 106 106394 112 107570
rect 146 106394 152 107570
rect 106 106382 152 106394
rect -96 106335 96 106341
rect -96 106301 -84 106335
rect 84 106301 96 106335
rect -96 106295 96 106301
rect -96 106227 96 106233
rect -96 106193 -84 106227
rect 84 106193 96 106227
rect -96 106187 96 106193
rect -152 106134 -106 106146
rect -152 104958 -146 106134
rect -112 104958 -106 106134
rect -152 104946 -106 104958
rect 106 106134 152 106146
rect 106 104958 112 106134
rect 146 104958 152 106134
rect 106 104946 152 104958
rect -96 104899 96 104905
rect -96 104865 -84 104899
rect 84 104865 96 104899
rect -96 104859 96 104865
rect -96 104791 96 104797
rect -96 104757 -84 104791
rect 84 104757 96 104791
rect -96 104751 96 104757
rect -152 104698 -106 104710
rect -152 103522 -146 104698
rect -112 103522 -106 104698
rect -152 103510 -106 103522
rect 106 104698 152 104710
rect 106 103522 112 104698
rect 146 103522 152 104698
rect 106 103510 152 103522
rect -96 103463 96 103469
rect -96 103429 -84 103463
rect 84 103429 96 103463
rect -96 103423 96 103429
rect -96 103355 96 103361
rect -96 103321 -84 103355
rect 84 103321 96 103355
rect -96 103315 96 103321
rect -152 103262 -106 103274
rect -152 102086 -146 103262
rect -112 102086 -106 103262
rect -152 102074 -106 102086
rect 106 103262 152 103274
rect 106 102086 112 103262
rect 146 102086 152 103262
rect 106 102074 152 102086
rect -96 102027 96 102033
rect -96 101993 -84 102027
rect 84 101993 96 102027
rect -96 101987 96 101993
rect -96 101919 96 101925
rect -96 101885 -84 101919
rect 84 101885 96 101919
rect -96 101879 96 101885
rect -152 101826 -106 101838
rect -152 100650 -146 101826
rect -112 100650 -106 101826
rect -152 100638 -106 100650
rect 106 101826 152 101838
rect 106 100650 112 101826
rect 146 100650 152 101826
rect 106 100638 152 100650
rect -96 100591 96 100597
rect -96 100557 -84 100591
rect 84 100557 96 100591
rect -96 100551 96 100557
rect -96 100483 96 100489
rect -96 100449 -84 100483
rect 84 100449 96 100483
rect -96 100443 96 100449
rect -152 100390 -106 100402
rect -152 99214 -146 100390
rect -112 99214 -106 100390
rect -152 99202 -106 99214
rect 106 100390 152 100402
rect 106 99214 112 100390
rect 146 99214 152 100390
rect 106 99202 152 99214
rect -96 99155 96 99161
rect -96 99121 -84 99155
rect 84 99121 96 99155
rect -96 99115 96 99121
rect -96 99047 96 99053
rect -96 99013 -84 99047
rect 84 99013 96 99047
rect -96 99007 96 99013
rect -152 98954 -106 98966
rect -152 97778 -146 98954
rect -112 97778 -106 98954
rect -152 97766 -106 97778
rect 106 98954 152 98966
rect 106 97778 112 98954
rect 146 97778 152 98954
rect 106 97766 152 97778
rect -96 97719 96 97725
rect -96 97685 -84 97719
rect 84 97685 96 97719
rect -96 97679 96 97685
rect -96 97611 96 97617
rect -96 97577 -84 97611
rect 84 97577 96 97611
rect -96 97571 96 97577
rect -152 97518 -106 97530
rect -152 96342 -146 97518
rect -112 96342 -106 97518
rect -152 96330 -106 96342
rect 106 97518 152 97530
rect 106 96342 112 97518
rect 146 96342 152 97518
rect 106 96330 152 96342
rect -96 96283 96 96289
rect -96 96249 -84 96283
rect 84 96249 96 96283
rect -96 96243 96 96249
rect -96 96175 96 96181
rect -96 96141 -84 96175
rect 84 96141 96 96175
rect -96 96135 96 96141
rect -152 96082 -106 96094
rect -152 94906 -146 96082
rect -112 94906 -106 96082
rect -152 94894 -106 94906
rect 106 96082 152 96094
rect 106 94906 112 96082
rect 146 94906 152 96082
rect 106 94894 152 94906
rect -96 94847 96 94853
rect -96 94813 -84 94847
rect 84 94813 96 94847
rect -96 94807 96 94813
rect -96 94739 96 94745
rect -96 94705 -84 94739
rect 84 94705 96 94739
rect -96 94699 96 94705
rect -152 94646 -106 94658
rect -152 93470 -146 94646
rect -112 93470 -106 94646
rect -152 93458 -106 93470
rect 106 94646 152 94658
rect 106 93470 112 94646
rect 146 93470 152 94646
rect 106 93458 152 93470
rect -96 93411 96 93417
rect -96 93377 -84 93411
rect 84 93377 96 93411
rect -96 93371 96 93377
rect -96 93303 96 93309
rect -96 93269 -84 93303
rect 84 93269 96 93303
rect -96 93263 96 93269
rect -152 93210 -106 93222
rect -152 92034 -146 93210
rect -112 92034 -106 93210
rect -152 92022 -106 92034
rect 106 93210 152 93222
rect 106 92034 112 93210
rect 146 92034 152 93210
rect 106 92022 152 92034
rect -96 91975 96 91981
rect -96 91941 -84 91975
rect 84 91941 96 91975
rect -96 91935 96 91941
rect -96 91867 96 91873
rect -96 91833 -84 91867
rect 84 91833 96 91867
rect -96 91827 96 91833
rect -152 91774 -106 91786
rect -152 90598 -146 91774
rect -112 90598 -106 91774
rect -152 90586 -106 90598
rect 106 91774 152 91786
rect 106 90598 112 91774
rect 146 90598 152 91774
rect 106 90586 152 90598
rect -96 90539 96 90545
rect -96 90505 -84 90539
rect 84 90505 96 90539
rect -96 90499 96 90505
rect -96 90431 96 90437
rect -96 90397 -84 90431
rect 84 90397 96 90431
rect -96 90391 96 90397
rect -152 90338 -106 90350
rect -152 89162 -146 90338
rect -112 89162 -106 90338
rect -152 89150 -106 89162
rect 106 90338 152 90350
rect 106 89162 112 90338
rect 146 89162 152 90338
rect 106 89150 152 89162
rect -96 89103 96 89109
rect -96 89069 -84 89103
rect 84 89069 96 89103
rect -96 89063 96 89069
rect -96 88995 96 89001
rect -96 88961 -84 88995
rect 84 88961 96 88995
rect -96 88955 96 88961
rect -152 88902 -106 88914
rect -152 87726 -146 88902
rect -112 87726 -106 88902
rect -152 87714 -106 87726
rect 106 88902 152 88914
rect 106 87726 112 88902
rect 146 87726 152 88902
rect 106 87714 152 87726
rect -96 87667 96 87673
rect -96 87633 -84 87667
rect 84 87633 96 87667
rect -96 87627 96 87633
rect -96 87559 96 87565
rect -96 87525 -84 87559
rect 84 87525 96 87559
rect -96 87519 96 87525
rect -152 87466 -106 87478
rect -152 86290 -146 87466
rect -112 86290 -106 87466
rect -152 86278 -106 86290
rect 106 87466 152 87478
rect 106 86290 112 87466
rect 146 86290 152 87466
rect 106 86278 152 86290
rect -96 86231 96 86237
rect -96 86197 -84 86231
rect 84 86197 96 86231
rect -96 86191 96 86197
rect -96 86123 96 86129
rect -96 86089 -84 86123
rect 84 86089 96 86123
rect -96 86083 96 86089
rect -152 86030 -106 86042
rect -152 84854 -146 86030
rect -112 84854 -106 86030
rect -152 84842 -106 84854
rect 106 86030 152 86042
rect 106 84854 112 86030
rect 146 84854 152 86030
rect 106 84842 152 84854
rect -96 84795 96 84801
rect -96 84761 -84 84795
rect 84 84761 96 84795
rect -96 84755 96 84761
rect -96 84687 96 84693
rect -96 84653 -84 84687
rect 84 84653 96 84687
rect -96 84647 96 84653
rect -152 84594 -106 84606
rect -152 83418 -146 84594
rect -112 83418 -106 84594
rect -152 83406 -106 83418
rect 106 84594 152 84606
rect 106 83418 112 84594
rect 146 83418 152 84594
rect 106 83406 152 83418
rect -96 83359 96 83365
rect -96 83325 -84 83359
rect 84 83325 96 83359
rect -96 83319 96 83325
rect -96 83251 96 83257
rect -96 83217 -84 83251
rect 84 83217 96 83251
rect -96 83211 96 83217
rect -152 83158 -106 83170
rect -152 81982 -146 83158
rect -112 81982 -106 83158
rect -152 81970 -106 81982
rect 106 83158 152 83170
rect 106 81982 112 83158
rect 146 81982 152 83158
rect 106 81970 152 81982
rect -96 81923 96 81929
rect -96 81889 -84 81923
rect 84 81889 96 81923
rect -96 81883 96 81889
rect -96 81815 96 81821
rect -96 81781 -84 81815
rect 84 81781 96 81815
rect -96 81775 96 81781
rect -152 81722 -106 81734
rect -152 80546 -146 81722
rect -112 80546 -106 81722
rect -152 80534 -106 80546
rect 106 81722 152 81734
rect 106 80546 112 81722
rect 146 80546 152 81722
rect 106 80534 152 80546
rect -96 80487 96 80493
rect -96 80453 -84 80487
rect 84 80453 96 80487
rect -96 80447 96 80453
rect -96 80379 96 80385
rect -96 80345 -84 80379
rect 84 80345 96 80379
rect -96 80339 96 80345
rect -152 80286 -106 80298
rect -152 79110 -146 80286
rect -112 79110 -106 80286
rect -152 79098 -106 79110
rect 106 80286 152 80298
rect 106 79110 112 80286
rect 146 79110 152 80286
rect 106 79098 152 79110
rect -96 79051 96 79057
rect -96 79017 -84 79051
rect 84 79017 96 79051
rect -96 79011 96 79017
rect -96 78943 96 78949
rect -96 78909 -84 78943
rect 84 78909 96 78943
rect -96 78903 96 78909
rect -152 78850 -106 78862
rect -152 77674 -146 78850
rect -112 77674 -106 78850
rect -152 77662 -106 77674
rect 106 78850 152 78862
rect 106 77674 112 78850
rect 146 77674 152 78850
rect 106 77662 152 77674
rect -96 77615 96 77621
rect -96 77581 -84 77615
rect 84 77581 96 77615
rect -96 77575 96 77581
rect -96 77507 96 77513
rect -96 77473 -84 77507
rect 84 77473 96 77507
rect -96 77467 96 77473
rect -152 77414 -106 77426
rect -152 76238 -146 77414
rect -112 76238 -106 77414
rect -152 76226 -106 76238
rect 106 77414 152 77426
rect 106 76238 112 77414
rect 146 76238 152 77414
rect 106 76226 152 76238
rect -96 76179 96 76185
rect -96 76145 -84 76179
rect 84 76145 96 76179
rect -96 76139 96 76145
rect -96 76071 96 76077
rect -96 76037 -84 76071
rect 84 76037 96 76071
rect -96 76031 96 76037
rect -152 75978 -106 75990
rect -152 74802 -146 75978
rect -112 74802 -106 75978
rect -152 74790 -106 74802
rect 106 75978 152 75990
rect 106 74802 112 75978
rect 146 74802 152 75978
rect 106 74790 152 74802
rect -96 74743 96 74749
rect -96 74709 -84 74743
rect 84 74709 96 74743
rect -96 74703 96 74709
rect -96 74635 96 74641
rect -96 74601 -84 74635
rect 84 74601 96 74635
rect -96 74595 96 74601
rect -152 74542 -106 74554
rect -152 73366 -146 74542
rect -112 73366 -106 74542
rect -152 73354 -106 73366
rect 106 74542 152 74554
rect 106 73366 112 74542
rect 146 73366 152 74542
rect 106 73354 152 73366
rect -96 73307 96 73313
rect -96 73273 -84 73307
rect 84 73273 96 73307
rect -96 73267 96 73273
rect -96 73199 96 73205
rect -96 73165 -84 73199
rect 84 73165 96 73199
rect -96 73159 96 73165
rect -152 73106 -106 73118
rect -152 71930 -146 73106
rect -112 71930 -106 73106
rect -152 71918 -106 71930
rect 106 73106 152 73118
rect 106 71930 112 73106
rect 146 71930 152 73106
rect 106 71918 152 71930
rect -96 71871 96 71877
rect -96 71837 -84 71871
rect 84 71837 96 71871
rect -96 71831 96 71837
rect -96 71763 96 71769
rect -96 71729 -84 71763
rect 84 71729 96 71763
rect -96 71723 96 71729
rect -152 71670 -106 71682
rect -152 70494 -146 71670
rect -112 70494 -106 71670
rect -152 70482 -106 70494
rect 106 71670 152 71682
rect 106 70494 112 71670
rect 146 70494 152 71670
rect 106 70482 152 70494
rect -96 70435 96 70441
rect -96 70401 -84 70435
rect 84 70401 96 70435
rect -96 70395 96 70401
rect -96 70327 96 70333
rect -96 70293 -84 70327
rect 84 70293 96 70327
rect -96 70287 96 70293
rect -152 70234 -106 70246
rect -152 69058 -146 70234
rect -112 69058 -106 70234
rect -152 69046 -106 69058
rect 106 70234 152 70246
rect 106 69058 112 70234
rect 146 69058 152 70234
rect 106 69046 152 69058
rect -96 68999 96 69005
rect -96 68965 -84 68999
rect 84 68965 96 68999
rect -96 68959 96 68965
rect -96 68891 96 68897
rect -96 68857 -84 68891
rect 84 68857 96 68891
rect -96 68851 96 68857
rect -152 68798 -106 68810
rect -152 67622 -146 68798
rect -112 67622 -106 68798
rect -152 67610 -106 67622
rect 106 68798 152 68810
rect 106 67622 112 68798
rect 146 67622 152 68798
rect 106 67610 152 67622
rect -96 67563 96 67569
rect -96 67529 -84 67563
rect 84 67529 96 67563
rect -96 67523 96 67529
rect -96 67455 96 67461
rect -96 67421 -84 67455
rect 84 67421 96 67455
rect -96 67415 96 67421
rect -152 67362 -106 67374
rect -152 66186 -146 67362
rect -112 66186 -106 67362
rect -152 66174 -106 66186
rect 106 67362 152 67374
rect 106 66186 112 67362
rect 146 66186 152 67362
rect 106 66174 152 66186
rect -96 66127 96 66133
rect -96 66093 -84 66127
rect 84 66093 96 66127
rect -96 66087 96 66093
rect -96 66019 96 66025
rect -96 65985 -84 66019
rect 84 65985 96 66019
rect -96 65979 96 65985
rect -152 65926 -106 65938
rect -152 64750 -146 65926
rect -112 64750 -106 65926
rect -152 64738 -106 64750
rect 106 65926 152 65938
rect 106 64750 112 65926
rect 146 64750 152 65926
rect 106 64738 152 64750
rect -96 64691 96 64697
rect -96 64657 -84 64691
rect 84 64657 96 64691
rect -96 64651 96 64657
rect -96 64583 96 64589
rect -96 64549 -84 64583
rect 84 64549 96 64583
rect -96 64543 96 64549
rect -152 64490 -106 64502
rect -152 63314 -146 64490
rect -112 63314 -106 64490
rect -152 63302 -106 63314
rect 106 64490 152 64502
rect 106 63314 112 64490
rect 146 63314 152 64490
rect 106 63302 152 63314
rect -96 63255 96 63261
rect -96 63221 -84 63255
rect 84 63221 96 63255
rect -96 63215 96 63221
rect -96 63147 96 63153
rect -96 63113 -84 63147
rect 84 63113 96 63147
rect -96 63107 96 63113
rect -152 63054 -106 63066
rect -152 61878 -146 63054
rect -112 61878 -106 63054
rect -152 61866 -106 61878
rect 106 63054 152 63066
rect 106 61878 112 63054
rect 146 61878 152 63054
rect 106 61866 152 61878
rect -96 61819 96 61825
rect -96 61785 -84 61819
rect 84 61785 96 61819
rect -96 61779 96 61785
rect -96 61711 96 61717
rect -96 61677 -84 61711
rect 84 61677 96 61711
rect -96 61671 96 61677
rect -152 61618 -106 61630
rect -152 60442 -146 61618
rect -112 60442 -106 61618
rect -152 60430 -106 60442
rect 106 61618 152 61630
rect 106 60442 112 61618
rect 146 60442 152 61618
rect 106 60430 152 60442
rect -96 60383 96 60389
rect -96 60349 -84 60383
rect 84 60349 96 60383
rect -96 60343 96 60349
rect -96 60275 96 60281
rect -96 60241 -84 60275
rect 84 60241 96 60275
rect -96 60235 96 60241
rect -152 60182 -106 60194
rect -152 59006 -146 60182
rect -112 59006 -106 60182
rect -152 58994 -106 59006
rect 106 60182 152 60194
rect 106 59006 112 60182
rect 146 59006 152 60182
rect 106 58994 152 59006
rect -96 58947 96 58953
rect -96 58913 -84 58947
rect 84 58913 96 58947
rect -96 58907 96 58913
rect -96 58839 96 58845
rect -96 58805 -84 58839
rect 84 58805 96 58839
rect -96 58799 96 58805
rect -152 58746 -106 58758
rect -152 57570 -146 58746
rect -112 57570 -106 58746
rect -152 57558 -106 57570
rect 106 58746 152 58758
rect 106 57570 112 58746
rect 146 57570 152 58746
rect 106 57558 152 57570
rect -96 57511 96 57517
rect -96 57477 -84 57511
rect 84 57477 96 57511
rect -96 57471 96 57477
rect -96 57403 96 57409
rect -96 57369 -84 57403
rect 84 57369 96 57403
rect -96 57363 96 57369
rect -152 57310 -106 57322
rect -152 56134 -146 57310
rect -112 56134 -106 57310
rect -152 56122 -106 56134
rect 106 57310 152 57322
rect 106 56134 112 57310
rect 146 56134 152 57310
rect 106 56122 152 56134
rect -96 56075 96 56081
rect -96 56041 -84 56075
rect 84 56041 96 56075
rect -96 56035 96 56041
rect -96 55967 96 55973
rect -96 55933 -84 55967
rect 84 55933 96 55967
rect -96 55927 96 55933
rect -152 55874 -106 55886
rect -152 54698 -146 55874
rect -112 54698 -106 55874
rect -152 54686 -106 54698
rect 106 55874 152 55886
rect 106 54698 112 55874
rect 146 54698 152 55874
rect 106 54686 152 54698
rect -96 54639 96 54645
rect -96 54605 -84 54639
rect 84 54605 96 54639
rect -96 54599 96 54605
rect -96 54531 96 54537
rect -96 54497 -84 54531
rect 84 54497 96 54531
rect -96 54491 96 54497
rect -152 54438 -106 54450
rect -152 53262 -146 54438
rect -112 53262 -106 54438
rect -152 53250 -106 53262
rect 106 54438 152 54450
rect 106 53262 112 54438
rect 146 53262 152 54438
rect 106 53250 152 53262
rect -96 53203 96 53209
rect -96 53169 -84 53203
rect 84 53169 96 53203
rect -96 53163 96 53169
rect -96 53095 96 53101
rect -96 53061 -84 53095
rect 84 53061 96 53095
rect -96 53055 96 53061
rect -152 53002 -106 53014
rect -152 51826 -146 53002
rect -112 51826 -106 53002
rect -152 51814 -106 51826
rect 106 53002 152 53014
rect 106 51826 112 53002
rect 146 51826 152 53002
rect 106 51814 152 51826
rect -96 51767 96 51773
rect -96 51733 -84 51767
rect 84 51733 96 51767
rect -96 51727 96 51733
rect -96 51659 96 51665
rect -96 51625 -84 51659
rect 84 51625 96 51659
rect -96 51619 96 51625
rect -152 51566 -106 51578
rect -152 50390 -146 51566
rect -112 50390 -106 51566
rect -152 50378 -106 50390
rect 106 51566 152 51578
rect 106 50390 112 51566
rect 146 50390 152 51566
rect 106 50378 152 50390
rect -96 50331 96 50337
rect -96 50297 -84 50331
rect 84 50297 96 50331
rect -96 50291 96 50297
rect -96 50223 96 50229
rect -96 50189 -84 50223
rect 84 50189 96 50223
rect -96 50183 96 50189
rect -152 50130 -106 50142
rect -152 48954 -146 50130
rect -112 48954 -106 50130
rect -152 48942 -106 48954
rect 106 50130 152 50142
rect 106 48954 112 50130
rect 146 48954 152 50130
rect 106 48942 152 48954
rect -96 48895 96 48901
rect -96 48861 -84 48895
rect 84 48861 96 48895
rect -96 48855 96 48861
rect -96 48787 96 48793
rect -96 48753 -84 48787
rect 84 48753 96 48787
rect -96 48747 96 48753
rect -152 48694 -106 48706
rect -152 47518 -146 48694
rect -112 47518 -106 48694
rect -152 47506 -106 47518
rect 106 48694 152 48706
rect 106 47518 112 48694
rect 146 47518 152 48694
rect 106 47506 152 47518
rect -96 47459 96 47465
rect -96 47425 -84 47459
rect 84 47425 96 47459
rect -96 47419 96 47425
rect -96 47351 96 47357
rect -96 47317 -84 47351
rect 84 47317 96 47351
rect -96 47311 96 47317
rect -152 47258 -106 47270
rect -152 46082 -146 47258
rect -112 46082 -106 47258
rect -152 46070 -106 46082
rect 106 47258 152 47270
rect 106 46082 112 47258
rect 146 46082 152 47258
rect 106 46070 152 46082
rect -96 46023 96 46029
rect -96 45989 -84 46023
rect 84 45989 96 46023
rect -96 45983 96 45989
rect -96 45915 96 45921
rect -96 45881 -84 45915
rect 84 45881 96 45915
rect -96 45875 96 45881
rect -152 45822 -106 45834
rect -152 44646 -146 45822
rect -112 44646 -106 45822
rect -152 44634 -106 44646
rect 106 45822 152 45834
rect 106 44646 112 45822
rect 146 44646 152 45822
rect 106 44634 152 44646
rect -96 44587 96 44593
rect -96 44553 -84 44587
rect 84 44553 96 44587
rect -96 44547 96 44553
rect -96 44479 96 44485
rect -96 44445 -84 44479
rect 84 44445 96 44479
rect -96 44439 96 44445
rect -152 44386 -106 44398
rect -152 43210 -146 44386
rect -112 43210 -106 44386
rect -152 43198 -106 43210
rect 106 44386 152 44398
rect 106 43210 112 44386
rect 146 43210 152 44386
rect 106 43198 152 43210
rect -96 43151 96 43157
rect -96 43117 -84 43151
rect 84 43117 96 43151
rect -96 43111 96 43117
rect -96 43043 96 43049
rect -96 43009 -84 43043
rect 84 43009 96 43043
rect -96 43003 96 43009
rect -152 42950 -106 42962
rect -152 41774 -146 42950
rect -112 41774 -106 42950
rect -152 41762 -106 41774
rect 106 42950 152 42962
rect 106 41774 112 42950
rect 146 41774 152 42950
rect 106 41762 152 41774
rect -96 41715 96 41721
rect -96 41681 -84 41715
rect 84 41681 96 41715
rect -96 41675 96 41681
rect -96 41607 96 41613
rect -96 41573 -84 41607
rect 84 41573 96 41607
rect -96 41567 96 41573
rect -152 41514 -106 41526
rect -152 40338 -146 41514
rect -112 40338 -106 41514
rect -152 40326 -106 40338
rect 106 41514 152 41526
rect 106 40338 112 41514
rect 146 40338 152 41514
rect 106 40326 152 40338
rect -96 40279 96 40285
rect -96 40245 -84 40279
rect 84 40245 96 40279
rect -96 40239 96 40245
rect -96 40171 96 40177
rect -96 40137 -84 40171
rect 84 40137 96 40171
rect -96 40131 96 40137
rect -152 40078 -106 40090
rect -152 38902 -146 40078
rect -112 38902 -106 40078
rect -152 38890 -106 38902
rect 106 40078 152 40090
rect 106 38902 112 40078
rect 146 38902 152 40078
rect 106 38890 152 38902
rect -96 38843 96 38849
rect -96 38809 -84 38843
rect 84 38809 96 38843
rect -96 38803 96 38809
rect -96 38735 96 38741
rect -96 38701 -84 38735
rect 84 38701 96 38735
rect -96 38695 96 38701
rect -152 38642 -106 38654
rect -152 37466 -146 38642
rect -112 37466 -106 38642
rect -152 37454 -106 37466
rect 106 38642 152 38654
rect 106 37466 112 38642
rect 146 37466 152 38642
rect 106 37454 152 37466
rect -96 37407 96 37413
rect -96 37373 -84 37407
rect 84 37373 96 37407
rect -96 37367 96 37373
rect -96 37299 96 37305
rect -96 37265 -84 37299
rect 84 37265 96 37299
rect -96 37259 96 37265
rect -152 37206 -106 37218
rect -152 36030 -146 37206
rect -112 36030 -106 37206
rect -152 36018 -106 36030
rect 106 37206 152 37218
rect 106 36030 112 37206
rect 146 36030 152 37206
rect 106 36018 152 36030
rect -96 35971 96 35977
rect -96 35937 -84 35971
rect 84 35937 96 35971
rect -96 35931 96 35937
rect -96 35863 96 35869
rect -96 35829 -84 35863
rect 84 35829 96 35863
rect -96 35823 96 35829
rect -152 35770 -106 35782
rect -152 34594 -146 35770
rect -112 34594 -106 35770
rect -152 34582 -106 34594
rect 106 35770 152 35782
rect 106 34594 112 35770
rect 146 34594 152 35770
rect 106 34582 152 34594
rect -96 34535 96 34541
rect -96 34501 -84 34535
rect 84 34501 96 34535
rect -96 34495 96 34501
rect -96 34427 96 34433
rect -96 34393 -84 34427
rect 84 34393 96 34427
rect -96 34387 96 34393
rect -152 34334 -106 34346
rect -152 33158 -146 34334
rect -112 33158 -106 34334
rect -152 33146 -106 33158
rect 106 34334 152 34346
rect 106 33158 112 34334
rect 146 33158 152 34334
rect 106 33146 152 33158
rect -96 33099 96 33105
rect -96 33065 -84 33099
rect 84 33065 96 33099
rect -96 33059 96 33065
rect -96 32991 96 32997
rect -96 32957 -84 32991
rect 84 32957 96 32991
rect -96 32951 96 32957
rect -152 32898 -106 32910
rect -152 31722 -146 32898
rect -112 31722 -106 32898
rect -152 31710 -106 31722
rect 106 32898 152 32910
rect 106 31722 112 32898
rect 146 31722 152 32898
rect 106 31710 152 31722
rect -96 31663 96 31669
rect -96 31629 -84 31663
rect 84 31629 96 31663
rect -96 31623 96 31629
rect -96 31555 96 31561
rect -96 31521 -84 31555
rect 84 31521 96 31555
rect -96 31515 96 31521
rect -152 31462 -106 31474
rect -152 30286 -146 31462
rect -112 30286 -106 31462
rect -152 30274 -106 30286
rect 106 31462 152 31474
rect 106 30286 112 31462
rect 146 30286 152 31462
rect 106 30274 152 30286
rect -96 30227 96 30233
rect -96 30193 -84 30227
rect 84 30193 96 30227
rect -96 30187 96 30193
rect -96 30119 96 30125
rect -96 30085 -84 30119
rect 84 30085 96 30119
rect -96 30079 96 30085
rect -152 30026 -106 30038
rect -152 28850 -146 30026
rect -112 28850 -106 30026
rect -152 28838 -106 28850
rect 106 30026 152 30038
rect 106 28850 112 30026
rect 146 28850 152 30026
rect 106 28838 152 28850
rect -96 28791 96 28797
rect -96 28757 -84 28791
rect 84 28757 96 28791
rect -96 28751 96 28757
rect -96 28683 96 28689
rect -96 28649 -84 28683
rect 84 28649 96 28683
rect -96 28643 96 28649
rect -152 28590 -106 28602
rect -152 27414 -146 28590
rect -112 27414 -106 28590
rect -152 27402 -106 27414
rect 106 28590 152 28602
rect 106 27414 112 28590
rect 146 27414 152 28590
rect 106 27402 152 27414
rect -96 27355 96 27361
rect -96 27321 -84 27355
rect 84 27321 96 27355
rect -96 27315 96 27321
rect -96 27247 96 27253
rect -96 27213 -84 27247
rect 84 27213 96 27247
rect -96 27207 96 27213
rect -152 27154 -106 27166
rect -152 25978 -146 27154
rect -112 25978 -106 27154
rect -152 25966 -106 25978
rect 106 27154 152 27166
rect 106 25978 112 27154
rect 146 25978 152 27154
rect 106 25966 152 25978
rect -96 25919 96 25925
rect -96 25885 -84 25919
rect 84 25885 96 25919
rect -96 25879 96 25885
rect -96 25811 96 25817
rect -96 25777 -84 25811
rect 84 25777 96 25811
rect -96 25771 96 25777
rect -152 25718 -106 25730
rect -152 24542 -146 25718
rect -112 24542 -106 25718
rect -152 24530 -106 24542
rect 106 25718 152 25730
rect 106 24542 112 25718
rect 146 24542 152 25718
rect 106 24530 152 24542
rect -96 24483 96 24489
rect -96 24449 -84 24483
rect 84 24449 96 24483
rect -96 24443 96 24449
rect -96 24375 96 24381
rect -96 24341 -84 24375
rect 84 24341 96 24375
rect -96 24335 96 24341
rect -152 24282 -106 24294
rect -152 23106 -146 24282
rect -112 23106 -106 24282
rect -152 23094 -106 23106
rect 106 24282 152 24294
rect 106 23106 112 24282
rect 146 23106 152 24282
rect 106 23094 152 23106
rect -96 23047 96 23053
rect -96 23013 -84 23047
rect 84 23013 96 23047
rect -96 23007 96 23013
rect -96 22939 96 22945
rect -96 22905 -84 22939
rect 84 22905 96 22939
rect -96 22899 96 22905
rect -152 22846 -106 22858
rect -152 21670 -146 22846
rect -112 21670 -106 22846
rect -152 21658 -106 21670
rect 106 22846 152 22858
rect 106 21670 112 22846
rect 146 21670 152 22846
rect 106 21658 152 21670
rect -96 21611 96 21617
rect -96 21577 -84 21611
rect 84 21577 96 21611
rect -96 21571 96 21577
rect -96 21503 96 21509
rect -96 21469 -84 21503
rect 84 21469 96 21503
rect -96 21463 96 21469
rect -152 21410 -106 21422
rect -152 20234 -146 21410
rect -112 20234 -106 21410
rect -152 20222 -106 20234
rect 106 21410 152 21422
rect 106 20234 112 21410
rect 146 20234 152 21410
rect 106 20222 152 20234
rect -96 20175 96 20181
rect -96 20141 -84 20175
rect 84 20141 96 20175
rect -96 20135 96 20141
rect -96 20067 96 20073
rect -96 20033 -84 20067
rect 84 20033 96 20067
rect -96 20027 96 20033
rect -152 19974 -106 19986
rect -152 18798 -146 19974
rect -112 18798 -106 19974
rect -152 18786 -106 18798
rect 106 19974 152 19986
rect 106 18798 112 19974
rect 146 18798 152 19974
rect 106 18786 152 18798
rect -96 18739 96 18745
rect -96 18705 -84 18739
rect 84 18705 96 18739
rect -96 18699 96 18705
rect -96 18631 96 18637
rect -96 18597 -84 18631
rect 84 18597 96 18631
rect -96 18591 96 18597
rect -152 18538 -106 18550
rect -152 17362 -146 18538
rect -112 17362 -106 18538
rect -152 17350 -106 17362
rect 106 18538 152 18550
rect 106 17362 112 18538
rect 146 17362 152 18538
rect 106 17350 152 17362
rect -96 17303 96 17309
rect -96 17269 -84 17303
rect 84 17269 96 17303
rect -96 17263 96 17269
rect -96 17195 96 17201
rect -96 17161 -84 17195
rect 84 17161 96 17195
rect -96 17155 96 17161
rect -152 17102 -106 17114
rect -152 15926 -146 17102
rect -112 15926 -106 17102
rect -152 15914 -106 15926
rect 106 17102 152 17114
rect 106 15926 112 17102
rect 146 15926 152 17102
rect 106 15914 152 15926
rect -96 15867 96 15873
rect -96 15833 -84 15867
rect 84 15833 96 15867
rect -96 15827 96 15833
rect -96 15759 96 15765
rect -96 15725 -84 15759
rect 84 15725 96 15759
rect -96 15719 96 15725
rect -152 15666 -106 15678
rect -152 14490 -146 15666
rect -112 14490 -106 15666
rect -152 14478 -106 14490
rect 106 15666 152 15678
rect 106 14490 112 15666
rect 146 14490 152 15666
rect 106 14478 152 14490
rect -96 14431 96 14437
rect -96 14397 -84 14431
rect 84 14397 96 14431
rect -96 14391 96 14397
rect -96 14323 96 14329
rect -96 14289 -84 14323
rect 84 14289 96 14323
rect -96 14283 96 14289
rect -152 14230 -106 14242
rect -152 13054 -146 14230
rect -112 13054 -106 14230
rect -152 13042 -106 13054
rect 106 14230 152 14242
rect 106 13054 112 14230
rect 146 13054 152 14230
rect 106 13042 152 13054
rect -96 12995 96 13001
rect -96 12961 -84 12995
rect 84 12961 96 12995
rect -96 12955 96 12961
rect -96 12887 96 12893
rect -96 12853 -84 12887
rect 84 12853 96 12887
rect -96 12847 96 12853
rect -152 12794 -106 12806
rect -152 11618 -146 12794
rect -112 11618 -106 12794
rect -152 11606 -106 11618
rect 106 12794 152 12806
rect 106 11618 112 12794
rect 146 11618 152 12794
rect 106 11606 152 11618
rect -96 11559 96 11565
rect -96 11525 -84 11559
rect 84 11525 96 11559
rect -96 11519 96 11525
rect -96 11451 96 11457
rect -96 11417 -84 11451
rect 84 11417 96 11451
rect -96 11411 96 11417
rect -152 11358 -106 11370
rect -152 10182 -146 11358
rect -112 10182 -106 11358
rect -152 10170 -106 10182
rect 106 11358 152 11370
rect 106 10182 112 11358
rect 146 10182 152 11358
rect 106 10170 152 10182
rect -96 10123 96 10129
rect -96 10089 -84 10123
rect 84 10089 96 10123
rect -96 10083 96 10089
rect -96 10015 96 10021
rect -96 9981 -84 10015
rect 84 9981 96 10015
rect -96 9975 96 9981
rect -152 9922 -106 9934
rect -152 8746 -146 9922
rect -112 8746 -106 9922
rect -152 8734 -106 8746
rect 106 9922 152 9934
rect 106 8746 112 9922
rect 146 8746 152 9922
rect 106 8734 152 8746
rect -96 8687 96 8693
rect -96 8653 -84 8687
rect 84 8653 96 8687
rect -96 8647 96 8653
rect -96 8579 96 8585
rect -96 8545 -84 8579
rect 84 8545 96 8579
rect -96 8539 96 8545
rect -152 8486 -106 8498
rect -152 7310 -146 8486
rect -112 7310 -106 8486
rect -152 7298 -106 7310
rect 106 8486 152 8498
rect 106 7310 112 8486
rect 146 7310 152 8486
rect 106 7298 152 7310
rect -96 7251 96 7257
rect -96 7217 -84 7251
rect 84 7217 96 7251
rect -96 7211 96 7217
rect -96 7143 96 7149
rect -96 7109 -84 7143
rect 84 7109 96 7143
rect -96 7103 96 7109
rect -152 7050 -106 7062
rect -152 5874 -146 7050
rect -112 5874 -106 7050
rect -152 5862 -106 5874
rect 106 7050 152 7062
rect 106 5874 112 7050
rect 146 5874 152 7050
rect 106 5862 152 5874
rect -96 5815 96 5821
rect -96 5781 -84 5815
rect 84 5781 96 5815
rect -96 5775 96 5781
rect -96 5707 96 5713
rect -96 5673 -84 5707
rect 84 5673 96 5707
rect -96 5667 96 5673
rect -152 5614 -106 5626
rect -152 4438 -146 5614
rect -112 4438 -106 5614
rect -152 4426 -106 4438
rect 106 5614 152 5626
rect 106 4438 112 5614
rect 146 4438 152 5614
rect 106 4426 152 4438
rect -96 4379 96 4385
rect -96 4345 -84 4379
rect 84 4345 96 4379
rect -96 4339 96 4345
rect -96 4271 96 4277
rect -96 4237 -84 4271
rect 84 4237 96 4271
rect -96 4231 96 4237
rect -152 4178 -106 4190
rect -152 3002 -146 4178
rect -112 3002 -106 4178
rect -152 2990 -106 3002
rect 106 4178 152 4190
rect 106 3002 112 4178
rect 146 3002 152 4178
rect 106 2990 152 3002
rect -96 2943 96 2949
rect -96 2909 -84 2943
rect 84 2909 96 2943
rect -96 2903 96 2909
rect -96 2835 96 2841
rect -96 2801 -84 2835
rect 84 2801 96 2835
rect -96 2795 96 2801
rect -152 2742 -106 2754
rect -152 1566 -146 2742
rect -112 1566 -106 2742
rect -152 1554 -106 1566
rect 106 2742 152 2754
rect 106 1566 112 2742
rect 146 1566 152 2742
rect 106 1554 152 1566
rect -96 1507 96 1513
rect -96 1473 -84 1507
rect 84 1473 96 1507
rect -96 1467 96 1473
rect -96 1399 96 1405
rect -96 1365 -84 1399
rect 84 1365 96 1399
rect -96 1359 96 1365
rect -152 1306 -106 1318
rect -152 130 -146 1306
rect -112 130 -106 1306
rect -152 118 -106 130
rect 106 1306 152 1318
rect 106 130 112 1306
rect 146 130 152 1306
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -1306 -146 -130
rect -112 -1306 -106 -130
rect -152 -1318 -106 -1306
rect 106 -130 152 -118
rect 106 -1306 112 -130
rect 146 -1306 152 -130
rect 106 -1318 152 -1306
rect -96 -1365 96 -1359
rect -96 -1399 -84 -1365
rect 84 -1399 96 -1365
rect -96 -1405 96 -1399
rect -96 -1473 96 -1467
rect -96 -1507 -84 -1473
rect 84 -1507 96 -1473
rect -96 -1513 96 -1507
rect -152 -1566 -106 -1554
rect -152 -2742 -146 -1566
rect -112 -2742 -106 -1566
rect -152 -2754 -106 -2742
rect 106 -1566 152 -1554
rect 106 -2742 112 -1566
rect 146 -2742 152 -1566
rect 106 -2754 152 -2742
rect -96 -2801 96 -2795
rect -96 -2835 -84 -2801
rect 84 -2835 96 -2801
rect -96 -2841 96 -2835
rect -96 -2909 96 -2903
rect -96 -2943 -84 -2909
rect 84 -2943 96 -2909
rect -96 -2949 96 -2943
rect -152 -3002 -106 -2990
rect -152 -4178 -146 -3002
rect -112 -4178 -106 -3002
rect -152 -4190 -106 -4178
rect 106 -3002 152 -2990
rect 106 -4178 112 -3002
rect 146 -4178 152 -3002
rect 106 -4190 152 -4178
rect -96 -4237 96 -4231
rect -96 -4271 -84 -4237
rect 84 -4271 96 -4237
rect -96 -4277 96 -4271
rect -96 -4345 96 -4339
rect -96 -4379 -84 -4345
rect 84 -4379 96 -4345
rect -96 -4385 96 -4379
rect -152 -4438 -106 -4426
rect -152 -5614 -146 -4438
rect -112 -5614 -106 -4438
rect -152 -5626 -106 -5614
rect 106 -4438 152 -4426
rect 106 -5614 112 -4438
rect 146 -5614 152 -4438
rect 106 -5626 152 -5614
rect -96 -5673 96 -5667
rect -96 -5707 -84 -5673
rect 84 -5707 96 -5673
rect -96 -5713 96 -5707
rect -96 -5781 96 -5775
rect -96 -5815 -84 -5781
rect 84 -5815 96 -5781
rect -96 -5821 96 -5815
rect -152 -5874 -106 -5862
rect -152 -7050 -146 -5874
rect -112 -7050 -106 -5874
rect -152 -7062 -106 -7050
rect 106 -5874 152 -5862
rect 106 -7050 112 -5874
rect 146 -7050 152 -5874
rect 106 -7062 152 -7050
rect -96 -7109 96 -7103
rect -96 -7143 -84 -7109
rect 84 -7143 96 -7109
rect -96 -7149 96 -7143
rect -96 -7217 96 -7211
rect -96 -7251 -84 -7217
rect 84 -7251 96 -7217
rect -96 -7257 96 -7251
rect -152 -7310 -106 -7298
rect -152 -8486 -146 -7310
rect -112 -8486 -106 -7310
rect -152 -8498 -106 -8486
rect 106 -7310 152 -7298
rect 106 -8486 112 -7310
rect 146 -8486 152 -7310
rect 106 -8498 152 -8486
rect -96 -8545 96 -8539
rect -96 -8579 -84 -8545
rect 84 -8579 96 -8545
rect -96 -8585 96 -8579
rect -96 -8653 96 -8647
rect -96 -8687 -84 -8653
rect 84 -8687 96 -8653
rect -96 -8693 96 -8687
rect -152 -8746 -106 -8734
rect -152 -9922 -146 -8746
rect -112 -9922 -106 -8746
rect -152 -9934 -106 -9922
rect 106 -8746 152 -8734
rect 106 -9922 112 -8746
rect 146 -9922 152 -8746
rect 106 -9934 152 -9922
rect -96 -9981 96 -9975
rect -96 -10015 -84 -9981
rect 84 -10015 96 -9981
rect -96 -10021 96 -10015
rect -96 -10089 96 -10083
rect -96 -10123 -84 -10089
rect 84 -10123 96 -10089
rect -96 -10129 96 -10123
rect -152 -10182 -106 -10170
rect -152 -11358 -146 -10182
rect -112 -11358 -106 -10182
rect -152 -11370 -106 -11358
rect 106 -10182 152 -10170
rect 106 -11358 112 -10182
rect 146 -11358 152 -10182
rect 106 -11370 152 -11358
rect -96 -11417 96 -11411
rect -96 -11451 -84 -11417
rect 84 -11451 96 -11417
rect -96 -11457 96 -11451
rect -96 -11525 96 -11519
rect -96 -11559 -84 -11525
rect 84 -11559 96 -11525
rect -96 -11565 96 -11559
rect -152 -11618 -106 -11606
rect -152 -12794 -146 -11618
rect -112 -12794 -106 -11618
rect -152 -12806 -106 -12794
rect 106 -11618 152 -11606
rect 106 -12794 112 -11618
rect 146 -12794 152 -11618
rect 106 -12806 152 -12794
rect -96 -12853 96 -12847
rect -96 -12887 -84 -12853
rect 84 -12887 96 -12853
rect -96 -12893 96 -12887
rect -96 -12961 96 -12955
rect -96 -12995 -84 -12961
rect 84 -12995 96 -12961
rect -96 -13001 96 -12995
rect -152 -13054 -106 -13042
rect -152 -14230 -146 -13054
rect -112 -14230 -106 -13054
rect -152 -14242 -106 -14230
rect 106 -13054 152 -13042
rect 106 -14230 112 -13054
rect 146 -14230 152 -13054
rect 106 -14242 152 -14230
rect -96 -14289 96 -14283
rect -96 -14323 -84 -14289
rect 84 -14323 96 -14289
rect -96 -14329 96 -14323
rect -96 -14397 96 -14391
rect -96 -14431 -84 -14397
rect 84 -14431 96 -14397
rect -96 -14437 96 -14431
rect -152 -14490 -106 -14478
rect -152 -15666 -146 -14490
rect -112 -15666 -106 -14490
rect -152 -15678 -106 -15666
rect 106 -14490 152 -14478
rect 106 -15666 112 -14490
rect 146 -15666 152 -14490
rect 106 -15678 152 -15666
rect -96 -15725 96 -15719
rect -96 -15759 -84 -15725
rect 84 -15759 96 -15725
rect -96 -15765 96 -15759
rect -96 -15833 96 -15827
rect -96 -15867 -84 -15833
rect 84 -15867 96 -15833
rect -96 -15873 96 -15867
rect -152 -15926 -106 -15914
rect -152 -17102 -146 -15926
rect -112 -17102 -106 -15926
rect -152 -17114 -106 -17102
rect 106 -15926 152 -15914
rect 106 -17102 112 -15926
rect 146 -17102 152 -15926
rect 106 -17114 152 -17102
rect -96 -17161 96 -17155
rect -96 -17195 -84 -17161
rect 84 -17195 96 -17161
rect -96 -17201 96 -17195
rect -96 -17269 96 -17263
rect -96 -17303 -84 -17269
rect 84 -17303 96 -17269
rect -96 -17309 96 -17303
rect -152 -17362 -106 -17350
rect -152 -18538 -146 -17362
rect -112 -18538 -106 -17362
rect -152 -18550 -106 -18538
rect 106 -17362 152 -17350
rect 106 -18538 112 -17362
rect 146 -18538 152 -17362
rect 106 -18550 152 -18538
rect -96 -18597 96 -18591
rect -96 -18631 -84 -18597
rect 84 -18631 96 -18597
rect -96 -18637 96 -18631
rect -96 -18705 96 -18699
rect -96 -18739 -84 -18705
rect 84 -18739 96 -18705
rect -96 -18745 96 -18739
rect -152 -18798 -106 -18786
rect -152 -19974 -146 -18798
rect -112 -19974 -106 -18798
rect -152 -19986 -106 -19974
rect 106 -18798 152 -18786
rect 106 -19974 112 -18798
rect 146 -19974 152 -18798
rect 106 -19986 152 -19974
rect -96 -20033 96 -20027
rect -96 -20067 -84 -20033
rect 84 -20067 96 -20033
rect -96 -20073 96 -20067
rect -96 -20141 96 -20135
rect -96 -20175 -84 -20141
rect 84 -20175 96 -20141
rect -96 -20181 96 -20175
rect -152 -20234 -106 -20222
rect -152 -21410 -146 -20234
rect -112 -21410 -106 -20234
rect -152 -21422 -106 -21410
rect 106 -20234 152 -20222
rect 106 -21410 112 -20234
rect 146 -21410 152 -20234
rect 106 -21422 152 -21410
rect -96 -21469 96 -21463
rect -96 -21503 -84 -21469
rect 84 -21503 96 -21469
rect -96 -21509 96 -21503
rect -96 -21577 96 -21571
rect -96 -21611 -84 -21577
rect 84 -21611 96 -21577
rect -96 -21617 96 -21611
rect -152 -21670 -106 -21658
rect -152 -22846 -146 -21670
rect -112 -22846 -106 -21670
rect -152 -22858 -106 -22846
rect 106 -21670 152 -21658
rect 106 -22846 112 -21670
rect 146 -22846 152 -21670
rect 106 -22858 152 -22846
rect -96 -22905 96 -22899
rect -96 -22939 -84 -22905
rect 84 -22939 96 -22905
rect -96 -22945 96 -22939
rect -96 -23013 96 -23007
rect -96 -23047 -84 -23013
rect 84 -23047 96 -23013
rect -96 -23053 96 -23047
rect -152 -23106 -106 -23094
rect -152 -24282 -146 -23106
rect -112 -24282 -106 -23106
rect -152 -24294 -106 -24282
rect 106 -23106 152 -23094
rect 106 -24282 112 -23106
rect 146 -24282 152 -23106
rect 106 -24294 152 -24282
rect -96 -24341 96 -24335
rect -96 -24375 -84 -24341
rect 84 -24375 96 -24341
rect -96 -24381 96 -24375
rect -96 -24449 96 -24443
rect -96 -24483 -84 -24449
rect 84 -24483 96 -24449
rect -96 -24489 96 -24483
rect -152 -24542 -106 -24530
rect -152 -25718 -146 -24542
rect -112 -25718 -106 -24542
rect -152 -25730 -106 -25718
rect 106 -24542 152 -24530
rect 106 -25718 112 -24542
rect 146 -25718 152 -24542
rect 106 -25730 152 -25718
rect -96 -25777 96 -25771
rect -96 -25811 -84 -25777
rect 84 -25811 96 -25777
rect -96 -25817 96 -25811
rect -96 -25885 96 -25879
rect -96 -25919 -84 -25885
rect 84 -25919 96 -25885
rect -96 -25925 96 -25919
rect -152 -25978 -106 -25966
rect -152 -27154 -146 -25978
rect -112 -27154 -106 -25978
rect -152 -27166 -106 -27154
rect 106 -25978 152 -25966
rect 106 -27154 112 -25978
rect 146 -27154 152 -25978
rect 106 -27166 152 -27154
rect -96 -27213 96 -27207
rect -96 -27247 -84 -27213
rect 84 -27247 96 -27213
rect -96 -27253 96 -27247
rect -96 -27321 96 -27315
rect -96 -27355 -84 -27321
rect 84 -27355 96 -27321
rect -96 -27361 96 -27355
rect -152 -27414 -106 -27402
rect -152 -28590 -146 -27414
rect -112 -28590 -106 -27414
rect -152 -28602 -106 -28590
rect 106 -27414 152 -27402
rect 106 -28590 112 -27414
rect 146 -28590 152 -27414
rect 106 -28602 152 -28590
rect -96 -28649 96 -28643
rect -96 -28683 -84 -28649
rect 84 -28683 96 -28649
rect -96 -28689 96 -28683
rect -96 -28757 96 -28751
rect -96 -28791 -84 -28757
rect 84 -28791 96 -28757
rect -96 -28797 96 -28791
rect -152 -28850 -106 -28838
rect -152 -30026 -146 -28850
rect -112 -30026 -106 -28850
rect -152 -30038 -106 -30026
rect 106 -28850 152 -28838
rect 106 -30026 112 -28850
rect 146 -30026 152 -28850
rect 106 -30038 152 -30026
rect -96 -30085 96 -30079
rect -96 -30119 -84 -30085
rect 84 -30119 96 -30085
rect -96 -30125 96 -30119
rect -96 -30193 96 -30187
rect -96 -30227 -84 -30193
rect 84 -30227 96 -30193
rect -96 -30233 96 -30227
rect -152 -30286 -106 -30274
rect -152 -31462 -146 -30286
rect -112 -31462 -106 -30286
rect -152 -31474 -106 -31462
rect 106 -30286 152 -30274
rect 106 -31462 112 -30286
rect 146 -31462 152 -30286
rect 106 -31474 152 -31462
rect -96 -31521 96 -31515
rect -96 -31555 -84 -31521
rect 84 -31555 96 -31521
rect -96 -31561 96 -31555
rect -96 -31629 96 -31623
rect -96 -31663 -84 -31629
rect 84 -31663 96 -31629
rect -96 -31669 96 -31663
rect -152 -31722 -106 -31710
rect -152 -32898 -146 -31722
rect -112 -32898 -106 -31722
rect -152 -32910 -106 -32898
rect 106 -31722 152 -31710
rect 106 -32898 112 -31722
rect 146 -32898 152 -31722
rect 106 -32910 152 -32898
rect -96 -32957 96 -32951
rect -96 -32991 -84 -32957
rect 84 -32991 96 -32957
rect -96 -32997 96 -32991
rect -96 -33065 96 -33059
rect -96 -33099 -84 -33065
rect 84 -33099 96 -33065
rect -96 -33105 96 -33099
rect -152 -33158 -106 -33146
rect -152 -34334 -146 -33158
rect -112 -34334 -106 -33158
rect -152 -34346 -106 -34334
rect 106 -33158 152 -33146
rect 106 -34334 112 -33158
rect 146 -34334 152 -33158
rect 106 -34346 152 -34334
rect -96 -34393 96 -34387
rect -96 -34427 -84 -34393
rect 84 -34427 96 -34393
rect -96 -34433 96 -34427
rect -96 -34501 96 -34495
rect -96 -34535 -84 -34501
rect 84 -34535 96 -34501
rect -96 -34541 96 -34535
rect -152 -34594 -106 -34582
rect -152 -35770 -146 -34594
rect -112 -35770 -106 -34594
rect -152 -35782 -106 -35770
rect 106 -34594 152 -34582
rect 106 -35770 112 -34594
rect 146 -35770 152 -34594
rect 106 -35782 152 -35770
rect -96 -35829 96 -35823
rect -96 -35863 -84 -35829
rect 84 -35863 96 -35829
rect -96 -35869 96 -35863
rect -96 -35937 96 -35931
rect -96 -35971 -84 -35937
rect 84 -35971 96 -35937
rect -96 -35977 96 -35971
rect -152 -36030 -106 -36018
rect -152 -37206 -146 -36030
rect -112 -37206 -106 -36030
rect -152 -37218 -106 -37206
rect 106 -36030 152 -36018
rect 106 -37206 112 -36030
rect 146 -37206 152 -36030
rect 106 -37218 152 -37206
rect -96 -37265 96 -37259
rect -96 -37299 -84 -37265
rect 84 -37299 96 -37265
rect -96 -37305 96 -37299
rect -96 -37373 96 -37367
rect -96 -37407 -84 -37373
rect 84 -37407 96 -37373
rect -96 -37413 96 -37407
rect -152 -37466 -106 -37454
rect -152 -38642 -146 -37466
rect -112 -38642 -106 -37466
rect -152 -38654 -106 -38642
rect 106 -37466 152 -37454
rect 106 -38642 112 -37466
rect 146 -38642 152 -37466
rect 106 -38654 152 -38642
rect -96 -38701 96 -38695
rect -96 -38735 -84 -38701
rect 84 -38735 96 -38701
rect -96 -38741 96 -38735
rect -96 -38809 96 -38803
rect -96 -38843 -84 -38809
rect 84 -38843 96 -38809
rect -96 -38849 96 -38843
rect -152 -38902 -106 -38890
rect -152 -40078 -146 -38902
rect -112 -40078 -106 -38902
rect -152 -40090 -106 -40078
rect 106 -38902 152 -38890
rect 106 -40078 112 -38902
rect 146 -40078 152 -38902
rect 106 -40090 152 -40078
rect -96 -40137 96 -40131
rect -96 -40171 -84 -40137
rect 84 -40171 96 -40137
rect -96 -40177 96 -40171
rect -96 -40245 96 -40239
rect -96 -40279 -84 -40245
rect 84 -40279 96 -40245
rect -96 -40285 96 -40279
rect -152 -40338 -106 -40326
rect -152 -41514 -146 -40338
rect -112 -41514 -106 -40338
rect -152 -41526 -106 -41514
rect 106 -40338 152 -40326
rect 106 -41514 112 -40338
rect 146 -41514 152 -40338
rect 106 -41526 152 -41514
rect -96 -41573 96 -41567
rect -96 -41607 -84 -41573
rect 84 -41607 96 -41573
rect -96 -41613 96 -41607
rect -96 -41681 96 -41675
rect -96 -41715 -84 -41681
rect 84 -41715 96 -41681
rect -96 -41721 96 -41715
rect -152 -41774 -106 -41762
rect -152 -42950 -146 -41774
rect -112 -42950 -106 -41774
rect -152 -42962 -106 -42950
rect 106 -41774 152 -41762
rect 106 -42950 112 -41774
rect 146 -42950 152 -41774
rect 106 -42962 152 -42950
rect -96 -43009 96 -43003
rect -96 -43043 -84 -43009
rect 84 -43043 96 -43009
rect -96 -43049 96 -43043
rect -96 -43117 96 -43111
rect -96 -43151 -84 -43117
rect 84 -43151 96 -43117
rect -96 -43157 96 -43151
rect -152 -43210 -106 -43198
rect -152 -44386 -146 -43210
rect -112 -44386 -106 -43210
rect -152 -44398 -106 -44386
rect 106 -43210 152 -43198
rect 106 -44386 112 -43210
rect 146 -44386 152 -43210
rect 106 -44398 152 -44386
rect -96 -44445 96 -44439
rect -96 -44479 -84 -44445
rect 84 -44479 96 -44445
rect -96 -44485 96 -44479
rect -96 -44553 96 -44547
rect -96 -44587 -84 -44553
rect 84 -44587 96 -44553
rect -96 -44593 96 -44587
rect -152 -44646 -106 -44634
rect -152 -45822 -146 -44646
rect -112 -45822 -106 -44646
rect -152 -45834 -106 -45822
rect 106 -44646 152 -44634
rect 106 -45822 112 -44646
rect 146 -45822 152 -44646
rect 106 -45834 152 -45822
rect -96 -45881 96 -45875
rect -96 -45915 -84 -45881
rect 84 -45915 96 -45881
rect -96 -45921 96 -45915
rect -96 -45989 96 -45983
rect -96 -46023 -84 -45989
rect 84 -46023 96 -45989
rect -96 -46029 96 -46023
rect -152 -46082 -106 -46070
rect -152 -47258 -146 -46082
rect -112 -47258 -106 -46082
rect -152 -47270 -106 -47258
rect 106 -46082 152 -46070
rect 106 -47258 112 -46082
rect 146 -47258 152 -46082
rect 106 -47270 152 -47258
rect -96 -47317 96 -47311
rect -96 -47351 -84 -47317
rect 84 -47351 96 -47317
rect -96 -47357 96 -47351
rect -96 -47425 96 -47419
rect -96 -47459 -84 -47425
rect 84 -47459 96 -47425
rect -96 -47465 96 -47459
rect -152 -47518 -106 -47506
rect -152 -48694 -146 -47518
rect -112 -48694 -106 -47518
rect -152 -48706 -106 -48694
rect 106 -47518 152 -47506
rect 106 -48694 112 -47518
rect 146 -48694 152 -47518
rect 106 -48706 152 -48694
rect -96 -48753 96 -48747
rect -96 -48787 -84 -48753
rect 84 -48787 96 -48753
rect -96 -48793 96 -48787
rect -96 -48861 96 -48855
rect -96 -48895 -84 -48861
rect 84 -48895 96 -48861
rect -96 -48901 96 -48895
rect -152 -48954 -106 -48942
rect -152 -50130 -146 -48954
rect -112 -50130 -106 -48954
rect -152 -50142 -106 -50130
rect 106 -48954 152 -48942
rect 106 -50130 112 -48954
rect 146 -50130 152 -48954
rect 106 -50142 152 -50130
rect -96 -50189 96 -50183
rect -96 -50223 -84 -50189
rect 84 -50223 96 -50189
rect -96 -50229 96 -50223
rect -96 -50297 96 -50291
rect -96 -50331 -84 -50297
rect 84 -50331 96 -50297
rect -96 -50337 96 -50331
rect -152 -50390 -106 -50378
rect -152 -51566 -146 -50390
rect -112 -51566 -106 -50390
rect -152 -51578 -106 -51566
rect 106 -50390 152 -50378
rect 106 -51566 112 -50390
rect 146 -51566 152 -50390
rect 106 -51578 152 -51566
rect -96 -51625 96 -51619
rect -96 -51659 -84 -51625
rect 84 -51659 96 -51625
rect -96 -51665 96 -51659
rect -96 -51733 96 -51727
rect -96 -51767 -84 -51733
rect 84 -51767 96 -51733
rect -96 -51773 96 -51767
rect -152 -51826 -106 -51814
rect -152 -53002 -146 -51826
rect -112 -53002 -106 -51826
rect -152 -53014 -106 -53002
rect 106 -51826 152 -51814
rect 106 -53002 112 -51826
rect 146 -53002 152 -51826
rect 106 -53014 152 -53002
rect -96 -53061 96 -53055
rect -96 -53095 -84 -53061
rect 84 -53095 96 -53061
rect -96 -53101 96 -53095
rect -96 -53169 96 -53163
rect -96 -53203 -84 -53169
rect 84 -53203 96 -53169
rect -96 -53209 96 -53203
rect -152 -53262 -106 -53250
rect -152 -54438 -146 -53262
rect -112 -54438 -106 -53262
rect -152 -54450 -106 -54438
rect 106 -53262 152 -53250
rect 106 -54438 112 -53262
rect 146 -54438 152 -53262
rect 106 -54450 152 -54438
rect -96 -54497 96 -54491
rect -96 -54531 -84 -54497
rect 84 -54531 96 -54497
rect -96 -54537 96 -54531
rect -96 -54605 96 -54599
rect -96 -54639 -84 -54605
rect 84 -54639 96 -54605
rect -96 -54645 96 -54639
rect -152 -54698 -106 -54686
rect -152 -55874 -146 -54698
rect -112 -55874 -106 -54698
rect -152 -55886 -106 -55874
rect 106 -54698 152 -54686
rect 106 -55874 112 -54698
rect 146 -55874 152 -54698
rect 106 -55886 152 -55874
rect -96 -55933 96 -55927
rect -96 -55967 -84 -55933
rect 84 -55967 96 -55933
rect -96 -55973 96 -55967
rect -96 -56041 96 -56035
rect -96 -56075 -84 -56041
rect 84 -56075 96 -56041
rect -96 -56081 96 -56075
rect -152 -56134 -106 -56122
rect -152 -57310 -146 -56134
rect -112 -57310 -106 -56134
rect -152 -57322 -106 -57310
rect 106 -56134 152 -56122
rect 106 -57310 112 -56134
rect 146 -57310 152 -56134
rect 106 -57322 152 -57310
rect -96 -57369 96 -57363
rect -96 -57403 -84 -57369
rect 84 -57403 96 -57369
rect -96 -57409 96 -57403
rect -96 -57477 96 -57471
rect -96 -57511 -84 -57477
rect 84 -57511 96 -57477
rect -96 -57517 96 -57511
rect -152 -57570 -106 -57558
rect -152 -58746 -146 -57570
rect -112 -58746 -106 -57570
rect -152 -58758 -106 -58746
rect 106 -57570 152 -57558
rect 106 -58746 112 -57570
rect 146 -58746 152 -57570
rect 106 -58758 152 -58746
rect -96 -58805 96 -58799
rect -96 -58839 -84 -58805
rect 84 -58839 96 -58805
rect -96 -58845 96 -58839
rect -96 -58913 96 -58907
rect -96 -58947 -84 -58913
rect 84 -58947 96 -58913
rect -96 -58953 96 -58947
rect -152 -59006 -106 -58994
rect -152 -60182 -146 -59006
rect -112 -60182 -106 -59006
rect -152 -60194 -106 -60182
rect 106 -59006 152 -58994
rect 106 -60182 112 -59006
rect 146 -60182 152 -59006
rect 106 -60194 152 -60182
rect -96 -60241 96 -60235
rect -96 -60275 -84 -60241
rect 84 -60275 96 -60241
rect -96 -60281 96 -60275
rect -96 -60349 96 -60343
rect -96 -60383 -84 -60349
rect 84 -60383 96 -60349
rect -96 -60389 96 -60383
rect -152 -60442 -106 -60430
rect -152 -61618 -146 -60442
rect -112 -61618 -106 -60442
rect -152 -61630 -106 -61618
rect 106 -60442 152 -60430
rect 106 -61618 112 -60442
rect 146 -61618 152 -60442
rect 106 -61630 152 -61618
rect -96 -61677 96 -61671
rect -96 -61711 -84 -61677
rect 84 -61711 96 -61677
rect -96 -61717 96 -61711
rect -96 -61785 96 -61779
rect -96 -61819 -84 -61785
rect 84 -61819 96 -61785
rect -96 -61825 96 -61819
rect -152 -61878 -106 -61866
rect -152 -63054 -146 -61878
rect -112 -63054 -106 -61878
rect -152 -63066 -106 -63054
rect 106 -61878 152 -61866
rect 106 -63054 112 -61878
rect 146 -63054 152 -61878
rect 106 -63066 152 -63054
rect -96 -63113 96 -63107
rect -96 -63147 -84 -63113
rect 84 -63147 96 -63113
rect -96 -63153 96 -63147
rect -96 -63221 96 -63215
rect -96 -63255 -84 -63221
rect 84 -63255 96 -63221
rect -96 -63261 96 -63255
rect -152 -63314 -106 -63302
rect -152 -64490 -146 -63314
rect -112 -64490 -106 -63314
rect -152 -64502 -106 -64490
rect 106 -63314 152 -63302
rect 106 -64490 112 -63314
rect 146 -64490 152 -63314
rect 106 -64502 152 -64490
rect -96 -64549 96 -64543
rect -96 -64583 -84 -64549
rect 84 -64583 96 -64549
rect -96 -64589 96 -64583
rect -96 -64657 96 -64651
rect -96 -64691 -84 -64657
rect 84 -64691 96 -64657
rect -96 -64697 96 -64691
rect -152 -64750 -106 -64738
rect -152 -65926 -146 -64750
rect -112 -65926 -106 -64750
rect -152 -65938 -106 -65926
rect 106 -64750 152 -64738
rect 106 -65926 112 -64750
rect 146 -65926 152 -64750
rect 106 -65938 152 -65926
rect -96 -65985 96 -65979
rect -96 -66019 -84 -65985
rect 84 -66019 96 -65985
rect -96 -66025 96 -66019
rect -96 -66093 96 -66087
rect -96 -66127 -84 -66093
rect 84 -66127 96 -66093
rect -96 -66133 96 -66127
rect -152 -66186 -106 -66174
rect -152 -67362 -146 -66186
rect -112 -67362 -106 -66186
rect -152 -67374 -106 -67362
rect 106 -66186 152 -66174
rect 106 -67362 112 -66186
rect 146 -67362 152 -66186
rect 106 -67374 152 -67362
rect -96 -67421 96 -67415
rect -96 -67455 -84 -67421
rect 84 -67455 96 -67421
rect -96 -67461 96 -67455
rect -96 -67529 96 -67523
rect -96 -67563 -84 -67529
rect 84 -67563 96 -67529
rect -96 -67569 96 -67563
rect -152 -67622 -106 -67610
rect -152 -68798 -146 -67622
rect -112 -68798 -106 -67622
rect -152 -68810 -106 -68798
rect 106 -67622 152 -67610
rect 106 -68798 112 -67622
rect 146 -68798 152 -67622
rect 106 -68810 152 -68798
rect -96 -68857 96 -68851
rect -96 -68891 -84 -68857
rect 84 -68891 96 -68857
rect -96 -68897 96 -68891
rect -96 -68965 96 -68959
rect -96 -68999 -84 -68965
rect 84 -68999 96 -68965
rect -96 -69005 96 -68999
rect -152 -69058 -106 -69046
rect -152 -70234 -146 -69058
rect -112 -70234 -106 -69058
rect -152 -70246 -106 -70234
rect 106 -69058 152 -69046
rect 106 -70234 112 -69058
rect 146 -70234 152 -69058
rect 106 -70246 152 -70234
rect -96 -70293 96 -70287
rect -96 -70327 -84 -70293
rect 84 -70327 96 -70293
rect -96 -70333 96 -70327
rect -96 -70401 96 -70395
rect -96 -70435 -84 -70401
rect 84 -70435 96 -70401
rect -96 -70441 96 -70435
rect -152 -70494 -106 -70482
rect -152 -71670 -146 -70494
rect -112 -71670 -106 -70494
rect -152 -71682 -106 -71670
rect 106 -70494 152 -70482
rect 106 -71670 112 -70494
rect 146 -71670 152 -70494
rect 106 -71682 152 -71670
rect -96 -71729 96 -71723
rect -96 -71763 -84 -71729
rect 84 -71763 96 -71729
rect -96 -71769 96 -71763
rect -96 -71837 96 -71831
rect -96 -71871 -84 -71837
rect 84 -71871 96 -71837
rect -96 -71877 96 -71871
rect -152 -71930 -106 -71918
rect -152 -73106 -146 -71930
rect -112 -73106 -106 -71930
rect -152 -73118 -106 -73106
rect 106 -71930 152 -71918
rect 106 -73106 112 -71930
rect 146 -73106 152 -71930
rect 106 -73118 152 -73106
rect -96 -73165 96 -73159
rect -96 -73199 -84 -73165
rect 84 -73199 96 -73165
rect -96 -73205 96 -73199
rect -96 -73273 96 -73267
rect -96 -73307 -84 -73273
rect 84 -73307 96 -73273
rect -96 -73313 96 -73307
rect -152 -73366 -106 -73354
rect -152 -74542 -146 -73366
rect -112 -74542 -106 -73366
rect -152 -74554 -106 -74542
rect 106 -73366 152 -73354
rect 106 -74542 112 -73366
rect 146 -74542 152 -73366
rect 106 -74554 152 -74542
rect -96 -74601 96 -74595
rect -96 -74635 -84 -74601
rect 84 -74635 96 -74601
rect -96 -74641 96 -74635
rect -96 -74709 96 -74703
rect -96 -74743 -84 -74709
rect 84 -74743 96 -74709
rect -96 -74749 96 -74743
rect -152 -74802 -106 -74790
rect -152 -75978 -146 -74802
rect -112 -75978 -106 -74802
rect -152 -75990 -106 -75978
rect 106 -74802 152 -74790
rect 106 -75978 112 -74802
rect 146 -75978 152 -74802
rect 106 -75990 152 -75978
rect -96 -76037 96 -76031
rect -96 -76071 -84 -76037
rect 84 -76071 96 -76037
rect -96 -76077 96 -76071
rect -96 -76145 96 -76139
rect -96 -76179 -84 -76145
rect 84 -76179 96 -76145
rect -96 -76185 96 -76179
rect -152 -76238 -106 -76226
rect -152 -77414 -146 -76238
rect -112 -77414 -106 -76238
rect -152 -77426 -106 -77414
rect 106 -76238 152 -76226
rect 106 -77414 112 -76238
rect 146 -77414 152 -76238
rect 106 -77426 152 -77414
rect -96 -77473 96 -77467
rect -96 -77507 -84 -77473
rect 84 -77507 96 -77473
rect -96 -77513 96 -77507
rect -96 -77581 96 -77575
rect -96 -77615 -84 -77581
rect 84 -77615 96 -77581
rect -96 -77621 96 -77615
rect -152 -77674 -106 -77662
rect -152 -78850 -146 -77674
rect -112 -78850 -106 -77674
rect -152 -78862 -106 -78850
rect 106 -77674 152 -77662
rect 106 -78850 112 -77674
rect 146 -78850 152 -77674
rect 106 -78862 152 -78850
rect -96 -78909 96 -78903
rect -96 -78943 -84 -78909
rect 84 -78943 96 -78909
rect -96 -78949 96 -78943
rect -96 -79017 96 -79011
rect -96 -79051 -84 -79017
rect 84 -79051 96 -79017
rect -96 -79057 96 -79051
rect -152 -79110 -106 -79098
rect -152 -80286 -146 -79110
rect -112 -80286 -106 -79110
rect -152 -80298 -106 -80286
rect 106 -79110 152 -79098
rect 106 -80286 112 -79110
rect 146 -80286 152 -79110
rect 106 -80298 152 -80286
rect -96 -80345 96 -80339
rect -96 -80379 -84 -80345
rect 84 -80379 96 -80345
rect -96 -80385 96 -80379
rect -96 -80453 96 -80447
rect -96 -80487 -84 -80453
rect 84 -80487 96 -80453
rect -96 -80493 96 -80487
rect -152 -80546 -106 -80534
rect -152 -81722 -146 -80546
rect -112 -81722 -106 -80546
rect -152 -81734 -106 -81722
rect 106 -80546 152 -80534
rect 106 -81722 112 -80546
rect 146 -81722 152 -80546
rect 106 -81734 152 -81722
rect -96 -81781 96 -81775
rect -96 -81815 -84 -81781
rect 84 -81815 96 -81781
rect -96 -81821 96 -81815
rect -96 -81889 96 -81883
rect -96 -81923 -84 -81889
rect 84 -81923 96 -81889
rect -96 -81929 96 -81923
rect -152 -81982 -106 -81970
rect -152 -83158 -146 -81982
rect -112 -83158 -106 -81982
rect -152 -83170 -106 -83158
rect 106 -81982 152 -81970
rect 106 -83158 112 -81982
rect 146 -83158 152 -81982
rect 106 -83170 152 -83158
rect -96 -83217 96 -83211
rect -96 -83251 -84 -83217
rect 84 -83251 96 -83217
rect -96 -83257 96 -83251
rect -96 -83325 96 -83319
rect -96 -83359 -84 -83325
rect 84 -83359 96 -83325
rect -96 -83365 96 -83359
rect -152 -83418 -106 -83406
rect -152 -84594 -146 -83418
rect -112 -84594 -106 -83418
rect -152 -84606 -106 -84594
rect 106 -83418 152 -83406
rect 106 -84594 112 -83418
rect 146 -84594 152 -83418
rect 106 -84606 152 -84594
rect -96 -84653 96 -84647
rect -96 -84687 -84 -84653
rect 84 -84687 96 -84653
rect -96 -84693 96 -84687
rect -96 -84761 96 -84755
rect -96 -84795 -84 -84761
rect 84 -84795 96 -84761
rect -96 -84801 96 -84795
rect -152 -84854 -106 -84842
rect -152 -86030 -146 -84854
rect -112 -86030 -106 -84854
rect -152 -86042 -106 -86030
rect 106 -84854 152 -84842
rect 106 -86030 112 -84854
rect 146 -86030 152 -84854
rect 106 -86042 152 -86030
rect -96 -86089 96 -86083
rect -96 -86123 -84 -86089
rect 84 -86123 96 -86089
rect -96 -86129 96 -86123
rect -96 -86197 96 -86191
rect -96 -86231 -84 -86197
rect 84 -86231 96 -86197
rect -96 -86237 96 -86231
rect -152 -86290 -106 -86278
rect -152 -87466 -146 -86290
rect -112 -87466 -106 -86290
rect -152 -87478 -106 -87466
rect 106 -86290 152 -86278
rect 106 -87466 112 -86290
rect 146 -87466 152 -86290
rect 106 -87478 152 -87466
rect -96 -87525 96 -87519
rect -96 -87559 -84 -87525
rect 84 -87559 96 -87525
rect -96 -87565 96 -87559
rect -96 -87633 96 -87627
rect -96 -87667 -84 -87633
rect 84 -87667 96 -87633
rect -96 -87673 96 -87667
rect -152 -87726 -106 -87714
rect -152 -88902 -146 -87726
rect -112 -88902 -106 -87726
rect -152 -88914 -106 -88902
rect 106 -87726 152 -87714
rect 106 -88902 112 -87726
rect 146 -88902 152 -87726
rect 106 -88914 152 -88902
rect -96 -88961 96 -88955
rect -96 -88995 -84 -88961
rect 84 -88995 96 -88961
rect -96 -89001 96 -88995
rect -96 -89069 96 -89063
rect -96 -89103 -84 -89069
rect 84 -89103 96 -89069
rect -96 -89109 96 -89103
rect -152 -89162 -106 -89150
rect -152 -90338 -146 -89162
rect -112 -90338 -106 -89162
rect -152 -90350 -106 -90338
rect 106 -89162 152 -89150
rect 106 -90338 112 -89162
rect 146 -90338 152 -89162
rect 106 -90350 152 -90338
rect -96 -90397 96 -90391
rect -96 -90431 -84 -90397
rect 84 -90431 96 -90397
rect -96 -90437 96 -90431
rect -96 -90505 96 -90499
rect -96 -90539 -84 -90505
rect 84 -90539 96 -90505
rect -96 -90545 96 -90539
rect -152 -90598 -106 -90586
rect -152 -91774 -146 -90598
rect -112 -91774 -106 -90598
rect -152 -91786 -106 -91774
rect 106 -90598 152 -90586
rect 106 -91774 112 -90598
rect 146 -91774 152 -90598
rect 106 -91786 152 -91774
rect -96 -91833 96 -91827
rect -96 -91867 -84 -91833
rect 84 -91867 96 -91833
rect -96 -91873 96 -91867
rect -96 -91941 96 -91935
rect -96 -91975 -84 -91941
rect 84 -91975 96 -91941
rect -96 -91981 96 -91975
rect -152 -92034 -106 -92022
rect -152 -93210 -146 -92034
rect -112 -93210 -106 -92034
rect -152 -93222 -106 -93210
rect 106 -92034 152 -92022
rect 106 -93210 112 -92034
rect 146 -93210 152 -92034
rect 106 -93222 152 -93210
rect -96 -93269 96 -93263
rect -96 -93303 -84 -93269
rect 84 -93303 96 -93269
rect -96 -93309 96 -93303
rect -96 -93377 96 -93371
rect -96 -93411 -84 -93377
rect 84 -93411 96 -93377
rect -96 -93417 96 -93411
rect -152 -93470 -106 -93458
rect -152 -94646 -146 -93470
rect -112 -94646 -106 -93470
rect -152 -94658 -106 -94646
rect 106 -93470 152 -93458
rect 106 -94646 112 -93470
rect 146 -94646 152 -93470
rect 106 -94658 152 -94646
rect -96 -94705 96 -94699
rect -96 -94739 -84 -94705
rect 84 -94739 96 -94705
rect -96 -94745 96 -94739
rect -96 -94813 96 -94807
rect -96 -94847 -84 -94813
rect 84 -94847 96 -94813
rect -96 -94853 96 -94847
rect -152 -94906 -106 -94894
rect -152 -96082 -146 -94906
rect -112 -96082 -106 -94906
rect -152 -96094 -106 -96082
rect 106 -94906 152 -94894
rect 106 -96082 112 -94906
rect 146 -96082 152 -94906
rect 106 -96094 152 -96082
rect -96 -96141 96 -96135
rect -96 -96175 -84 -96141
rect 84 -96175 96 -96141
rect -96 -96181 96 -96175
rect -96 -96249 96 -96243
rect -96 -96283 -84 -96249
rect 84 -96283 96 -96249
rect -96 -96289 96 -96283
rect -152 -96342 -106 -96330
rect -152 -97518 -146 -96342
rect -112 -97518 -106 -96342
rect -152 -97530 -106 -97518
rect 106 -96342 152 -96330
rect 106 -97518 112 -96342
rect 146 -97518 152 -96342
rect 106 -97530 152 -97518
rect -96 -97577 96 -97571
rect -96 -97611 -84 -97577
rect 84 -97611 96 -97577
rect -96 -97617 96 -97611
rect -96 -97685 96 -97679
rect -96 -97719 -84 -97685
rect 84 -97719 96 -97685
rect -96 -97725 96 -97719
rect -152 -97778 -106 -97766
rect -152 -98954 -146 -97778
rect -112 -98954 -106 -97778
rect -152 -98966 -106 -98954
rect 106 -97778 152 -97766
rect 106 -98954 112 -97778
rect 146 -98954 152 -97778
rect 106 -98966 152 -98954
rect -96 -99013 96 -99007
rect -96 -99047 -84 -99013
rect 84 -99047 96 -99013
rect -96 -99053 96 -99047
rect -96 -99121 96 -99115
rect -96 -99155 -84 -99121
rect 84 -99155 96 -99121
rect -96 -99161 96 -99155
rect -152 -99214 -106 -99202
rect -152 -100390 -146 -99214
rect -112 -100390 -106 -99214
rect -152 -100402 -106 -100390
rect 106 -99214 152 -99202
rect 106 -100390 112 -99214
rect 146 -100390 152 -99214
rect 106 -100402 152 -100390
rect -96 -100449 96 -100443
rect -96 -100483 -84 -100449
rect 84 -100483 96 -100449
rect -96 -100489 96 -100483
rect -96 -100557 96 -100551
rect -96 -100591 -84 -100557
rect 84 -100591 96 -100557
rect -96 -100597 96 -100591
rect -152 -100650 -106 -100638
rect -152 -101826 -146 -100650
rect -112 -101826 -106 -100650
rect -152 -101838 -106 -101826
rect 106 -100650 152 -100638
rect 106 -101826 112 -100650
rect 146 -101826 152 -100650
rect 106 -101838 152 -101826
rect -96 -101885 96 -101879
rect -96 -101919 -84 -101885
rect 84 -101919 96 -101885
rect -96 -101925 96 -101919
rect -96 -101993 96 -101987
rect -96 -102027 -84 -101993
rect 84 -102027 96 -101993
rect -96 -102033 96 -102027
rect -152 -102086 -106 -102074
rect -152 -103262 -146 -102086
rect -112 -103262 -106 -102086
rect -152 -103274 -106 -103262
rect 106 -102086 152 -102074
rect 106 -103262 112 -102086
rect 146 -103262 152 -102086
rect 106 -103274 152 -103262
rect -96 -103321 96 -103315
rect -96 -103355 -84 -103321
rect 84 -103355 96 -103321
rect -96 -103361 96 -103355
rect -96 -103429 96 -103423
rect -96 -103463 -84 -103429
rect 84 -103463 96 -103429
rect -96 -103469 96 -103463
rect -152 -103522 -106 -103510
rect -152 -104698 -146 -103522
rect -112 -104698 -106 -103522
rect -152 -104710 -106 -104698
rect 106 -103522 152 -103510
rect 106 -104698 112 -103522
rect 146 -104698 152 -103522
rect 106 -104710 152 -104698
rect -96 -104757 96 -104751
rect -96 -104791 -84 -104757
rect 84 -104791 96 -104757
rect -96 -104797 96 -104791
rect -96 -104865 96 -104859
rect -96 -104899 -84 -104865
rect 84 -104899 96 -104865
rect -96 -104905 96 -104899
rect -152 -104958 -106 -104946
rect -152 -106134 -146 -104958
rect -112 -106134 -106 -104958
rect -152 -106146 -106 -106134
rect 106 -104958 152 -104946
rect 106 -106134 112 -104958
rect 146 -106134 152 -104958
rect 106 -106146 152 -106134
rect -96 -106193 96 -106187
rect -96 -106227 -84 -106193
rect 84 -106227 96 -106193
rect -96 -106233 96 -106227
rect -96 -106301 96 -106295
rect -96 -106335 -84 -106301
rect 84 -106335 96 -106301
rect -96 -106341 96 -106335
rect -152 -106394 -106 -106382
rect -152 -107570 -146 -106394
rect -112 -107570 -106 -106394
rect -152 -107582 -106 -107570
rect 106 -106394 152 -106382
rect 106 -107570 112 -106394
rect 146 -107570 152 -106394
rect 106 -107582 152 -107570
rect -96 -107629 96 -107623
rect -96 -107663 -84 -107629
rect 84 -107663 96 -107629
rect -96 -107669 96 -107663
rect -96 -107737 96 -107731
rect -96 -107771 -84 -107737
rect 84 -107771 96 -107737
rect -96 -107777 96 -107771
rect -152 -107830 -106 -107818
rect -152 -109006 -146 -107830
rect -112 -109006 -106 -107830
rect -152 -109018 -106 -109006
rect 106 -107830 152 -107818
rect 106 -109006 112 -107830
rect 146 -109006 152 -107830
rect 106 -109018 152 -109006
rect -96 -109065 96 -109059
rect -96 -109099 -84 -109065
rect 84 -109099 96 -109065
rect -96 -109105 96 -109099
rect -96 -109173 96 -109167
rect -96 -109207 -84 -109173
rect 84 -109207 96 -109173
rect -96 -109213 96 -109207
rect -152 -109266 -106 -109254
rect -152 -110442 -146 -109266
rect -112 -110442 -106 -109266
rect -152 -110454 -106 -110442
rect 106 -109266 152 -109254
rect 106 -110442 112 -109266
rect 146 -110442 152 -109266
rect 106 -110454 152 -110442
rect -96 -110501 96 -110495
rect -96 -110535 -84 -110501
rect 84 -110535 96 -110501
rect -96 -110541 96 -110535
rect -96 -110609 96 -110603
rect -96 -110643 -84 -110609
rect 84 -110643 96 -110609
rect -96 -110649 96 -110643
rect -152 -110702 -106 -110690
rect -152 -111878 -146 -110702
rect -112 -111878 -106 -110702
rect -152 -111890 -106 -111878
rect 106 -110702 152 -110690
rect 106 -111878 112 -110702
rect 146 -111878 152 -110702
rect 106 -111890 152 -111878
rect -96 -111937 96 -111931
rect -96 -111971 -84 -111937
rect 84 -111971 96 -111937
rect -96 -111977 96 -111971
rect -96 -112045 96 -112039
rect -96 -112079 -84 -112045
rect 84 -112079 96 -112045
rect -96 -112085 96 -112079
rect -152 -112138 -106 -112126
rect -152 -113314 -146 -112138
rect -112 -113314 -106 -112138
rect -152 -113326 -106 -113314
rect 106 -112138 152 -112126
rect 106 -113314 112 -112138
rect 146 -113314 152 -112138
rect 106 -113326 152 -113314
rect -96 -113373 96 -113367
rect -96 -113407 -84 -113373
rect 84 -113407 96 -113373
rect -96 -113413 96 -113407
rect -96 -113481 96 -113475
rect -96 -113515 -84 -113481
rect 84 -113515 96 -113481
rect -96 -113521 96 -113515
rect -152 -113574 -106 -113562
rect -152 -114750 -146 -113574
rect -112 -114750 -106 -113574
rect -152 -114762 -106 -114750
rect 106 -113574 152 -113562
rect 106 -114750 112 -113574
rect 146 -114750 152 -113574
rect 106 -114762 152 -114750
rect -96 -114809 96 -114803
rect -96 -114843 -84 -114809
rect 84 -114843 96 -114809
rect -96 -114849 96 -114843
rect -96 -114917 96 -114911
rect -96 -114951 -84 -114917
rect 84 -114951 96 -114917
rect -96 -114957 96 -114951
rect -152 -115010 -106 -114998
rect -152 -116186 -146 -115010
rect -112 -116186 -106 -115010
rect -152 -116198 -106 -116186
rect 106 -115010 152 -114998
rect 106 -116186 112 -115010
rect 146 -116186 152 -115010
rect 106 -116198 152 -116186
rect -96 -116245 96 -116239
rect -96 -116279 -84 -116245
rect 84 -116279 96 -116245
rect -96 -116285 96 -116279
rect -96 -116353 96 -116347
rect -96 -116387 -84 -116353
rect 84 -116387 96 -116353
rect -96 -116393 96 -116387
rect -152 -116446 -106 -116434
rect -152 -117622 -146 -116446
rect -112 -117622 -106 -116446
rect -152 -117634 -106 -117622
rect 106 -116446 152 -116434
rect 106 -117622 112 -116446
rect 146 -117622 152 -116446
rect 106 -117634 152 -117622
rect -96 -117681 96 -117675
rect -96 -117715 -84 -117681
rect 84 -117715 96 -117681
rect -96 -117721 96 -117715
rect -96 -117789 96 -117783
rect -96 -117823 -84 -117789
rect 84 -117823 96 -117789
rect -96 -117829 96 -117823
rect -152 -117882 -106 -117870
rect -152 -119058 -146 -117882
rect -112 -119058 -106 -117882
rect -152 -119070 -106 -119058
rect 106 -117882 152 -117870
rect 106 -119058 112 -117882
rect 146 -119058 152 -117882
rect 106 -119070 152 -119058
rect -96 -119117 96 -119111
rect -96 -119151 -84 -119117
rect 84 -119151 96 -119117
rect -96 -119157 96 -119151
rect -96 -119225 96 -119219
rect -96 -119259 -84 -119225
rect 84 -119259 96 -119225
rect -96 -119265 96 -119259
rect -152 -119318 -106 -119306
rect -152 -120494 -146 -119318
rect -112 -120494 -106 -119318
rect -152 -120506 -106 -120494
rect 106 -119318 152 -119306
rect 106 -120494 112 -119318
rect 146 -120494 152 -119318
rect 106 -120506 152 -120494
rect -96 -120553 96 -120547
rect -96 -120587 -84 -120553
rect 84 -120587 96 -120553
rect -96 -120593 96 -120587
rect -96 -120661 96 -120655
rect -96 -120695 -84 -120661
rect 84 -120695 96 -120661
rect -96 -120701 96 -120695
rect -152 -120754 -106 -120742
rect -152 -121930 -146 -120754
rect -112 -121930 -106 -120754
rect -152 -121942 -106 -121930
rect 106 -120754 152 -120742
rect 106 -121930 112 -120754
rect 146 -121930 152 -120754
rect 106 -121942 152 -121930
rect -96 -121989 96 -121983
rect -96 -122023 -84 -121989
rect 84 -122023 96 -121989
rect -96 -122029 96 -122023
rect -96 -122097 96 -122091
rect -96 -122131 -84 -122097
rect 84 -122131 96 -122097
rect -96 -122137 96 -122131
rect -152 -122190 -106 -122178
rect -152 -123366 -146 -122190
rect -112 -123366 -106 -122190
rect -152 -123378 -106 -123366
rect 106 -122190 152 -122178
rect 106 -123366 112 -122190
rect 146 -123366 152 -122190
rect 106 -123378 152 -123366
rect -96 -123425 96 -123419
rect -96 -123459 -84 -123425
rect 84 -123459 96 -123425
rect -96 -123465 96 -123459
rect -96 -123533 96 -123527
rect -96 -123567 -84 -123533
rect 84 -123567 96 -123533
rect -96 -123573 96 -123567
rect -152 -123626 -106 -123614
rect -152 -124802 -146 -123626
rect -112 -124802 -106 -123626
rect -152 -124814 -106 -124802
rect 106 -123626 152 -123614
rect 106 -124802 112 -123626
rect 146 -124802 152 -123626
rect 106 -124814 152 -124802
rect -96 -124861 96 -124855
rect -96 -124895 -84 -124861
rect 84 -124895 96 -124861
rect -96 -124901 96 -124895
rect -96 -124969 96 -124963
rect -96 -125003 -84 -124969
rect 84 -125003 96 -124969
rect -96 -125009 96 -125003
rect -152 -125062 -106 -125050
rect -152 -126238 -146 -125062
rect -112 -126238 -106 -125062
rect -152 -126250 -106 -126238
rect 106 -125062 152 -125050
rect 106 -126238 112 -125062
rect 146 -126238 152 -125062
rect 106 -126250 152 -126238
rect -96 -126297 96 -126291
rect -96 -126331 -84 -126297
rect 84 -126331 96 -126297
rect -96 -126337 96 -126331
rect -96 -126405 96 -126399
rect -96 -126439 -84 -126405
rect 84 -126439 96 -126405
rect -96 -126445 96 -126439
rect -152 -126498 -106 -126486
rect -152 -127674 -146 -126498
rect -112 -127674 -106 -126498
rect -152 -127686 -106 -127674
rect 106 -126498 152 -126486
rect 106 -127674 112 -126498
rect 146 -127674 152 -126498
rect 106 -127686 152 -127674
rect -96 -127733 96 -127727
rect -96 -127767 -84 -127733
rect 84 -127767 96 -127733
rect -96 -127773 96 -127767
rect -96 -127841 96 -127835
rect -96 -127875 -84 -127841
rect 84 -127875 96 -127841
rect -96 -127881 96 -127875
rect -152 -127934 -106 -127922
rect -152 -129110 -146 -127934
rect -112 -129110 -106 -127934
rect -152 -129122 -106 -129110
rect 106 -127934 152 -127922
rect 106 -129110 112 -127934
rect 146 -129110 152 -127934
rect 106 -129122 152 -129110
rect -96 -129169 96 -129163
rect -96 -129203 -84 -129169
rect 84 -129203 96 -129169
rect -96 -129209 96 -129203
rect -96 -129277 96 -129271
rect -96 -129311 -84 -129277
rect 84 -129311 96 -129277
rect -96 -129317 96 -129311
rect -152 -129370 -106 -129358
rect -152 -130546 -146 -129370
rect -112 -130546 -106 -129370
rect -152 -130558 -106 -130546
rect 106 -129370 152 -129358
rect 106 -130546 112 -129370
rect 146 -130546 152 -129370
rect 106 -130558 152 -130546
rect -96 -130605 96 -130599
rect -96 -130639 -84 -130605
rect 84 -130639 96 -130605
rect -96 -130645 96 -130639
rect -96 -130713 96 -130707
rect -96 -130747 -84 -130713
rect 84 -130747 96 -130713
rect -96 -130753 96 -130747
rect -152 -130806 -106 -130794
rect -152 -131982 -146 -130806
rect -112 -131982 -106 -130806
rect -152 -131994 -106 -131982
rect 106 -130806 152 -130794
rect 106 -131982 112 -130806
rect 146 -131982 152 -130806
rect 106 -131994 152 -131982
rect -96 -132041 96 -132035
rect -96 -132075 -84 -132041
rect 84 -132075 96 -132041
rect -96 -132081 96 -132075
rect -96 -132149 96 -132143
rect -96 -132183 -84 -132149
rect 84 -132183 96 -132149
rect -96 -132189 96 -132183
rect -152 -132242 -106 -132230
rect -152 -133418 -146 -132242
rect -112 -133418 -106 -132242
rect -152 -133430 -106 -133418
rect 106 -132242 152 -132230
rect 106 -133418 112 -132242
rect 146 -133418 152 -132242
rect 106 -133430 152 -133418
rect -96 -133477 96 -133471
rect -96 -133511 -84 -133477
rect 84 -133511 96 -133477
rect -96 -133517 96 -133511
rect -96 -133585 96 -133579
rect -96 -133619 -84 -133585
rect 84 -133619 96 -133585
rect -96 -133625 96 -133619
rect -152 -133678 -106 -133666
rect -152 -134854 -146 -133678
rect -112 -134854 -106 -133678
rect -152 -134866 -106 -134854
rect 106 -133678 152 -133666
rect 106 -134854 112 -133678
rect 146 -134854 152 -133678
rect 106 -134866 152 -134854
rect -96 -134913 96 -134907
rect -96 -134947 -84 -134913
rect 84 -134947 96 -134913
rect -96 -134953 96 -134947
rect -96 -135021 96 -135015
rect -96 -135055 -84 -135021
rect 84 -135055 96 -135021
rect -96 -135061 96 -135055
rect -152 -135114 -106 -135102
rect -152 -136290 -146 -135114
rect -112 -136290 -106 -135114
rect -152 -136302 -106 -136290
rect 106 -135114 152 -135102
rect 106 -136290 112 -135114
rect 146 -136290 152 -135114
rect 106 -136302 152 -136290
rect -96 -136349 96 -136343
rect -96 -136383 -84 -136349
rect 84 -136383 96 -136349
rect -96 -136389 96 -136383
rect -96 -136457 96 -136451
rect -96 -136491 -84 -136457
rect 84 -136491 96 -136457
rect -96 -136497 96 -136491
rect -152 -136550 -106 -136538
rect -152 -137726 -146 -136550
rect -112 -137726 -106 -136550
rect -152 -137738 -106 -137726
rect 106 -136550 152 -136538
rect 106 -137726 112 -136550
rect 146 -137726 152 -136550
rect 106 -137738 152 -137726
rect -96 -137785 96 -137779
rect -96 -137819 -84 -137785
rect 84 -137819 96 -137785
rect -96 -137825 96 -137819
rect -96 -137893 96 -137887
rect -96 -137927 -84 -137893
rect 84 -137927 96 -137893
rect -96 -137933 96 -137927
rect -152 -137986 -106 -137974
rect -152 -139162 -146 -137986
rect -112 -139162 -106 -137986
rect -152 -139174 -106 -139162
rect 106 -137986 152 -137974
rect 106 -139162 112 -137986
rect 146 -139162 152 -137986
rect 106 -139174 152 -139162
rect -96 -139221 96 -139215
rect -96 -139255 -84 -139221
rect 84 -139255 96 -139221
rect -96 -139261 96 -139255
rect -96 -139329 96 -139323
rect -96 -139363 -84 -139329
rect 84 -139363 96 -139329
rect -96 -139369 96 -139363
rect -152 -139422 -106 -139410
rect -152 -140598 -146 -139422
rect -112 -140598 -106 -139422
rect -152 -140610 -106 -140598
rect 106 -139422 152 -139410
rect 106 -140598 112 -139422
rect 146 -140598 152 -139422
rect 106 -140610 152 -140598
rect -96 -140657 96 -140651
rect -96 -140691 -84 -140657
rect 84 -140691 96 -140657
rect -96 -140697 96 -140691
rect -96 -140765 96 -140759
rect -96 -140799 -84 -140765
rect 84 -140799 96 -140765
rect -96 -140805 96 -140799
rect -152 -140858 -106 -140846
rect -152 -142034 -146 -140858
rect -112 -142034 -106 -140858
rect -152 -142046 -106 -142034
rect 106 -140858 152 -140846
rect 106 -142034 112 -140858
rect 146 -142034 152 -140858
rect 106 -142046 152 -142034
rect -96 -142093 96 -142087
rect -96 -142127 -84 -142093
rect 84 -142127 96 -142093
rect -96 -142133 96 -142127
rect -96 -142201 96 -142195
rect -96 -142235 -84 -142201
rect 84 -142235 96 -142201
rect -96 -142241 96 -142235
rect -152 -142294 -106 -142282
rect -152 -143470 -146 -142294
rect -112 -143470 -106 -142294
rect -152 -143482 -106 -143470
rect 106 -142294 152 -142282
rect 106 -143470 112 -142294
rect 146 -143470 152 -142294
rect 106 -143482 152 -143470
rect -96 -143529 96 -143523
rect -96 -143563 -84 -143529
rect 84 -143563 96 -143529
rect -96 -143569 96 -143563
rect -96 -143637 96 -143631
rect -96 -143671 -84 -143637
rect 84 -143671 96 -143637
rect -96 -143677 96 -143671
rect -152 -143730 -106 -143718
rect -152 -144906 -146 -143730
rect -112 -144906 -106 -143730
rect -152 -144918 -106 -144906
rect 106 -143730 152 -143718
rect 106 -144906 112 -143730
rect 146 -144906 152 -143730
rect 106 -144918 152 -144906
rect -96 -144965 96 -144959
rect -96 -144999 -84 -144965
rect 84 -144999 96 -144965
rect -96 -145005 96 -144999
rect -96 -145073 96 -145067
rect -96 -145107 -84 -145073
rect 84 -145107 96 -145073
rect -96 -145113 96 -145107
rect -152 -145166 -106 -145154
rect -152 -146342 -146 -145166
rect -112 -146342 -106 -145166
rect -152 -146354 -106 -146342
rect 106 -145166 152 -145154
rect 106 -146342 112 -145166
rect 146 -146342 152 -145166
rect 106 -146354 152 -146342
rect -96 -146401 96 -146395
rect -96 -146435 -84 -146401
rect 84 -146435 96 -146401
rect -96 -146441 96 -146435
rect -96 -146509 96 -146503
rect -96 -146543 -84 -146509
rect 84 -146543 96 -146509
rect -96 -146549 96 -146543
rect -152 -146602 -106 -146590
rect -152 -147778 -146 -146602
rect -112 -147778 -106 -146602
rect -152 -147790 -106 -147778
rect 106 -146602 152 -146590
rect 106 -147778 112 -146602
rect 146 -147778 152 -146602
rect 106 -147790 152 -147778
rect -96 -147837 96 -147831
rect -96 -147871 -84 -147837
rect 84 -147871 96 -147837
rect -96 -147877 96 -147871
rect -96 -147945 96 -147939
rect -96 -147979 -84 -147945
rect 84 -147979 96 -147945
rect -96 -147985 96 -147979
rect -152 -148038 -106 -148026
rect -152 -149214 -146 -148038
rect -112 -149214 -106 -148038
rect -152 -149226 -106 -149214
rect 106 -148038 152 -148026
rect 106 -149214 112 -148038
rect 146 -149214 152 -148038
rect 106 -149226 152 -149214
rect -96 -149273 96 -149267
rect -96 -149307 -84 -149273
rect 84 -149307 96 -149273
rect -96 -149313 96 -149307
rect -96 -149381 96 -149375
rect -96 -149415 -84 -149381
rect 84 -149415 96 -149381
rect -96 -149421 96 -149415
rect -152 -149474 -106 -149462
rect -152 -150650 -146 -149474
rect -112 -150650 -106 -149474
rect -152 -150662 -106 -150650
rect 106 -149474 152 -149462
rect 106 -150650 112 -149474
rect 146 -150650 152 -149474
rect 106 -150662 152 -150650
rect -96 -150709 96 -150703
rect -96 -150743 -84 -150709
rect 84 -150743 96 -150709
rect -96 -150749 96 -150743
rect -96 -150817 96 -150811
rect -96 -150851 -84 -150817
rect 84 -150851 96 -150817
rect -96 -150857 96 -150851
rect -152 -150910 -106 -150898
rect -152 -152086 -146 -150910
rect -112 -152086 -106 -150910
rect -152 -152098 -106 -152086
rect 106 -150910 152 -150898
rect 106 -152086 112 -150910
rect 146 -152086 152 -150910
rect 106 -152098 152 -152086
rect -96 -152145 96 -152139
rect -96 -152179 -84 -152145
rect 84 -152179 96 -152145
rect -96 -152185 96 -152179
rect -96 -152253 96 -152247
rect -96 -152287 -84 -152253
rect 84 -152287 96 -152253
rect -96 -152293 96 -152287
rect -152 -152346 -106 -152334
rect -152 -153522 -146 -152346
rect -112 -153522 -106 -152346
rect -152 -153534 -106 -153522
rect 106 -152346 152 -152334
rect 106 -153522 112 -152346
rect 146 -153522 152 -152346
rect 106 -153534 152 -153522
rect -96 -153581 96 -153575
rect -96 -153615 -84 -153581
rect 84 -153615 96 -153581
rect -96 -153621 96 -153615
rect -96 -153689 96 -153683
rect -96 -153723 -84 -153689
rect 84 -153723 96 -153689
rect -96 -153729 96 -153723
rect -152 -153782 -106 -153770
rect -152 -154958 -146 -153782
rect -112 -154958 -106 -153782
rect -152 -154970 -106 -154958
rect 106 -153782 152 -153770
rect 106 -154958 112 -153782
rect 146 -154958 152 -153782
rect 106 -154970 152 -154958
rect -96 -155017 96 -155011
rect -96 -155051 -84 -155017
rect 84 -155051 96 -155017
rect -96 -155057 96 -155051
rect -96 -155125 96 -155119
rect -96 -155159 -84 -155125
rect 84 -155159 96 -155125
rect -96 -155165 96 -155159
rect -152 -155218 -106 -155206
rect -152 -156394 -146 -155218
rect -112 -156394 -106 -155218
rect -152 -156406 -106 -156394
rect 106 -155218 152 -155206
rect 106 -156394 112 -155218
rect 146 -156394 152 -155218
rect 106 -156406 152 -156394
rect -96 -156453 96 -156447
rect -96 -156487 -84 -156453
rect 84 -156487 96 -156453
rect -96 -156493 96 -156487
rect -96 -156561 96 -156555
rect -96 -156595 -84 -156561
rect 84 -156595 96 -156561
rect -96 -156601 96 -156595
rect -152 -156654 -106 -156642
rect -152 -157830 -146 -156654
rect -112 -157830 -106 -156654
rect -152 -157842 -106 -157830
rect 106 -156654 152 -156642
rect 106 -157830 112 -156654
rect 146 -157830 152 -156654
rect 106 -157842 152 -157830
rect -96 -157889 96 -157883
rect -96 -157923 -84 -157889
rect 84 -157923 96 -157889
rect -96 -157929 96 -157923
rect -96 -157997 96 -157991
rect -96 -158031 -84 -157997
rect 84 -158031 96 -157997
rect -96 -158037 96 -158031
rect -152 -158090 -106 -158078
rect -152 -159266 -146 -158090
rect -112 -159266 -106 -158090
rect -152 -159278 -106 -159266
rect 106 -158090 152 -158078
rect 106 -159266 112 -158090
rect 146 -159266 152 -158090
rect 106 -159278 152 -159266
rect -96 -159325 96 -159319
rect -96 -159359 -84 -159325
rect 84 -159359 96 -159325
rect -96 -159365 96 -159359
rect -96 -159433 96 -159427
rect -96 -159467 -84 -159433
rect 84 -159467 96 -159433
rect -96 -159473 96 -159467
rect -152 -159526 -106 -159514
rect -152 -160702 -146 -159526
rect -112 -160702 -106 -159526
rect -152 -160714 -106 -160702
rect 106 -159526 152 -159514
rect 106 -160702 112 -159526
rect 146 -160702 152 -159526
rect 106 -160714 152 -160702
rect -96 -160761 96 -160755
rect -96 -160795 -84 -160761
rect 84 -160795 96 -160761
rect -96 -160801 96 -160795
rect -96 -160869 96 -160863
rect -96 -160903 -84 -160869
rect 84 -160903 96 -160869
rect -96 -160909 96 -160903
rect -152 -160962 -106 -160950
rect -152 -162138 -146 -160962
rect -112 -162138 -106 -160962
rect -152 -162150 -106 -162138
rect 106 -160962 152 -160950
rect 106 -162138 112 -160962
rect 146 -162138 152 -160962
rect 106 -162150 152 -162138
rect -96 -162197 96 -162191
rect -96 -162231 -84 -162197
rect 84 -162231 96 -162197
rect -96 -162237 96 -162231
rect -96 -162305 96 -162299
rect -96 -162339 -84 -162305
rect 84 -162339 96 -162305
rect -96 -162345 96 -162339
rect -152 -162398 -106 -162386
rect -152 -163574 -146 -162398
rect -112 -163574 -106 -162398
rect -152 -163586 -106 -163574
rect 106 -162398 152 -162386
rect 106 -163574 112 -162398
rect 146 -163574 152 -162398
rect 106 -163586 152 -163574
rect -96 -163633 96 -163627
rect -96 -163667 -84 -163633
rect 84 -163667 96 -163633
rect -96 -163673 96 -163667
rect -96 -163741 96 -163735
rect -96 -163775 -84 -163741
rect 84 -163775 96 -163741
rect -96 -163781 96 -163775
rect -152 -163834 -106 -163822
rect -152 -165010 -146 -163834
rect -112 -165010 -106 -163834
rect -152 -165022 -106 -165010
rect 106 -163834 152 -163822
rect 106 -165010 112 -163834
rect 146 -165010 152 -163834
rect 106 -165022 152 -165010
rect -96 -165069 96 -165063
rect -96 -165103 -84 -165069
rect 84 -165103 96 -165069
rect -96 -165109 96 -165103
rect -96 -165177 96 -165171
rect -96 -165211 -84 -165177
rect 84 -165211 96 -165177
rect -96 -165217 96 -165211
rect -152 -165270 -106 -165258
rect -152 -166446 -146 -165270
rect -112 -166446 -106 -165270
rect -152 -166458 -106 -166446
rect 106 -165270 152 -165258
rect 106 -166446 112 -165270
rect 146 -166446 152 -165270
rect 106 -166458 152 -166446
rect -96 -166505 96 -166499
rect -96 -166539 -84 -166505
rect 84 -166539 96 -166505
rect -96 -166545 96 -166539
rect -96 -166613 96 -166607
rect -96 -166647 -84 -166613
rect 84 -166647 96 -166613
rect -96 -166653 96 -166647
rect -152 -166706 -106 -166694
rect -152 -167882 -146 -166706
rect -112 -167882 -106 -166706
rect -152 -167894 -106 -167882
rect 106 -166706 152 -166694
rect 106 -167882 112 -166706
rect 146 -167882 152 -166706
rect 106 -167894 152 -167882
rect -96 -167941 96 -167935
rect -96 -167975 -84 -167941
rect 84 -167975 96 -167941
rect -96 -167981 96 -167975
rect -96 -168049 96 -168043
rect -96 -168083 -84 -168049
rect 84 -168083 96 -168049
rect -96 -168089 96 -168083
rect -152 -168142 -106 -168130
rect -152 -169318 -146 -168142
rect -112 -169318 -106 -168142
rect -152 -169330 -106 -169318
rect 106 -168142 152 -168130
rect 106 -169318 112 -168142
rect 146 -169318 152 -168142
rect 106 -169330 152 -169318
rect -96 -169377 96 -169371
rect -96 -169411 -84 -169377
rect 84 -169411 96 -169377
rect -96 -169417 96 -169411
rect -96 -169485 96 -169479
rect -96 -169519 -84 -169485
rect 84 -169519 96 -169485
rect -96 -169525 96 -169519
rect -152 -169578 -106 -169566
rect -152 -170754 -146 -169578
rect -112 -170754 -106 -169578
rect -152 -170766 -106 -170754
rect 106 -169578 152 -169566
rect 106 -170754 112 -169578
rect 146 -170754 152 -169578
rect 106 -170766 152 -170754
rect -96 -170813 96 -170807
rect -96 -170847 -84 -170813
rect 84 -170847 96 -170813
rect -96 -170853 96 -170847
rect -96 -170921 96 -170915
rect -96 -170955 -84 -170921
rect 84 -170955 96 -170921
rect -96 -170961 96 -170955
rect -152 -171014 -106 -171002
rect -152 -172190 -146 -171014
rect -112 -172190 -106 -171014
rect -152 -172202 -106 -172190
rect 106 -171014 152 -171002
rect 106 -172190 112 -171014
rect 146 -172190 152 -171014
rect 106 -172202 152 -172190
rect -96 -172249 96 -172243
rect -96 -172283 -84 -172249
rect 84 -172283 96 -172249
rect -96 -172289 96 -172283
rect -96 -172357 96 -172351
rect -96 -172391 -84 -172357
rect 84 -172391 96 -172357
rect -96 -172397 96 -172391
rect -152 -172450 -106 -172438
rect -152 -173626 -146 -172450
rect -112 -173626 -106 -172450
rect -152 -173638 -106 -173626
rect 106 -172450 152 -172438
rect 106 -173626 112 -172450
rect 146 -173626 152 -172450
rect 106 -173638 152 -173626
rect -96 -173685 96 -173679
rect -96 -173719 -84 -173685
rect 84 -173719 96 -173685
rect -96 -173725 96 -173719
rect -96 -173793 96 -173787
rect -96 -173827 -84 -173793
rect 84 -173827 96 -173793
rect -96 -173833 96 -173827
rect -152 -173886 -106 -173874
rect -152 -175062 -146 -173886
rect -112 -175062 -106 -173886
rect -152 -175074 -106 -175062
rect 106 -173886 152 -173874
rect 106 -175062 112 -173886
rect 146 -175062 152 -173886
rect 106 -175074 152 -175062
rect -96 -175121 96 -175115
rect -96 -175155 -84 -175121
rect 84 -175155 96 -175121
rect -96 -175161 96 -175155
rect -96 -175229 96 -175223
rect -96 -175263 -84 -175229
rect 84 -175263 96 -175229
rect -96 -175269 96 -175263
rect -152 -175322 -106 -175310
rect -152 -176498 -146 -175322
rect -112 -176498 -106 -175322
rect -152 -176510 -106 -176498
rect 106 -175322 152 -175310
rect 106 -176498 112 -175322
rect 146 -176498 152 -175322
rect 106 -176510 152 -176498
rect -96 -176557 96 -176551
rect -96 -176591 -84 -176557
rect 84 -176591 96 -176557
rect -96 -176597 96 -176591
rect -96 -176665 96 -176659
rect -96 -176699 -84 -176665
rect 84 -176699 96 -176665
rect -96 -176705 96 -176699
rect -152 -176758 -106 -176746
rect -152 -177934 -146 -176758
rect -112 -177934 -106 -176758
rect -152 -177946 -106 -177934
rect 106 -176758 152 -176746
rect 106 -177934 112 -176758
rect 146 -177934 152 -176758
rect 106 -177946 152 -177934
rect -96 -177993 96 -177987
rect -96 -178027 -84 -177993
rect 84 -178027 96 -177993
rect -96 -178033 96 -178027
rect -96 -178101 96 -178095
rect -96 -178135 -84 -178101
rect 84 -178135 96 -178101
rect -96 -178141 96 -178135
rect -152 -178194 -106 -178182
rect -152 -179370 -146 -178194
rect -112 -179370 -106 -178194
rect -152 -179382 -106 -179370
rect 106 -178194 152 -178182
rect 106 -179370 112 -178194
rect 146 -179370 152 -178194
rect 106 -179382 152 -179370
rect -96 -179429 96 -179423
rect -96 -179463 -84 -179429
rect 84 -179463 96 -179429
rect -96 -179469 96 -179463
rect -96 -179537 96 -179531
rect -96 -179571 -84 -179537
rect 84 -179571 96 -179537
rect -96 -179577 96 -179571
rect -152 -179630 -106 -179618
rect -152 -180806 -146 -179630
rect -112 -180806 -106 -179630
rect -152 -180818 -106 -180806
rect 106 -179630 152 -179618
rect 106 -180806 112 -179630
rect 146 -180806 152 -179630
rect 106 -180818 152 -180806
rect -96 -180865 96 -180859
rect -96 -180899 -84 -180865
rect 84 -180899 96 -180865
rect -96 -180905 96 -180899
rect -96 -180973 96 -180967
rect -96 -181007 -84 -180973
rect 84 -181007 96 -180973
rect -96 -181013 96 -181007
rect -152 -181066 -106 -181054
rect -152 -182242 -146 -181066
rect -112 -182242 -106 -181066
rect -152 -182254 -106 -182242
rect 106 -181066 152 -181054
rect 106 -182242 112 -181066
rect 146 -182242 152 -181066
rect 106 -182254 152 -182242
rect -96 -182301 96 -182295
rect -96 -182335 -84 -182301
rect 84 -182335 96 -182301
rect -96 -182341 96 -182335
rect -96 -182409 96 -182403
rect -96 -182443 -84 -182409
rect 84 -182443 96 -182409
rect -96 -182449 96 -182443
rect -152 -182502 -106 -182490
rect -152 -183678 -146 -182502
rect -112 -183678 -106 -182502
rect -152 -183690 -106 -183678
rect 106 -182502 152 -182490
rect 106 -183678 112 -182502
rect 146 -183678 152 -182502
rect 106 -183690 152 -183678
rect -96 -183737 96 -183731
rect -96 -183771 -84 -183737
rect 84 -183771 96 -183737
rect -96 -183777 96 -183771
<< properties >>
string FIXED_BBOX -263 -183892 263 183892
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 6.0 l 1.0 m 256 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
