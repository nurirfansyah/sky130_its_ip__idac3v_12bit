* NGSPICE file created from pcell256scs.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_BK8KVU a_n158_n84606# a_n158_60430# a_n100_n31571#
+ a_n100_n45931# a_n158_n111890# a_n100_38793# a_n158_n15678# a_n158_n71682# a_n158_n136302#
+ a_100_4426# a_n100_76129# a_n100_n106243# a_n100_n14339# a_n158_n27166# a_n100_n70343#
+ a_n158_n83170# a_n158_158078# a_n100_n84703# a_n158_n97530# a_n100_n133527# a_n158_17350#
+ a_100_5862# a_100_123614# a_n158_n150662# a_n100_77565# a_n100_123517# a_n158_30274#
+ a_n158_44634# a_n100_n15775# a_n100_90489# a_100_86278# a_n100_n134963# a_100_110690#
+ a_n158_71918# a_n100_110593# a_n158_n55886# a_n100_124953# a_n100_n145015# a_100_135102#
+ a_n158_n106146# a_n100_89053# a_n100_135005# a_n158_n176510# a_n158_n162150# a_n158_n1318#
+ a_n158_56122# a_n100_n27263# a_n100_n132091# a_n100_n146451# a_n158_n107582# a_n100_122081#
+ a_n100_n40187# a_n158_83406# a_n100_136441# a_n158_n2754# a_n100_n54547# a_n158_n67374#
+ a_n100_n68907# a_100_107818# a_100_n32910# a_n100_n173735# a_100_163822# a_n158_n134866#
+ a_n100_163725# a_n158_n80298# a_n158_n94658# a_n158_14478# a_n158_28838# a_n158_70482#
+ a_n158_84842# a_n100_n55983# a_n158_n119070# a_n100_n66035# a_n100_n129219# a_100_119306#
+ a_n158_n146354# a_n100_119209# a_100_175310# a_100_n120506# a_n100_175213# a_n100_n93319#
+ a_n100_n67471# a_n158_96330# a_n100_n116295# a_n158_n173638# a_100_106382# a_n100_106285#
+ a_n158_n147790# a_n100_n80395# a_n100_n94755# a_100_n121942# a_n100_n157939# a_n100_n143579#
+ a_100_133666# a_n100_133569# a_n100_147929# a_n158_54686# a_100_11606# a_100_n133430#
+ a_100_n14242# a_n100_n155067# a_100_n28602# a_n158_n116198# a_n100_n169427# a_100_145154#
+ a_100_159514# a_n100_145057# a_n100_159417# a_100_n160714# a_100_n41526# a_n158_66174#
+ a_100_172438# a_100_146590# a_n158_93458# a_n100_146493# a_n100_n64599# a_n158_123614#
+ a_n100_n78959# a_n100_n183787# a_100_n42962# a_100_10170# a_100_24530# a_100_173874#
+ a_100_n172202# a_n100_173777# a_100_n53014# a_n158_94894# a_n158_110690# a_100_51814#
+ a_n100_n76087# a_100_n103274# a_n158_135102# a_100_n117634# a_100_n40090# a_100_129358#
+ a_100_n54450# a_100_n68810# a_100_n130558# a_100_n144918# a_n100_11509# a_100_n81734#
+ a_100_63302# a_100_n129122# a_n158_107818# a_n158_n32910# a_100_n131994# a_n158_163822#
+ a_n100_12945# a_100_n142046# a_100_n156406# a_100_n37218# a_100_n93222# a_100_21658#
+ a_n100_7201# a_n158_119306# a_n158_n8498# a_n158_175310# a_100_n157842# a_100_n143482#
+ a_100_n24294# a_100_n38654# a_n100_n179479# a_n100_10073# a_n100_24433# a_100_169566#
+ a_n100_169469# a_100_n170766# a_100_n51578# a_n158_106382# a_100_n65938# a_100_33146#
+ a_n100_51717# a_100_47506# a_n158_4426# a_100_n169330# a_n158_133666# a_n100_n4287#
+ a_100_34582# a_100_48942# a_100_n182254# a_n158_5862# a_100_n63066# a_100_n77426#
+ a_n100_63205# a_100_61866# a_n158_n14242# a_n158_145154# a_n158_n28602# a_100_n127686#
+ a_n158_159514# a_n100_n120603# a_100_n183690# a_100_n5626# a_n100_4329# a_n100_50281#
+ a_100_n78862# a_100_46070# a_n100_64641# a_n158_n41526# a_n158_172438# a_n158_31710#
+ a_100_n91786# a_n100_91925# a_n158_146590# a_100_73354# a_100_87714# a_100_n139174#
+ a_n100_5765# a_n158_n42962# a_n158_173874# a_n100_22997# a_n158_n53014# a_100_18786#
+ a_100_n166458# a_100_n152098# a_100_74790# a_n100_33049# a_n158_n120506# a_n100_47409#
+ a_100_n4190# a_100_99202# a_n158_n40090# a_n100_n41623# a_n158_129358# a_n158_n54450#
+ a_n158_n68810# a_n100_n104807# a_100_n167894# a_n100_n160811# a_n100_34485# a_n100_48845#
+ a_n158_n121942# a_n100_150801# a_n158_n81734# a_n158_118# a_n158_15914# a_n100_61769#
+ a_100_43198# a_100_57558# a_n100_21# a_n100_n53111# a_100_n179382# a_n158_n133430#
+ a_n158_n37218# a_n158_n93222# a_n158_13042# a_100_58994# a_100_1554# a_n158_27402#
+ a_100_n87478# a_n100_73257# a_n100_87617# a_n100_n103371# a_n158_n160714# a_100_69046#
+ a_n100_n117731# a_n100_n11467# a_n158_40326# a_n100_107721# a_n158_n24294# a_n100_n25827#
+ a_n158_n38654# a_n158_169566# a_n100_n81831# a_n100_n130655# a_100_2990# a_n100_18689#
+ a_100_120742# a_n100_74693# a_n100_120645# a_n158_n51578# a_n158_n65938# a_n158_41762#
+ a_n158_n172202# a_n100_99105# a_100_97766# a_n100_n37315# a_n100_n142143# a_n158_n103274#
+ a_n100_n156503# a_100_132230# a_n100_n50239# a_n158_n117634# a_n100_86181# a_n100_132133#
+ a_n158_n63066# a_n158_n77426# a_n100_n24391# a_n158_53250# a_n158_67610# a_n100_n38751#
+ a_n158_n130558# a_n158_n144918# a_n158_80534# a_n100_n51675# a_n158_n78862# a_n100_n100499#
+ a_n100_n114859# a_n158_n129122# a_n100_n170863# a_100_104946# a_n158_n131994# a_n100_58897#
+ a_n100_104849# a_100_160950# a_n100_160853# a_n158_n91786# a_n158_n142046# a_n158_25966#
+ a_100_171002# a_n158_n156406# a_n158_81970# w_n358_n183987# a_n158_36018# a_n100_n63163#
+ a_100_n104710# a_n158_92022# a_n100_n77523# a_n100_n126347# a_100_102074# a_100_116434#
+ a_n100_n182351# a_n100_116337# a_n158_n157842# a_n158_n143482# a_n100_172341# a_n100_n90447#
+ a_100_n12806# a_n158_23094# a_n158_37454# a_100_143718# a_n158_n170766# a_100_79098#
+ a_n100_97669# a_n100_n127783# a_n158_50378# a_100_117870# a_n100_n35879# a_n100_n89011#
+ a_n158_64738# a_n100_117773# a_n100_n91883# a_n158_38890# a_100_130794# a_n158_n169330#
+ a_n100_130697# a_n100_n165119# a_100_155206# a_n100_155109# a_n158_n182254# a_n100_n139271#
+ a_n158_76226# a_n100_129261# a_n100_n47367# a_n158_n9934# a_100_n11370# a_100_n25730#
+ a_n100_n166555# a_n100_n152195# a_100_142282# a_n158_n127686# a_n100_142185# a_100_156642#
+ a_100_n101838# a_n158_n183690# a_n100_156545# a_n158_n87478# a_100_20222# a_n158_77662#
+ a_n100_n167991# a_n158_n7062# a_n158_90586# a_n158_120742# a_n100_157981# a_n100_n178043#
+ a_100_114998# a_100_168130# a_100_n113326# a_n158_n139174# a_n100_168033# a_n100_n5723#
+ a_n100_n86139# a_100_7298# a_100_n50142# a_100_n64502# a_n158_89150# a_100_181054#
+ a_n158_n166458# a_n158_n152098# a_n158_132230# a_n100_n87575# a_100_n114762# a_n100_n136399#
+ a_100_126486# a_n100_126389# a_100_182490# a_n158_n167894# a_n100_182393# a_100_n22858#
+ a_100_60430# a_100_n126250# a_n158_104946# a_n100_n99063# a_n158_160950# a_n158_n179382#
+ a_n158_171002# a_100_n153534# a_100_n34346# a_n100_20125# a_100_n48706# a_100_n90350#
+ a_100_165258# a_100_179618# a_100_n180818# a_n158_102074# a_n158_86278# a_n158_116434#
+ a_100_n154970# a_100_n35782# a_100_n109018# a_n100_21561# a_n100_35921# a_100_166694#
+ a_n158_n12806# a_100_n165022# a_100_17350# a_n158_143718# a_n100_166597# a_n158_117870#
+ a_100_30274# a_100_44634# a_n158_1554# a_100_n73118# a_n158_130794# a_100_n47270#
+ a_100_71918# a_100_178182# a_100_n123378# a_100_n137738# a_n158_155206# a_n100_178085#
+ a_100_n1318# a_100_n60194# a_n158_2990# a_100_n74554# a_100_n88914# a_n100_60333#
+ a_100_56122# a_n158_n11370# a_n100_n12903# a_n158_n25730# a_n158_142282# a_n158_156642#
+ a_100_83406# a_100_n2754# a_100_n19986# a_100_n75990# a_n100_1457# a_100_n149226#
+ a_100_n86042# a_100_14478# a_100_28838# a_100_70482# a_100_84842# a_n100_n10031#
+ a_n100_2893# a_n158_114998# a_n158_168130# a_n100_17253# a_n158_n104710# a_n158_n50142#
+ a_n158_n64502# a_100_n163586# a_n158_181054# a_100_n177946# a_100_n44398# a_100_n58758#
+ a_n100_30177# a_n100_44537# a_100_96330# a_n158_11606# a_n158_126486# a_n158_182490#
+ a_n100_n101935# a_n100_45973# a_n158_n22858# a_100_n175074# a_n100_56025# a_100_54686#
+ a_n100_83309# a_n100_n113423# a_100_103510# a_n100_57461# a_n100_103413# a_n100_n21519#
+ a_n158_n34346# a_n158_n48706# a_n158_165258# a_n158_n90350# a_n158_179618# a_n100_n140707#
+ a_n158_10170# a_n158_24530# a_n158_n101838# a_n100_70385# a_100_n98966# a_100_66174#
+ a_n100_84745# a_n100_n22955# a_n158_51814# a_n158_n35782# a_n158_166694# a_100_93458#
+ a_n100_n33007# a_100_n159278# a_100_n96094# a_n158_n113326# a_n100_96233# a_n158_n73118#
+ a_100_94894# a_n100_n20083# a_n158_63302# a_n100_n34443# a_n158_n47270# a_n100_n48803#
+ a_n158_178182# a_n100_n153631# a_n158_n114762# a_n158_n60194# a_n100_n61727# a_n158_n74554#
+ a_n100_143621# a_n158_n88914# a_100_100638# a_n100_n180915# a_n100_54589# a_n100_68949#
+ a_n100_170905# a_n158_7298# a_n158_21658# a_n158_n19986# a_n100_n109115# a_n158_n75990#
+ a_n100_n111987# a_n158_n126250# a_100_n100402# a_n100_101977# a_n100_n73215# a_n158_n86042#
+ a_n100_n122039# a_100_8734# a_100_112126# a_n100_66077# a_n100_112029# a_n158_n153534#
+ a_n158_33146# a_n100_n18647# a_n158_47506# a_n100_n60291# a_n100_n74651# a_n100_n123475#
+ a_n158_n180818# a_100_113562# a_100_n8498# a_n100_n137835# a_100_127922# a_n158_n44398#
+ a_n100_113465# a_n100_127825# a_n158_n58758# a_n158_n154970# a_n158_n109018# a_n158_n165022#
+ a_n100_n150759# a_n158_34582# a_n158_48942# a_100_140846# a_n100_94797# a_n100_140749#
+ a_n158_61866# a_n100_n149323# a_100_125050# a_100_139410# a_n100_n43059# a_n100_n57419#
+ a_n100_139313# a_n158_n5626# a_100_n140610# a_100_n21422# a_n100_n162247# a_n158_46070#
+ a_100_152334# a_n158_n123378# a_n158_n137738# a_n100_n176607# a_n100_152237# a_n100_n44495#
+ a_n158_73354# a_n158_87714# a_n158_103510# a_n100_n58855# a_n100_n107679# a_n100_n163683#
+ a_100_153770# a_n100_153673# a_n100_n71779# a_n158_n98966# a_n158_18786# a_n158_n149226#
+ a_n158_74790# a_n100_n1415# a_100_31710# a_n100_180957# a_n158_99202# a_n158_n4190#
+ a_n100_n119167# a_100_109254# a_n100_n175171# a_n100_109157# a_n100_n2851# a_n100_n83267#
+ a_n158_n96094# a_100_n110454# a_100_n124814# a_n100_165161# a_n100_179521# a_n100_n97627#
+ a_100_122178# a_100_136538# a_100_n61630# a_n158_n163586# a_n158_n177946# a_n158_43198#
+ a_n158_57558# a_n100_n28699# a_100_n111890# a_n100_n147887# a_100_137974# a_n158_100638#
+ a_100_n136302# a_n100_137877# a_100_n17114# a_100_148026# a_100_150898# a_n158_n175074#
+ a_100_15914# a_n158_58994# a_100_n30038# a_n158_69046# a_n100_n96191# a_n100_n159375#
+ a_100_n18550# a_100_149462# a_n158_112126# a_n100_149365# a_100_n150662# a_n100_n172299#
+ a_100_n31474# a_100_n45834# a_100_13042# a_n100_31613# a_100_162386# a_100_176746#
+ a_100_27402# a_n100_162289# a_n100_176649# a_n158_113562# a_100_40326# a_n158_97766#
+ a_n158_127922# a_100_n106146# a_100_118# a_100_n176510# a_100_n162150# a_n158_140846#
+ a_n100_43101# a_100_n57322# a_n158_n159278# a_100_41762# a_100_n70246# a_100_n84606#
+ a_100_n107582# a_n158_125050# a_n158_139410# a_n158_n21422# a_n158_152334# a_100_n134866#
+ a_100_n15678# a_n100_15817# a_100_n71682# a_n100_71821# a_100_53250# a_100_67610#
+ a_100_n119070# a_100_80534# a_n158_153770# a_100_n146354# a_100_n27166# a_n158_n100402#
+ a_n100_27305# a_100_158078# a_100_n83170# a_100_n97530# a_100_25966# a_100_n173638#
+ a_100_81970# a_n100_40229# a_n158_79098# a_n158_109254# a_100_36018# a_100_n147790#
+ a_100_92022# a_n100_14381# a_n100_28741# a_n158_122178# a_n158_n61630# a_n158_136538#
+ a_n100_41665# a_n100_n7159# a_100_n55886# a_100_23094# a_100_37454# a_n158_8734#
+ a_100_50378# a_n158_137974# a_100_64738# a_n158_n17114# a_100_n116198# a_n158_148026#
+ a_n100_n8595# a_100_38890# a_n158_150898# a_100_n67374# a_n100_53153# a_n100_67513#
+ a_n158_n30038# a_n158_n140610# a_n158_20222# a_n158_n18550# a_100_n80298# a_n100_80437#
+ a_100_n94658# a_100_76226# a_n158_149462# a_n100_n110551# a_n100_n124911# a_100_n9934#
+ a_n100_8637# a_n158_n31474# a_n100_100541# a_n100_114901# a_n158_n45834# a_n158_162386#
+ a_n158_176746# a_n100_25869# a_n100_79001# a_n100_81873# a_100_77662# a_n100_n17211#
+ a_100_n7062# a_100_90586# VSUBS a_n100_n30135# a_n158_n57322# a_n100_37357# a_n158_n110454#
+ a_n158_n124814# a_n100_93361# a_n158_n70246# a_100_89150#
X0 a_100_169566# a_n100_169469# a_n158_169566# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X1 a_100_53250# a_n100_53153# a_n158_53250# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X2 a_100_n98966# a_n100_n99063# a_n158_n98966# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X3 a_100_90586# a_n100_90489# a_n158_90586# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X4 a_100_21658# a_n100_21561# a_n158_21658# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X5 a_100_67610# a_n100_67513# a_n158_67610# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X6 a_100_123614# a_n100_123517# a_n158_123614# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X7 a_100_n11370# a_n100_n11467# a_n158_n11370# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X8 a_100_n152098# a_n100_n152195# a_n158_n152098# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X9 a_100_n110454# a_n100_n110551# a_n158_n110454# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X10 a_100_n80298# a_n100_n80395# a_n158_n80298# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X11 a_100_165258# a_n100_165161# a_n158_165258# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X12 a_100_n57322# a_n100_n57419# a_n158_n57322# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X13 a_100_153770# a_n100_153673# a_n158_153770# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X14 a_100_n129122# a_n100_n129219# a_n158_n129122# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X15 a_100_n124814# a_n100_n124911# a_n158_n124814# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X16 a_100_n94658# a_n100_n94755# a_n158_n94658# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X17 a_100_179618# a_n100_179521# a_n158_179618# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X18 a_100_n25730# a_n100_n25827# a_n158_n25730# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X19 a_100_n166458# a_n100_n166555# a_n158_n166458# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X20 a_100_126486# a_n100_126389# a_n158_126486# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X21 a_100_63302# a_n100_63205# a_n158_63302# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X22 a_100_n7062# a_n100_n7159# a_n158_n7062# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X23 a_100_10170# a_n100_10073# a_n158_10170# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X24 a_100_n2754# a_n100_n2851# a_n158_n2754# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X25 a_100_36018# a_n100_35921# a_n158_36018# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X26 a_100_n55886# a_n100_n55983# a_n158_n55886# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X27 a_100_n127686# a_n100_n127783# a_n158_n127686# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X28 a_100_n53014# a_n100_n53111# a_n158_n53014# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X29 a_100_n120506# a_n100_n120603# a_n158_n120506# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X30 a_100_n90350# a_n100_n90447# a_n158_n90350# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X31 a_100_24530# a_n100_24433# a_n158_24530# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X32 a_100_n162150# a_n100_n162247# a_n158_n162150# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X33 a_100_122178# a_n100_122081# a_n158_122178# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X34 a_100_66174# a_n100_66077# a_n158_66174# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X35 a_100_61866# a_n100_61769# a_n158_61866# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X36 a_100_168130# a_n100_168033# a_n158_168130# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X37 a_100_n14242# a_n100_n14339# a_n158_n14242# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X38 a_100_163822# a_n100_163725# a_n158_163822# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X39 a_100_110690# a_n100_110593# a_n158_110690# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X40 a_100_n150662# a_n100_n150759# a_n158_n150662# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X41 a_100_n176510# a_n100_n176607# a_n158_n176510# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X42 a_100_n51578# a_n100_n51675# a_n158_n51578# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X43 a_100_136538# a_n100_136441# a_n158_136538# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X44 a_100_n123378# a_n100_n123475# a_n158_n123378# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X45 a_100_118# a_n100_21# a_n158_118# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X46 a_100_n28602# a_n100_n28699# a_n158_n28602# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X47 a_100_20222# a_n100_20125# a_n158_20222# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X48 a_100_n65938# a_n100_n66035# a_n158_n65938# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X49 a_100_166694# a_n100_166597# a_n158_166694# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X50 a_100_n137738# a_n100_n137835# a_n158_n137738# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X51 a_100_76226# a_n100_76129# a_n158_76226# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X52 a_100_71918# a_n100_71821# a_n158_71918# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X53 a_100_23094# a_n100_22997# a_n158_23094# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X54 a_100_n167894# a_n100_n167991# a_n158_n167894# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X55 a_100_n93222# a_n100_n93319# a_n158_n93222# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X56 a_100_n165022# a_n100_n165119# a_n158_n165022# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X57 a_100_n160714# a_n100_n160811# a_n158_n160714# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X58 a_100_125050# a_n100_124953# a_n158_125050# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X59 a_100_120742# a_n100_120645# a_n158_120742# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X60 a_100_n61630# a_n100_n61727# a_n158_n61630# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X61 a_100_162386# a_n100_162289# a_n158_162386# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X62 a_100_n133430# a_n100_n133527# a_n158_n133430# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X63 a_100_37454# a_n100_37357# a_n158_37454# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X64 a_100_139410# a_n100_139313# a_n158_139410# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X65 a_100_79098# a_n100_79001# a_n158_79098# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X66 a_100_n96094# a_n100_n96191# a_n158_n96094# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X67 a_100_n27166# a_n100_n27263# a_n158_n27166# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X68 a_100_n121942# a_n100_n122039# a_n158_n121942# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X69 a_100_n91786# a_n100_n91883# a_n158_n91786# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X70 a_100_176746# a_n100_176649# a_n158_176746# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X71 a_100_n22858# a_n100_n22955# a_n158_n22858# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X72 a_100_n163586# a_n100_n163683# a_n158_n163586# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X73 a_100_107818# a_n100_107721# a_n158_107818# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X74 a_100_60430# a_n100_60333# a_n158_60430# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X75 a_100_n177946# a_n100_n178043# a_n158_n177946# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X76 a_100_137974# a_n100_137877# a_n158_137974# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X77 a_100_33146# a_n100_33049# a_n158_33146# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X78 a_100_n50142# a_n100_n50239# a_n158_n50142# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X79 a_100_135102# a_n100_135005# a_n158_135102# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X80 a_100_172438# a_n100_172341# a_n158_172438# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X81 a_100_47506# a_n100_47409# a_n158_47506# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X82 a_100_8734# a_n100_8637# a_n158_8734# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X83 a_100_n64502# a_n100_n64599# a_n158_n64502# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X84 a_100_160950# a_n100_160853# a_n158_160950# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X85 a_100_n136302# a_n100_n136399# a_n158_n136302# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X86 a_100_n32910# a_n100_n33007# a_n158_n32910# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X87 a_100_n37218# a_n100_n37315# a_n158_n37218# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X88 a_100_n173638# a_n100_n173735# a_n158_n173638# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X89 a_100_133666# a_n100_133569# a_n158_133666# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X90 a_100_77662# a_n100_77565# a_n158_77662# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X91 a_100_n109018# a_n100_n109115# a_n158_n109018# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X92 a_100_n104710# a_n100_n104807# a_n158_n104710# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X93 a_100_n67374# a_n100_n67471# a_n158_n67374# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X94 a_100_n139174# a_n100_n139271# a_n158_n139174# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X95 a_100_38890# a_n100_38793# a_n158_38890# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X96 a_100_4426# a_n100_4329# a_n158_4426# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X97 a_100_n134866# a_n100_n134963# a_n158_n134866# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X98 a_100_31710# a_n100_31613# a_n158_31710# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X99 a_100_73354# a_n100_73257# a_n158_73354# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X100 a_100_175310# a_n100_175213# a_n158_175310# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X101 a_100_n21422# a_n100_n21519# a_n158_n21422# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X102 a_100_7298# a_n100_7201# a_n158_7298# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X103 a_100_n63066# a_n100_n63163# a_n158_n63066# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X104 a_100_148026# a_n100_147929# a_n158_148026# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X105 a_100_87714# a_n100_87617# a_n158_87714# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X106 a_100_143718# a_n100_143621# a_n158_143718# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X107 a_100_34582# a_n100_34485# a_n158_34582# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X108 a_100_n130558# a_n100_n130655# a_n158_n130558# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X109 a_100_n24294# a_n100_n24391# a_n158_n24294# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X110 a_100_n77426# a_n100_n77523# a_n158_n77426# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X111 a_100_178182# a_n100_178085# a_n158_178182# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X112 a_100_173874# a_n100_173777# a_n158_173874# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X113 a_100_n149226# a_n100_n149323# a_n158_n149226# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X114 a_100_n144918# a_n100_n145015# a_n158_n144918# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X115 a_100_171002# a_n100_170905# a_n158_171002# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X116 a_100_109254# a_n100_109157# a_n158_109254# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X117 a_100_104946# a_n100_104849# a_n158_104946# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X118 a_100_48942# a_n100_48845# a_n158_48942# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X119 a_100_83406# a_n100_83309# a_n158_83406# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X120 a_100_n38654# a_n100_n38751# a_n158_n38654# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X121 a_100_n179382# a_n100_n179479# a_n158_n179382# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X122 a_100_30274# a_n100_30177# a_n158_30274# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X123 a_100_n172202# a_n100_n172299# a_n158_n172202# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X124 a_100_n75990# a_n100_n76087# a_n158_n75990# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X125 a_100_132230# a_n100_132133# a_n158_132230# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X126 a_100_n147790# a_n100_n147887# a_n158_n147790# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X127 a_100_n73118# a_n100_n73215# a_n158_n73118# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X128 a_100_n140610# a_n100_n140707# a_n158_n140610# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X129 a_100_100638# a_n100_100541# a_n158_100638# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X130 a_100_44634# a_n100_44537# a_n158_44634# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X131 a_100_86278# a_n100_86181# a_n158_86278# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X132 a_100_5862# a_n100_5765# a_n158_5862# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X133 a_100_n34346# a_n100_n34443# a_n158_n34346# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X134 a_100_n175074# a_n100_n175171# a_n158_n175074# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X135 a_100_119306# a_n100_119209# a_n158_119306# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X136 a_100_74790# a_n100_74693# a_n158_74790# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X137 a_100_n170766# a_n100_n170863# a_n158_n170766# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X138 a_100_n106146# a_n100_n106243# a_n158_n106146# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X139 a_100_130794# a_n100_130697# a_n158_130794# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X140 a_100_n101838# a_n100_n101935# a_n158_n101838# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X141 a_100_n48706# a_n100_n48803# a_n158_n48706# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X142 a_100_149462# a_n100_149365# a_n158_149462# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X143 a_100_40326# a_n100_40229# a_n158_40326# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X144 a_100_1554# a_n100_1457# a_n158_1554# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X145 a_100_n131994# a_n100_n132091# a_n158_n131994# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X146 a_100_n30038# a_n100_n30135# a_n158_n30038# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X147 a_100_n78862# a_n100_n78959# a_n158_n78862# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X148 a_100_70482# a_n100_70385# a_n158_70482# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X149 a_100_43198# a_n100_43101# a_n158_43198# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X150 a_100_103510# a_n100_103413# a_n158_103510# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X151 a_100_89150# a_n100_89053# a_n158_89150# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X152 a_100_n180818# a_n100_n180915# a_n158_n180818# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X153 a_100_n60194# a_n100_n60291# a_n158_n60194# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X154 a_100_145154# a_n100_145057# a_n158_145154# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X155 a_100_140846# a_n100_140749# a_n158_140846# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X156 a_100_84842# a_n100_84745# a_n158_84842# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X157 a_100_15914# a_n100_15817# a_n158_15914# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X158 a_100_57558# a_n100_57461# a_n158_57558# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X159 a_100_n74554# a_n100_n74651# a_n158_n74554# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X160 a_100_159514# a_n100_159417# a_n158_159514# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X161 a_100_n146354# a_n100_n146451# a_n158_n146354# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X162 a_100_106382# a_n100_106285# a_n158_106382# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X163 a_100_n47270# a_n100_n47367# a_n158_n47270# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X164 a_100_n183690# a_n100_n183787# a_n158_n183690# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X165 a_100_n119070# a_n100_n119167# a_n158_n119070# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X166 a_100_18786# a_n100_18689# a_n158_18786# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X167 a_100_n88914# a_n100_n89011# a_n158_n88914# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X168 a_100_80534# a_n100_80437# a_n158_80534# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X169 a_100_n35782# a_n100_n35879# a_n158_n35782# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X170 a_100_11606# a_n100_11509# a_n158_11606# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X171 a_100_n107582# a_n100_n107679# a_n158_n107582# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X172 a_100_n100402# a_n100_n100499# a_n158_n100402# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X173 a_100_n70246# a_n100_n70343# a_n158_n70246# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X174 a_100_155206# a_n100_155109# a_n158_155206# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X175 a_100_99202# a_n100_99105# a_n158_99202# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X176 a_100_n142046# a_n100_n142143# a_n158_n142046# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X177 a_100_102074# a_n100_101977# a_n158_102074# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X178 a_100_46070# a_n100_45973# a_n158_46070# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X179 a_100_41762# a_n100_41665# a_n158_41762# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X180 a_100_2990# a_n100_2893# a_n158_2990# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X181 a_100_14478# a_n100_14381# a_n158_14478# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X182 a_100_n84606# a_n100_n84703# a_n158_n84606# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X183 a_100_n31474# a_n100_n31571# a_n158_n31474# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X184 a_100_n156406# a_n100_n156503# a_n158_n156406# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X185 a_100_n103274# a_n100_n103371# a_n158_n103274# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X186 a_100_116434# a_n100_116337# a_n158_116434# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X187 a_100_158078# a_n100_157981# a_n158_158078# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X188 a_100_97766# a_n100_97669# a_n158_97766# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X189 a_100_28838# a_n100_28741# a_n158_28838# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X190 a_100_n45834# a_n100_n45931# a_n158_n45834# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X191 a_100_146590# a_n100_146493# a_n158_146590# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X192 a_100_n117634# a_n100_n117731# a_n158_n117634# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X193 a_100_n87478# a_n100_n87575# a_n158_n87478# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X194 a_100_n18550# a_n100_n18647# a_n158_n18550# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X195 a_100_n159278# a_n100_n159375# a_n158_n159278# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X196 a_100_114998# a_n100_114901# a_n158_114998# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X197 a_100_58994# a_n100_58897# a_n158_58994# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X198 a_100_n154970# a_n100_n155067# a_n158_n154970# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X199 a_100_181054# a_n100_180957# a_n158_181054# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X200 a_100_56122# a_n100_56025# a_n158_56122# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X201 a_100_112126# a_n100_112029# a_n158_112126# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X202 a_100_51814# a_n100_51717# a_n158_51814# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X203 a_100_93458# a_n100_93361# a_n158_93458# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X204 a_100_n41526# a_n100_n41623# a_n158_n41526# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X205 a_100_n182254# a_n100_n182351# a_n158_n182254# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X206 a_100_142282# a_n100_142185# a_n158_142282# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X207 a_100_81970# a_n100_81873# a_n158_81970# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X208 a_100_n9934# a_n100_n10031# a_n158_n9934# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X209 a_100_n113326# a_n100_n113423# a_n158_n113326# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X210 a_100_n83170# a_n100_n83267# a_n158_n83170# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X211 a_100_17350# a_n100_17253# a_n158_17350# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X212 a_100_54686# a_n100_54589# a_n158_54686# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X213 a_100_n71682# a_n100_n71779# a_n158_n71682# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X214 a_100_156642# a_n100_156545# a_n158_156642# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X215 a_100_n44398# a_n100_n44495# a_n158_n44398# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X216 a_100_n143482# a_n100_n143579# a_n158_n143482# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X217 a_100_n97530# a_n100_n97627# a_n158_n97530# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X218 a_100_n169330# a_n100_n169427# a_n158_n169330# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X219 a_100_n116198# a_n100_n116295# a_n158_n116198# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X220 a_100_129358# a_n100_129261# a_n158_129358# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X221 a_100_n111890# a_n100_n111987# a_n158_n111890# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X222 a_100_n5626# a_n100_n5723# a_n158_n5626# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X223 a_100_n157842# a_n100_n157939# a_n158_n157842# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X224 a_100_117870# a_n100_117773# a_n158_117870# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X225 a_100_13042# a_n100_12945# a_n158_13042# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X226 a_100_n58758# a_n100_n58855# a_n158_n58758# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X227 a_100_50378# a_n100_50281# a_n158_50378# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X228 a_100_96330# a_n100_96233# a_n158_96330# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X229 a_100_152334# a_n100_152237# a_n158_152334# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X230 a_100_27402# a_n100_27305# a_n158_27402# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X231 a_100_n40090# a_n100_n40187# a_n158_n40090# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X232 a_100_69046# a_n100_68949# a_n158_69046# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X233 a_100_n8498# a_n100_n8595# a_n158_n8498# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X234 a_100_64738# a_n100_64641# a_n158_64738# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X235 a_100_n19986# a_n100_n20083# a_n158_n19986# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X236 a_100_n86042# a_n100_n86139# a_n158_n86042# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X237 a_100_n81734# a_n100_n81831# a_n158_n81734# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X238 a_100_182490# a_n100_182393# a_n158_182490# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X239 a_100_n1318# a_n100_n1415# a_n158_n1318# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X240 a_100_n12806# a_n100_n12903# a_n158_n12806# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X241 a_100_n17114# a_n100_n17211# a_n158_n17114# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X242 a_100_n153534# a_n100_n153631# a_n158_n153534# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X243 a_100_113562# a_n100_113465# a_n158_113562# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X244 a_100_n54450# a_n100_n54547# a_n158_n54450# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X245 a_100_94894# a_n100_94797# a_n158_94894# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X246 a_100_n126250# a_n100_n126347# a_n158_n126250# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X247 a_100_150898# a_n100_150801# a_n158_150898# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X248 a_100_92022# a_n100_91925# a_n158_92022# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X249 a_100_25966# a_n100_25869# a_n158_25966# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X250 a_100_n42962# a_n100_n43059# a_n158_n42962# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X251 a_100_127922# a_n100_127825# a_n158_127922# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X252 a_100_n4190# a_n100_n4287# a_n158_n4190# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X253 a_100_n15678# a_n100_n15775# a_n158_n15678# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X254 a_100_n114762# a_n100_n114859# a_n158_n114762# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
X255 a_100_n68810# a_n100_n68907# a_n158_n68810# w_n358_n183987# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=1
C0 w_n358_n183987# a_n100_n139271# 0.269531f
C1 a_n100_n147887# a_100_n147790# 0.133664f
C2 a_n100_117773# a_100_117870# 0.133664f
C3 w_n358_n183987# a_n100_126389# 0.269531f
C4 a_100_47506# a_100_46070# 0.010536f
C5 a_n100_45973# a_n158_46070# 0.133664f
C6 w_n358_n183987# a_n158_n50142# 0.352467f
C7 w_n358_n183987# a_100_162386# 0.352467f
C8 a_n158_n103274# a_100_n103274# 0.328443f
C9 a_n100_n103371# a_n100_n104807# 0.205388f
C10 a_n100_n175171# a_100_n175074# 0.133664f
C11 a_n100_90489# a_100_90586# 0.133664f
C12 w_n358_n183987# a_n100_71821# 0.269531f
C13 a_100_20222# a_100_18786# 0.010536f
C14 a_n100_18689# a_n158_18786# 0.133664f
C15 a_n158_n14242# a_n158_n15678# 0.010536f
C16 w_n358_n183987# a_n158_n104710# 0.352467f
C17 a_n158_n130558# a_100_n130558# 0.328443f
C18 a_n100_n130655# a_n100_n132091# 0.205388f
C19 a_n158_135102# a_100_135102# 0.328443f
C20 a_n100_135005# a_n100_133569# 0.205388f
C21 a_n100_63205# a_100_63302# 0.133664f
C22 w_n358_n183987# a_100_n15678# 0.352467f
C23 w_n358_n183987# a_n100_17253# 0.269531f
C24 a_n158_n157842# a_100_n157842# 0.328443f
C25 a_n100_n157939# a_n100_n159375# 0.205388f
C26 a_n158_107818# a_100_107818# 0.328443f
C27 a_n100_107721# a_n100_106285# 0.205388f
C28 w_n358_n183987# a_n158_106382# 0.352467f
C29 a_n158_n41526# a_n158_n42962# 0.010536f
C30 w_n358_n183987# a_n158_n159278# 0.352467f
C31 a_n100_179521# a_n100_178085# 0.205388f
C32 a_n100_35921# a_100_36018# 0.133664f
C33 w_n358_n183987# a_100_n70246# 0.352467f
C34 a_n158_80534# a_100_80534# 0.328443f
C35 a_n100_80437# a_n100_79001# 0.205388f
C36 w_n358_n183987# a_n158_51814# 0.352467f
C37 a_n100_8637# a_100_8734# 0.133664f
C38 a_n158_n68810# a_n158_n70246# 0.010536f
C39 w_n358_n183987# a_100_n124814# 0.352467f
C40 w_n358_n183987# a_100_140846# 0.352467f
C41 a_n158_53250# a_100_53250# 0.328443f
C42 a_n100_53153# a_n100_51717# 0.205388f
C43 w_n358_n183987# a_n100_n37315# 0.269531f
C44 a_n158_173874# a_100_173874# 0.328443f
C45 a_n158_n96094# a_n158_n97530# 0.010536f
C46 w_n358_n183987# a_100_n179382# 0.352467f
C47 w_n358_n183987# a_100_86278# 0.352467f
C48 a_n100_159417# a_100_159514# 0.133664f
C49 a_n158_25966# a_100_25966# 0.328443f
C50 a_n100_25869# a_n100_24433# 0.205388f
C51 a_n158_n123378# a_n158_n124814# 0.010536f
C52 a_n158_142282# a_n158_140846# 0.010536f
C53 a_100_n7062# a_100_n8498# 0.010536f
C54 a_n100_n8595# a_n158_n8498# 0.133664f
C55 w_n358_n183987# a_n100_n91883# 0.269531f
C56 w_n358_n183987# a_n158_n2754# 0.352467f
C57 w_n358_n183987# a_100_31710# 0.352467f
C58 a_n158_n150662# a_n158_n152098# 0.010536f
C59 a_n158_114998# a_n158_113562# 0.010536f
C60 w_n358_n183987# a_n100_119209# 0.269531f
C61 a_100_n34346# a_100_n35782# 0.010536f
C62 a_n100_n35879# a_n158_n35782# 0.133664f
C63 w_n358_n183987# a_n100_n146451# 0.269531f
C64 a_n158_166694# a_100_166694# 0.328443f
C65 w_n358_n183987# a_n158_n57322# 0.352467f
C66 w_n358_n183987# a_n100_178085# 0.269531f
C67 a_n158_n177946# a_n158_n179382# 0.010536f
C68 a_n158_87714# a_n158_86278# 0.010536f
C69 w_n358_n183987# a_n100_64641# 0.269531f
C70 a_100_n61630# a_100_n63066# 0.010536f
C71 a_n100_n63163# a_n158_n63066# 0.133664f
C72 a_100_176746# a_n100_176649# 0.133664f
C73 w_n358_n183987# a_n158_n111890# 0.352467f
C74 w_n358_n183987# a_100_5862# 0.352467f
C75 w_n358_n183987# a_n158_153770# 0.352467f
C76 a_n100_n18647# a_100_n18550# 0.133664f
C77 a_n158_60430# a_n158_58994# 0.010536f
C78 w_n358_n183987# a_n100_10073# 0.269531f
C79 a_100_n88914# a_100_n90350# 0.010536f
C80 a_n100_n90447# a_n158_n90350# 0.133664f
C81 w_n358_n183987# a_100_n22858# 0.352467f
C82 w_n358_n183987# a_n158_n166458# 0.352467f
C83 w_n358_n183987# a_n158_99202# 0.352467f
C84 a_n100_n45931# a_100_n45834# 0.133664f
C85 a_n158_33146# a_n158_31710# 0.010536f
C86 a_100_n116198# a_100_n117634# 0.010536f
C87 a_n100_n117731# a_n158_n117634# 0.133664f
C88 a_100_149462# a_100_148026# 0.010536f
C89 a_n100_147929# a_n158_148026# 0.133664f
C90 a_n158_n1318# a_100_n1318# 0.328443f
C91 a_n100_n1415# a_n100_n2851# 0.205388f
C92 w_n358_n183987# a_100_n77426# 0.352467f
C93 a_n100_n73215# a_100_n73118# 0.133664f
C94 w_n358_n183987# a_n158_44634# 0.352467f
C95 w_n358_n183987# a_100_n131994# 0.352467f
C96 a_100_n143482# a_100_n144918# 0.010536f
C97 a_n100_n145015# a_n158_n144918# 0.133664f
C98 a_100_122178# a_100_120742# 0.010536f
C99 a_n100_120645# a_n158_120742# 0.133664f
C100 w_n358_n183987# a_100_133666# 0.352467f
C101 a_n158_n28602# a_100_n28602# 0.328443f
C102 a_n100_n28699# a_n100_n30135# 0.205388f
C103 a_n100_n100499# a_100_n100402# 0.133664f
C104 w_n358_n183987# a_n100_n44495# 0.269531f
C105 a_n158_n55886# a_100_n55886# 0.328443f
C106 a_n100_n55983# a_n100_n57419# 0.205388f
C107 a_100_n170766# a_100_n172202# 0.010536f
C108 a_n100_n172299# a_n158_n172202# 0.133664f
C109 a_100_94894# a_100_93458# 0.010536f
C110 a_n100_93361# a_n158_93458# 0.133664f
C111 w_n358_n183987# a_100_79098# 0.352467f
C112 w_n358_n183987# a_n100_n99063# 0.269531f
C113 a_n100_n127783# a_100_n127686# 0.133664f
C114 a_n100_137877# a_100_137974# 0.133664f
C115 w_n358_n183987# a_100_172438# 0.352467f
C116 a_n158_n83170# a_100_n83170# 0.328443f
C117 a_n100_n83267# a_n100_n84703# 0.205388f
C118 a_100_67610# a_100_66174# 0.010536f
C119 a_n100_66077# a_n158_66174# 0.133664f
C120 w_n358_n183987# a_100_24530# 0.352467f
C121 w_n358_n183987# a_n158_n9934# 0.352467f
C122 w_n358_n183987# a_n100_n153631# 0.269531f
C123 a_n100_n155067# a_100_n154970# 0.133664f
C124 a_n100_110593# a_100_110690# 0.133664f
C125 w_n358_n183987# a_n100_112029# 0.269531f
C126 a_100_40326# a_100_38890# 0.010536f
C127 a_n100_38793# a_n158_38890# 0.133664f
C128 w_n358_n183987# a_n158_n64502# 0.352467f
C129 a_n158_n110454# a_100_n110454# 0.328443f
C130 a_n100_n110551# a_n100_n111987# 0.205388f
C131 a_n158_155206# a_100_155206# 0.328443f
C132 a_n100_n182351# a_100_n182254# 0.133664f
C133 a_n100_83309# a_100_83406# 0.133664f
C134 w_n358_n183987# a_n100_57461# 0.269531f
C135 a_100_13042# a_100_11606# 0.010536f
C136 a_n100_11509# a_n158_11606# 0.133664f
C137 a_n158_n21422# a_n158_n22858# 0.010536f
C138 w_n358_n183987# a_n158_n119070# 0.352467f
C139 a_n158_n137738# a_100_n137738# 0.328443f
C140 a_n100_n137835# a_n100_n139271# 0.205388f
C141 a_n158_127922# a_100_127922# 0.328443f
C142 a_n100_127825# a_n100_126389# 0.205388f
C143 w_n358_n183987# a_n158_146590# 0.352467f
C144 a_n100_56025# a_100_56122# 0.133664f
C145 w_n358_n183987# a_100_n30038# 0.352467f
C146 a_n158_n48706# a_n158_n50142# 0.010536f
C147 w_n358_n183987# a_n158_n173638# 0.352467f
C148 a_n158_n165022# a_100_n165022# 0.328443f
C149 a_n100_n165119# a_n100_n166555# 0.205388f
C150 a_n158_100638# a_100_100638# 0.328443f
C151 a_n100_100541# a_n100_99105# 0.205388f
C152 w_n358_n183987# a_n158_92022# 0.352467f
C153 a_n100_28741# a_100_28838# 0.133664f
C154 a_100_163822# a_100_162386# 0.010536f
C155 a_n100_162289# a_n158_162386# 0.133664f
C156 w_n358_n183987# a_100_n84606# 0.352467f
C157 w_n358_n183987# a_n158_37454# 0.352467f
C158 a_n158_n75990# a_n158_n77426# 0.010536f
C159 a_n158_73354# a_100_73354# 0.328443f
C160 a_n100_73257# a_n100_71821# 0.205388f
C161 a_n100_21# a_100_118# 0.133664f
C162 w_n358_n183987# a_100_n139174# 0.352467f
C163 w_n358_n183987# a_100_126486# 0.352467f
C164 a_n158_46070# a_100_46070# 0.328443f
C165 a_n100_45973# a_n100_44537# 0.205388f
C166 a_n158_n103274# a_n158_n104710# 0.010536f
C167 a_n100_169469# a_100_169566# 0.133664f
C168 w_n358_n183987# a_n100_n51675# 0.269531f
C169 w_n358_n183987# a_n158_160950# 0.352467f
C170 w_n358_n183987# a_100_71918# 0.352467f
C171 a_n158_18786# a_100_18786# 0.328443f
C172 a_n100_18689# a_n100_17253# 0.205388f
C173 a_100_n14242# a_100_n15678# 0.010536f
C174 a_n100_n15775# a_n158_n15678# 0.133664f
C175 w_n358_n183987# a_n100_n106243# 0.269531f
C176 a_n158_n130558# a_n158_n131994# 0.010536f
C177 a_n158_135102# a_n158_133666# 0.010536f
C178 a_n100_4329# a_n100_2893# 0.205388f
C179 w_n358_n183987# a_n158_n17114# 0.352467f
C180 w_n358_n183987# a_100_17350# 0.352467f
C181 w_n358_n183987# a_n100_104849# 0.269531f
C182 a_100_n41526# a_100_n42962# 0.010536f
C183 a_n100_n43059# a_n158_n42962# 0.133664f
C184 w_n358_n183987# a_n100_n160811# 0.269531f
C185 a_n158_179618# a_n158_178182# 0.010536f
C186 a_n158_n157842# a_n158_n159278# 0.010536f
C187 a_n158_107818# a_n158_106382# 0.010536f
C188 w_n358_n183987# a_n158_n71682# 0.352467f
C189 a_n158_80534# a_n158_79098# 0.010536f
C190 w_n358_n183987# a_n100_50281# 0.269531f
C191 a_100_n68810# a_100_n70246# 0.010536f
C192 a_n100_n70343# a_n158_n70246# 0.133664f
C193 w_n358_n183987# a_n158_n126250# 0.352467f
C194 w_n358_n183987# a_n158_139410# 0.352467f
C195 a_n100_n25827# a_100_n25730# 0.133664f
C196 a_n158_53250# a_n158_51814# 0.010536f
C197 a_100_n96094# a_100_n97530# 0.010536f
C198 a_n100_n97627# a_n158_n97530# 0.133664f
C199 w_n358_n183987# a_100_n37218# 0.352467f
C200 a_n158_173874# a_n158_172438# 0.010536f
C201 w_n358_n183987# a_n158_n180818# 0.352467f
C202 w_n358_n183987# a_n158_84842# 0.352467f
C203 a_n100_n53111# a_100_n53014# 0.133664f
C204 a_n158_25966# a_n158_24530# 0.010536f
C205 a_100_n123378# a_100_n124814# 0.010536f
C206 a_n100_n124911# a_n158_n124814# 0.133664f
C207 a_n158_n8498# a_100_n8498# 0.328443f
C208 a_n100_n8595# a_n100_n10031# 0.205388f
C209 w_n358_n183987# a_100_n91786# 0.352467f
C210 a_100_142282# a_100_140846# 0.010536f
C211 a_n100_140749# a_n158_140846# 0.133664f
C212 w_n358_n183987# a_n100_n4287# 0.269531f
C213 w_n358_n183987# a_n158_30274# 0.352467f
C214 a_n100_n80395# a_100_n80298# 0.133664f
C215 a_100_n150662# a_100_n152098# 0.010536f
C216 a_n100_n152195# a_n158_n152098# 0.133664f
C217 a_100_114998# a_100_113562# 0.010536f
C218 a_n100_113465# a_n158_113562# 0.133664f
C219 w_n358_n183987# a_100_119306# 0.352467f
C220 a_n158_n35782# a_100_n35782# 0.328443f
C221 a_n100_n35879# a_n100_n37315# 0.205388f
C222 w_n358_n183987# a_100_n146354# 0.352467f
C223 a_n100_1457# a_n158_1554# 0.133664f
C224 w_n358_n183987# a_100_178182# 0.352467f
C225 a_100_182490# a_100_181054# 0.010536f
C226 w_n358_n183987# a_n100_n58855# 0.269531f
C227 a_n100_n107679# a_100_n107582# 0.133664f
C228 a_100_n177946# a_100_n179382# 0.010536f
C229 a_n100_n179479# a_n158_n179382# 0.133664f
C230 a_100_87714# a_100_86278# 0.010536f
C231 a_n100_86181# a_n158_86278# 0.133664f
C232 w_n358_n183987# a_100_64738# 0.352467f
C233 a_n158_n63066# a_100_n63066# 0.328443f
C234 a_n100_n63163# a_n100_n64599# 0.205388f
C235 a_n100_n134963# a_100_n134866# 0.133664f
C236 a_n100_130697# a_100_130794# 0.133664f
C237 w_n358_n183987# a_n100_152237# 0.269531f
C238 w_n358_n183987# a_n100_n113423# 0.269531f
C239 a_100_60430# a_100_58994# 0.010536f
C240 a_n100_58897# a_n158_58994# 0.133664f
C241 w_n358_n183987# a_100_10170# 0.352467f
C242 a_n158_n90350# a_100_n90350# 0.328443f
C243 a_n100_n90447# a_n100_n91883# 0.205388f
C244 w_n358_n183987# a_n158_n24294# 0.352467f
C245 a_n100_n162247# a_100_n162150# 0.133664f
C246 a_n100_103413# a_100_103510# 0.133664f
C247 w_n358_n183987# a_n100_n167991# 0.269531f
C248 a_n100_8637# a_n100_7201# 0.205388f
C249 w_n358_n183987# a_n100_97669# 0.269531f
C250 a_n158_n117634# a_100_n117634# 0.328443f
C251 a_n100_n117731# a_n100_n119167# 0.205388f
C252 a_100_33146# a_100_31710# 0.010536f
C253 a_n100_31613# a_n158_31710# 0.133664f
C254 a_n158_172438# a_n158_171002# 0.010536f
C255 a_n158_148026# a_100_148026# 0.328443f
C256 a_n100_147929# a_n100_146493# 0.205388f
C257 a_n158_n1318# a_n158_n2754# 0.010536f
C258 w_n358_n183987# a_n158_n78862# 0.352467f
C259 a_n100_76129# a_100_76226# 0.133664f
C260 w_n358_n183987# a_n100_43101# 0.269531f
C261 a_n158_n144918# a_100_n144918# 0.328443f
C262 a_n100_n145015# a_n100_n146451# 0.205388f
C263 a_n158_120742# a_100_120742# 0.328443f
C264 a_n100_120645# a_n100_119209# 0.205388f
C265 w_n358_n183987# a_n158_132230# 0.352467f
C266 a_n158_n28602# a_n158_n30038# 0.010536f
C267 w_n358_n183987# a_n158_n133430# 0.352467f
C268 a_n100_48845# a_100_48942# 0.133664f
C269 w_n358_n183987# a_100_n44398# 0.352467f
C270 a_n100_159417# a_n100_157981# 0.205388f
C271 a_n158_n172202# a_100_n172202# 0.328443f
C272 a_n100_n172299# a_n100_n173735# 0.205388f
C273 a_n158_93458# a_100_93458# 0.328443f
C274 a_n100_93361# a_n100_91925# 0.205388f
C275 w_n358_n183987# a_n158_77662# 0.352467f
C276 a_n158_n55886# a_n158_n57322# 0.010536f
C277 a_n100_182393# a_n158_182490# 0.133664f
C278 a_n100_21561# a_100_21658# 0.133664f
C279 w_n358_n183987# a_100_n98966# 0.352467f
C280 a_n158_n83170# a_n158_n84606# 0.010536f
C281 a_n158_66174# a_100_66174# 0.328443f
C282 a_n100_66077# a_n100_64641# 0.205388f
C283 w_n358_n183987# a_n158_23094# 0.352467f
C284 w_n358_n183987# a_n100_n11467# 0.269531f
C285 w_n358_n183987# a_100_n153534# 0.352467f
C286 w_n358_n183987# a_100_112126# 0.352467f
C287 a_n158_n110454# a_n158_n111890# 0.010536f
C288 a_n158_38890# a_100_38890# 0.328443f
C289 a_n100_38793# a_n100_37357# 0.205388f
C290 w_n358_n183987# a_n100_4329# 0.269531f
C291 a_n158_155206# a_n158_153770# 0.010536f
C292 w_n358_n183987# a_n100_n66035# 0.269531f
C293 a_n100_5765# a_n158_5862# 0.133664f
C294 w_n358_n183987# a_100_57558# 0.352467f
C295 a_n158_n137738# a_n158_n139174# 0.010536f
C296 a_n158_11606# a_100_11606# 0.328443f
C297 a_n100_11509# a_n100_10073# 0.205388f
C298 w_n358_n183987# a_n100_n120603# 0.269531f
C299 a_n158_127922# a_n158_126486# 0.010536f
C300 w_n358_n183987# a_n100_145057# 0.269531f
C301 a_100_n21422# a_100_n22858# 0.010536f
C302 a_n100_n22955# a_n158_n22858# 0.133664f
C303 w_n358_n183987# a_n158_n31474# 0.352467f
C304 w_n358_n183987# a_100_171002# 0.352467f
C305 a_n158_n165022# a_n158_n166458# 0.010536f
C306 a_100_n48706# a_100_n50142# 0.010536f
C307 a_n100_n50239# a_n158_n50142# 0.133664f
C308 w_n358_n183987# a_n100_n175171# 0.269531f
C309 a_n158_100638# a_n158_99202# 0.010536f
C310 w_n358_n183987# a_n100_90489# 0.269531f
C311 a_n158_162386# a_100_162386# 0.328443f
C312 a_n100_162289# a_n100_160853# 0.205388f
C313 w_n358_n183987# a_n158_n86042# 0.352467f
C314 a_n100_n5723# a_100_n5626# 0.133664f
C315 a_100_n75990# a_100_n77426# 0.010536f
C316 a_n100_n77523# a_n158_n77426# 0.133664f
C317 a_n158_73354# a_n158_71918# 0.010536f
C318 w_n358_n183987# a_n100_35921# 0.269531f
C319 w_n358_n183987# a_n158_n140610# 0.352467f
C320 w_n358_n183987# a_n158_125050# 0.352467f
C321 a_n100_n33007# a_100_n32910# 0.133664f
C322 a_100_n103274# a_100_n104710# 0.010536f
C323 a_n100_n104807# a_n158_n104710# 0.133664f
C324 a_n100_180957# a_n100_182393# 0.205388f
C325 a_n158_46070# a_n158_44634# 0.010536f
C326 w_n358_n183987# a_100_n51578# 0.352467f
C327 w_n358_n183987# a_n100_159417# 0.269531f
C328 w_n358_n183987# a_n158_70482# 0.352467f
C329 a_n100_n60291# a_100_n60194# 0.133664f
C330 a_n158_18786# a_n158_17350# 0.010536f
C331 a_100_n130558# a_100_n131994# 0.010536f
C332 a_n100_n132091# a_n158_n131994# 0.133664f
C333 a_n158_n15678# a_100_n15678# 0.328443f
C334 a_n100_n15775# a_n100_n17211# 0.205388f
C335 w_n358_n183987# a_100_n106146# 0.352467f
C336 a_100_135102# a_100_133666# 0.010536f
C337 a_n100_133569# a_n158_133666# 0.133664f
C338 a_n158_4426# a_n158_2990# 0.010536f
C339 w_n358_n183987# a_n100_n18647# 0.269531f
C340 w_n358_n183987# a_n158_15914# 0.352467f
C341 a_n100_n87575# a_100_n87478# 0.133664f
C342 a_100_n157842# a_100_n159278# 0.010536f
C343 a_n100_n159375# a_n158_n159278# 0.133664f
C344 a_100_179618# a_100_178182# 0.010536f
C345 a_n158_n42962# a_100_n42962# 0.328443f
C346 a_n100_n43059# a_n100_n44495# 0.205388f
C347 w_n358_n183987# a_100_n160714# 0.352467f
C348 a_100_107818# a_100_106382# 0.010536f
C349 a_n100_106285# a_n158_106382# 0.133664f
C350 w_n358_n183987# a_100_104946# 0.352467f
C351 w_n358_n183987# a_n100_n73215# 0.269531f
C352 a_n100_n114859# a_100_n114762# 0.133664f
C353 a_n100_150801# a_100_150898# 0.133664f
C354 w_n358_n183987# a_100_50378# 0.352467f
C355 a_n158_n70246# a_100_n70246# 0.328443f
C356 a_n100_n70343# a_n100_n71779# 0.205388f
C357 a_n158_156642# a_100_156642# 0.328443f
C358 a_n100_156545# a_n100_155109# 0.205388f
C359 a_100_80534# a_100_79098# 0.010536f
C360 a_n100_79001# a_n158_79098# 0.133664f
C361 w_n358_n183987# a_n100_n127783# 0.269531f
C362 a_n100_n142143# a_100_n142046# 0.133664f
C363 a_n100_123517# a_100_123614# 0.133664f
C364 w_n358_n183987# a_n100_137877# 0.269531f
C365 a_100_53250# a_100_51814# 0.010536f
C366 a_n100_51717# a_n158_51814# 0.133664f
C367 a_n158_n97530# a_100_n97530# 0.328443f
C368 a_n100_n97627# a_n100_n99063# 0.205388f
C369 a_100_159514# a_100_158078# 0.010536f
C370 w_n358_n183987# a_n158_n38654# 0.352467f
C371 a_n100_172341# a_n158_172438# 0.133664f
C372 a_100_173874# a_100_172438# 0.010536f
C373 w_n358_n183987# a_n100_83309# 0.269531f
C374 a_n158_118# a_100_118# 0.328443f
C375 a_n100_21# a_n100_n1415# 0.205388f
C376 w_n358_n183987# a_n100_n182351# 0.269531f
C377 a_n100_n169427# a_100_n169330# 0.133664f
C378 a_n100_96233# a_100_96330# 0.133664f
C379 a_100_25966# a_100_24530# 0.010536f
C380 a_n100_24433# a_n158_24530# 0.133664f
C381 a_n158_n124814# a_100_n124814# 0.328443f
C382 a_n100_n124911# a_n100_n126347# 0.205388f
C383 w_n358_n183987# a_n158_182490# 0.35701f
C384 a_n158_n8498# a_n158_n9934# 0.010536f
C385 w_n358_n183987# a_n158_n93222# 0.352467f
C386 a_n158_140846# a_100_140846# 0.328443f
C387 a_n100_140749# a_n100_139313# 0.205388f
C388 a_n100_68949# a_100_69046# 0.133664f
C389 w_n358_n183987# a_n100_28741# 0.269531f
C390 w_n358_n183987# a_100_n4190# 0.352467f
C391 a_n158_n152098# a_100_n152098# 0.328443f
C392 a_n100_n152195# a_n100_n153631# 0.205388f
C393 w_n358_n183987# a_n158_117870# 0.352467f
C394 a_n158_n35782# a_n158_n37218# 0.010536f
C395 w_n358_n183987# a_n158_n147790# 0.352467f
C396 a_n158_1554# a_100_1554# 0.328443f
C397 a_n158_113562# a_100_113562# 0.328443f
C398 a_n100_113465# a_n100_112029# 0.205388f
C399 a_n100_41665# a_100_41762# 0.133664f
C400 w_n358_n183987# a_n158_176746# 0.352467f
C401 a_n100_180957# a_n100_179521# 0.205388f
C402 w_n358_n183987# a_100_n58758# 0.352467f
C403 a_n100_156545# a_100_156642# 0.133664f
C404 a_n158_181054# a_100_181054# 0.328443f
C405 a_n158_n179382# a_100_n179382# 0.328443f
C406 a_n100_n179479# a_n100_n180915# 0.205388f
C407 a_n158_86278# a_100_86278# 0.328443f
C408 a_n100_86181# a_n100_84745# 0.205388f
C409 w_n358_n183987# a_n158_63302# 0.352467f
C410 a_n158_n63066# a_n158_n64502# 0.010536f
C411 a_n100_14381# a_100_14478# 0.133664f
C412 w_n358_n183987# a_100_152334# 0.352467f
C413 w_n358_n183987# a_100_n113326# 0.352467f
C414 a_n158_58994# a_100_58994# 0.328443f
C415 a_n100_58897# a_n100_57461# 0.205388f
C416 w_n358_n183987# a_n158_8734# 0.352467f
C417 a_n158_n90350# a_n158_n91786# 0.010536f
C418 w_n358_n183987# a_n100_n25827# 0.269531f
C419 w_n358_n183987# a_100_97766# 0.352467f
C420 w_n358_n183987# a_100_n167894# 0.352467f
C421 a_n158_8734# a_n158_7298# 0.010536f
C422 a_n100_165161# a_100_165258# 0.133664f
C423 a_n158_31710# a_100_31710# 0.328443f
C424 a_n100_31613# a_n100_30177# 0.205388f
C425 a_n100_170905# a_n158_171002# 0.133664f
C426 a_n158_n117634# a_n158_n119070# 0.010536f
C427 a_100_n1318# a_100_n2754# 0.010536f
C428 a_n100_n2851# a_n158_n2754# 0.133664f
C429 w_n358_n183987# a_n100_n80395# 0.269531f
C430 a_n158_148026# a_n158_146590# 0.010536f
C431 w_n358_n183987# a_100_43198# 0.352467f
C432 a_n158_n144918# a_n158_n146354# 0.010536f
C433 a_100_158078# a_100_156642# 0.010536f
C434 a_n100_156545# a_n158_156642# 0.133664f
C435 a_n158_120742# a_n158_119306# 0.010536f
C436 w_n358_n183987# a_n100_130697# 0.269531f
C437 a_100_n28602# a_100_n30038# 0.010536f
C438 a_n100_n30135# a_n158_n30038# 0.133664f
C439 w_n358_n183987# a_n100_n134963# 0.269531f
C440 w_n358_n183987# a_n158_n45834# 0.352467f
C441 a_n158_n172202# a_n158_n173638# 0.010536f
C442 w_n358_n183987# a_n100_180957# 0.269531f
C443 a_n158_93458# a_n158_92022# 0.010536f
C444 w_n358_n183987# a_n100_76129# 0.269531f
C445 a_100_n55886# a_100_n57322# 0.010536f
C446 a_n100_n57419# a_n158_n57322# 0.133664f
C447 w_n358_n183987# a_n158_n100402# 0.352467f
C448 a_n100_n12903# a_100_n12806# 0.133664f
C449 a_n158_66174# a_n158_64738# 0.010536f
C450 w_n358_n183987# a_n100_21561# 0.269531f
C451 a_100_n83170# a_100_n84606# 0.010536f
C452 a_n100_n84703# a_n158_n84606# 0.133664f
C453 w_n358_n183987# a_100_n11370# 0.352467f
C454 w_n358_n183987# a_n158_110690# 0.352467f
C455 w_n358_n183987# a_n158_n154970# 0.352467f
C456 a_n100_n40187# a_100_n40090# 0.133664f
C457 a_100_n110454# a_100_n111890# 0.010536f
C458 a_n100_n111987# a_n158_n111890# 0.133664f
C459 a_n158_38890# a_n158_37454# 0.010536f
C460 w_n358_n183987# a_100_4426# 0.352467f
C461 a_100_155206# a_100_153770# 0.010536f
C462 a_n100_153673# a_n158_153770# 0.133664f
C463 w_n358_n183987# a_100_n65938# 0.352467f
C464 a_n158_5862# a_100_5862# 0.328443f
C465 w_n358_n183987# a_n158_56122# 0.352467f
C466 a_n100_n67471# a_100_n67374# 0.133664f
C467 a_100_n137738# a_100_n139174# 0.010536f
C468 a_n100_n139271# a_n158_n139174# 0.133664f
C469 a_n158_11606# a_n158_10170# 0.010536f
C470 a_100_127922# a_100_126486# 0.010536f
C471 a_n100_126389# a_n158_126486# 0.133664f
C472 w_n358_n183987# a_100_145154# 0.352467f
C473 a_n158_n22858# a_100_n22858# 0.328443f
C474 a_n100_n22955# a_n100_n24391# 0.205388f
C475 w_n358_n183987# a_100_n120506# 0.352467f
C476 a_n100_n94755# a_100_n94658# 0.133664f
C477 w_n358_n183987# a_n100_n33007# 0.269531f
C478 w_n358_n183987# a_n158_169566# 0.352467f
C479 a_100_n165022# a_100_n166458# 0.010536f
C480 a_n100_n166555# a_n158_n166458# 0.133664f
C481 w_n358_n183987# a_100_n175074# 0.352467f
C482 a_100_100638# a_100_99202# 0.010536f
C483 a_n100_99105# a_n158_99202# 0.133664f
C484 w_n358_n183987# a_100_90586# 0.352467f
C485 a_n158_n50142# a_100_n50142# 0.328443f
C486 a_n100_n50239# a_n100_n51675# 0.205388f
C487 a_n158_162386# a_n158_160950# 0.010536f
C488 a_n100_n122039# a_100_n121942# 0.133664f
C489 a_n100_143621# a_100_143718# 0.133664f
C490 w_n358_n183987# a_n100_n87575# 0.269531f
C491 a_n158_n77426# a_100_n77426# 0.328443f
C492 a_n100_n77523# a_n100_n78959# 0.205388f
C493 a_100_73354# a_100_71918# 0.010536f
C494 a_n100_71821# a_n158_71918# 0.133664f
C495 w_n358_n183987# a_100_36018# 0.352467f
C496 w_n358_n183987# a_n100_n142143# 0.269531f
C497 a_n100_n149323# a_100_n149226# 0.133664f
C498 a_n100_116337# a_100_116434# 0.133664f
C499 w_n358_n183987# a_n100_123517# 0.269531f
C500 a_n158_158078# a_n158_156642# 0.010536f
C501 a_n158_n104710# a_100_n104710# 0.328443f
C502 a_n100_n104807# a_n100_n106243# 0.205388f
C503 a_100_46070# a_100_44634# 0.010536f
C504 a_n100_44537# a_n158_44634# 0.133664f
C505 w_n358_n183987# a_100_159514# 0.352467f
C506 w_n358_n183987# a_n158_n53014# 0.352467f
C507 a_n100_n176607# a_100_n176510# 0.133664f
C508 a_n100_89053# a_100_89150# 0.133664f
C509 w_n358_n183987# a_n100_68949# 0.269531f
C510 a_n158_n131994# a_100_n131994# 0.328443f
C511 a_n100_n132091# a_n100_n133527# 0.205388f
C512 a_100_18786# a_100_17350# 0.010536f
C513 a_n100_17253# a_n158_17350# 0.133664f
C514 w_n358_n183987# a_n158_n107582# 0.352467f
C515 a_100_4426# a_100_2990# 0.010536f
C516 a_n158_133666# a_100_133666# 0.328443f
C517 a_n100_133569# a_n100_132133# 0.205388f
C518 a_n158_n15678# a_n158_n17114# 0.010536f
C519 a_n100_61769# a_100_61866# 0.133664f
C520 w_n358_n183987# a_n100_14381# 0.269531f
C521 w_n358_n183987# a_100_n18550# 0.352467f
C522 a_n158_n159278# a_100_n159278# 0.328443f
C523 a_n100_n159375# a_n100_n160811# 0.205388f
C524 a_n158_n42962# a_n158_n44398# 0.010536f
C525 w_n358_n183987# a_n158_n162150# 0.352467f
C526 a_n158_106382# a_100_106382# 0.328443f
C527 a_n100_106285# a_n100_104849# 0.205388f
C528 w_n358_n183987# a_n158_103510# 0.352467f
C529 a_n100_34485# a_100_34582# 0.133664f
C530 w_n358_n183987# a_100_n73118# 0.352467f
C531 w_n358_n183987# a_n100_155109# 0.269531f
C532 a_n158_n70246# a_n158_n71682# 0.010536f
C533 a_n158_79098# a_100_79098# 0.328443f
C534 a_n100_79001# a_n100_77565# 0.205388f
C535 w_n358_n183987# a_n158_48942# 0.352467f
C536 w_n358_n183987# a_100_n127686# 0.352467f
C537 w_n358_n183987# a_100_137974# 0.352467f
C538 a_n158_n97530# a_n158_n98966# 0.010536f
C539 a_n158_51814# a_100_51814# 0.328443f
C540 a_n100_51717# a_n100_50281# 0.205388f
C541 w_n358_n183987# a_n100_n40187# 0.269531f
C542 a_n100_172341# a_n100_170905# 0.205388f
C543 a_n158_172438# a_100_172438# 0.328443f
C544 w_n358_n183987# a_100_n182254# 0.352467f
C545 w_n358_n183987# a_100_83406# 0.352467f
C546 a_n158_24530# a_100_24530# 0.328443f
C547 a_n100_24433# a_n100_22997# 0.205388f
C548 a_n158_n124814# a_n158_n126250# 0.010536f
C549 a_100_n8498# a_100_n9934# 0.010536f
C550 a_n100_n10031# a_n158_n9934# 0.133664f
C551 w_n358_n183987# a_n100_n94755# 0.269531f
C552 a_n158_140846# a_n158_139410# 0.010536f
C553 w_n358_n183987# a_100_28838# 0.352467f
C554 w_n358_n183987# a_n158_n5626# 0.352467f
C555 a_n158_n152098# a_n158_n153534# 0.010536f
C556 a_100_n35782# a_100_n37218# 0.010536f
C557 a_n100_n37315# a_n158_n37218# 0.133664f
C558 w_n358_n183987# a_100_156642# 0.352467f
C559 w_n358_n183987# a_n100_n149323# 0.269531f
C560 a_n158_113562# a_n158_112126# 0.010536f
C561 w_n358_n183987# a_n100_116337# 0.269531f
C562 a_n158_181054# a_n158_179618# 0.010536f
C563 w_n358_n183987# a_n158_n60194# 0.352467f
C564 a_n158_158078# a_100_158078# 0.328443f
C565 a_n100_157981# a_n100_156545# 0.205388f
C566 a_n158_n179382# a_n158_n180818# 0.010536f
C567 w_n358_n183987# a_n100_61769# 0.269531f
C568 a_100_n63066# a_100_n64502# 0.010536f
C569 a_n100_n64599# a_n158_n64502# 0.133664f
C570 a_n158_86278# a_n158_84842# 0.010536f
C571 w_n358_n183987# a_n158_n114762# 0.352467f
C572 w_n358_n183987# a_n158_150898# 0.352467f
C573 a_n100_n20083# a_100_n19986# 0.133664f
C574 a_n158_58994# a_n158_57558# 0.010536f
C575 a_100_n90350# a_100_n91786# 0.010536f
C576 a_n100_n91883# a_n158_n91786# 0.133664f
C577 w_n358_n183987# a_100_n25730# 0.352467f
C578 w_n358_n183987# a_n158_96330# 0.352467f
C579 w_n358_n183987# a_n158_n169330# 0.352467f
C580 a_100_8734# a_100_7298# 0.010536f
C581 a_n100_n47367# a_100_n47270# 0.133664f
C582 a_n158_31710# a_n158_30274# 0.010536f
C583 a_100_n117634# a_100_n119070# 0.010536f
C584 a_n100_n119167# a_n158_n119070# 0.133664f
C585 a_n158_n2754# a_100_n2754# 0.328443f
C586 a_n100_n2851# a_n100_n4287# 0.205388f
C587 w_n358_n183987# a_100_n80298# 0.352467f
C588 a_100_148026# a_100_146590# 0.010536f
C589 a_n100_146493# a_n158_146590# 0.133664f
C590 w_n358_n183987# a_n158_41762# 0.352467f
C591 a_n100_n74651# a_100_n74554# 0.133664f
C592 w_n358_n183987# a_n158_156642# 0.352467f
C593 a_100_n144918# a_100_n146354# 0.010536f
C594 a_n100_n146451# a_n158_n146354# 0.133664f
C595 w_n358_n183987# a_100_130794# 0.352467f
C596 a_n158_n30038# a_100_n30038# 0.328443f
C597 a_n100_n30135# a_n100_n31571# 0.205388f
C598 w_n358_n183987# a_100_n134866# 0.352467f
C599 a_n100_157981# a_100_158078# 0.133664f
C600 a_100_120742# a_100_119306# 0.010536f
C601 a_n100_119209# a_n158_119306# 0.133664f
C602 w_n358_n183987# a_n158_165258# 0.352467f
C603 w_n358_n183987# a_n100_n47367# 0.269531f
C604 a_n100_n101935# a_100_n101838# 0.133664f
C605 a_100_n172202# a_100_n173638# 0.010536f
C606 a_n100_n173735# a_n158_n173638# 0.133664f
C607 a_n100_178085# a_n158_178182# 0.133664f
C608 a_100_93458# a_100_92022# 0.010536f
C609 a_n100_91925# a_n158_92022# 0.133664f
C610 w_n358_n183987# a_100_76226# 0.352467f
C611 a_n158_n57322# a_100_n57322# 0.328443f
C612 a_n100_n57419# a_n100_n58855# 0.205388f
C613 w_n358_n183987# a_n100_n101935# 0.269531f
C614 a_n100_n129219# a_100_n129122# 0.133664f
C615 a_n100_136441# a_100_136538# 0.133664f
C616 a_100_66174# a_100_64738# 0.010536f
C617 a_n100_64641# a_n158_64738# 0.133664f
C618 w_n358_n183987# a_100_21658# 0.352467f
C619 a_n158_n84606# a_100_n84606# 0.328443f
C620 a_n100_n84703# a_n100_n86139# 0.205388f
C621 w_n358_n183987# a_n158_n12806# 0.352467f
C622 a_n100_n156503# a_100_n156406# 0.133664f
C623 a_n100_109157# a_100_109254# 0.133664f
C624 w_n358_n183987# a_n100_109157# 0.269531f
C625 w_n358_n183987# a_n100_n156503# 0.269531f
C626 a_n100_165161# a_n100_166597# 0.205388f
C627 a_100_38890# a_100_37454# 0.010536f
C628 a_n100_37357# a_n158_37454# 0.133664f
C629 w_n358_n183987# a_n100_156545# 0.269531f
C630 a_n158_n111890# a_100_n111890# 0.328443f
C631 a_n100_n111987# a_n100_n113423# 0.205388f
C632 w_n358_n183987# a_n158_n67374# 0.352467f
C633 a_n158_153770# a_100_153770# 0.328443f
C634 a_n100_153673# a_n100_152237# 0.205388f
C635 a_n100_n183787# a_100_n183690# 0.133664f
C636 a_n100_81873# a_100_81970# 0.133664f
C637 w_n358_n183987# a_n100_54589# 0.269531f
C638 a_n100_157981# a_n158_158078# 0.133664f
C639 w_n358_n183987# a_n100_175213# 0.269531f
C640 a_n158_n139174# a_100_n139174# 0.328443f
C641 a_n100_n139271# a_n100_n140707# 0.205388f
C642 a_100_11606# a_100_10170# 0.010536f
C643 a_n100_10073# a_n158_10170# 0.133664f
C644 a_n158_126486# a_100_126486# 0.328443f
C645 a_n100_126389# a_n100_124953# 0.205388f
C646 w_n358_n183987# a_n158_143718# 0.352467f
C647 a_n158_n22858# a_n158_n24294# 0.010536f
C648 w_n358_n183987# a_n158_n121942# 0.352467f
C649 a_n100_54589# a_100_54686# 0.133664f
C650 w_n358_n183987# a_100_n32910# 0.352467f
C651 a_n158_n166458# a_100_n166458# 0.328443f
C652 a_n100_n166555# a_n100_n167991# 0.205388f
C653 w_n358_n183987# a_n100_168033# 0.269531f
C654 a_n100_175213# a_100_175310# 0.133664f
C655 a_n158_99202# a_100_99202# 0.328443f
C656 a_n100_99105# a_n100_97669# 0.205388f
C657 w_n358_n183987# a_n158_89150# 0.352467f
C658 a_n158_n50142# a_n158_n51578# 0.010536f
C659 a_100_162386# a_100_160950# 0.010536f
C660 a_n100_160853# a_n158_160950# 0.133664f
C661 w_n358_n183987# a_n158_n176510# 0.352467f
C662 a_n100_27305# a_100_27402# 0.133664f
C663 w_n358_n183987# a_100_n87478# 0.352467f
C664 a_n158_71918# a_100_71918# 0.328443f
C665 a_n100_71821# a_n100_70385# 0.205388f
C666 w_n358_n183987# a_n158_34582# 0.352467f
C667 a_n158_n77426# a_n158_n78862# 0.010536f
C668 w_n358_n183987# a_100_158078# 0.352467f
C669 w_n358_n183987# a_100_123614# 0.352467f
C670 w_n358_n183987# a_100_n142046# 0.352467f
C671 a_n158_n104710# a_n158_n106146# 0.010536f
C672 a_n158_44634# a_100_44634# 0.328443f
C673 a_n100_44537# a_n100_43101# 0.205388f
C674 a_n100_168033# a_100_168130# 0.133664f
C675 w_n358_n183987# a_n100_n54547# 0.269531f
C676 w_n358_n183987# a_100_69046# 0.352467f
C677 w_n358_n183987# a_n100_2893# 0.269531f
C678 a_n158_n131994# a_n158_n133430# 0.010536f
C679 a_n158_17350# a_100_17350# 0.328443f
C680 a_n100_17253# a_n100_15817# 0.205388f
C681 a_n158_133666# a_n158_132230# 0.010536f
C682 a_100_n15678# a_100_n17114# 0.010536f
C683 a_n100_n17211# a_n158_n17114# 0.133664f
C684 w_n358_n183987# a_n100_n109115# 0.269531f
C685 w_n358_n183987# a_100_14478# 0.352467f
C686 w_n358_n183987# a_n158_n19986# 0.352467f
C687 a_n158_n159278# a_n158_n160714# 0.010536f
C688 w_n358_n183987# a_n100_182393# 0.349164f
C689 w_n358_n183987# a_n100_n163683# 0.269531f
C690 a_n158_106382# a_n158_104946# 0.010536f
C691 w_n358_n183987# a_n100_101977# 0.269531f
C692 a_100_n42962# a_100_n44398# 0.010536f
C693 a_n100_n44495# a_n158_n44398# 0.133664f
C694 w_n358_n183987# a_n158_n74554# 0.352467f
C695 w_n358_n183987# a_n158_158078# 0.352467f
C696 a_100_n70246# a_100_n71682# 0.010536f
C697 a_n100_n71779# a_n158_n71682# 0.133664f
C698 a_n158_79098# a_n158_77662# 0.010536f
C699 w_n358_n183987# a_n100_47409# 0.269531f
C700 w_n358_n183987# a_n158_n129122# 0.352467f
C701 w_n358_n183987# a_n158_136538# 0.352467f
C702 a_n100_n27263# a_100_n27166# 0.133664f
C703 a_100_n97530# a_100_n98966# 0.010536f
C704 a_n100_n99063# a_n158_n98966# 0.133664f
C705 a_n158_51814# a_n158_50378# 0.010536f
C706 w_n358_n183987# a_100_n40090# 0.352467f
C707 w_n358_n183987# a_n158_n183690# 0.35701f
C708 w_n358_n183987# a_n158_81970# 0.352467f
C709 a_n100_n54547# a_100_n54450# 0.133664f
C710 a_100_n124814# a_100_n126250# 0.010536f
C711 a_n100_n126347# a_n158_n126250# 0.133664f
C712 a_n158_24530# a_n158_23094# 0.010536f
C713 w_n358_n183987# a_100_n94658# 0.352467f
C714 a_100_140846# a_100_139410# 0.010536f
C715 a_n100_139313# a_n158_139410# 0.133664f
C716 a_n158_n9934# a_100_n9934# 0.328443f
C717 a_n100_n10031# a_n100_n11467# 0.205388f
C718 w_n358_n183987# a_n158_27402# 0.352467f
C719 a_n100_n81831# a_100_n81734# 0.133664f
C720 w_n358_n183987# a_n100_n7159# 0.269531f
C721 a_100_n152098# a_100_n153534# 0.010536f
C722 a_n100_n153631# a_n158_n153534# 0.133664f
C723 a_n158_n37218# a_100_n37218# 0.328443f
C724 a_n100_n37315# a_n100_n38751# 0.205388f
C725 w_n358_n183987# a_100_n149226# 0.352467f
C726 a_100_113562# a_100_112126# 0.010536f
C727 a_n100_112029# a_n158_112126# 0.133664f
C728 w_n358_n183987# a_100_116434# 0.352467f
C729 w_n358_n183987# a_n100_157981# 0.269531f
C730 a_n100_2893# a_100_2990# 0.133664f
C731 w_n358_n183987# a_n100_n61727# 0.269531f
C732 a_n100_n109115# a_100_n109018# 0.133664f
C733 a_100_n179382# a_100_n180818# 0.010536f
C734 a_n100_n180915# a_n158_n180818# 0.133664f
C735 a_n158_n64502# a_100_n64502# 0.328443f
C736 a_n100_n64599# a_n100_n66035# 0.205388f
C737 a_100_86278# a_100_84842# 0.010536f
C738 a_n100_84745# a_n158_84842# 0.133664f
C739 w_n358_n183987# a_100_61866# 0.352467f
C740 w_n358_n183987# a_n100_n116295# 0.269531f
C741 a_n100_n136399# a_100_n136302# 0.133664f
C742 a_n100_129261# a_100_129358# 0.133664f
C743 w_n358_n183987# a_n100_149365# 0.269531f
C744 a_n158_n91786# a_100_n91786# 0.328443f
C745 a_n100_n91883# a_n100_n93319# 0.205388f
C746 a_100_58994# a_100_57558# 0.010536f
C747 a_n100_57461# a_n158_57558# 0.133664f
C748 w_n358_n183987# a_n158_n27166# 0.352467f
C749 w_n358_n183987# a_n100_179521# 0.269531f
C750 a_n100_155109# a_n158_155206# 0.133664f
C751 w_n358_n183987# a_n100_n170863# 0.269531f
C752 a_n100_n163683# a_100_n163586# 0.133664f
C753 a_n100_101977# a_100_102074# 0.133664f
C754 w_n358_n183987# a_n100_94797# 0.269531f
C755 a_100_31710# a_100_30274# 0.010536f
C756 a_n100_30177# a_n158_30274# 0.133664f
C757 a_n158_n119070# a_100_n119070# 0.328443f
C758 a_n100_n119167# a_n100_n120603# 0.205388f
C759 a_n158_146590# a_100_146590# 0.328443f
C760 a_n100_146493# a_n100_145057# 0.205388f
C761 a_n158_n2754# a_n158_n4190# 0.010536f
C762 w_n358_n183987# a_n158_n81734# 0.352467f
C763 w_n358_n183987# a_n100_40229# 0.269531f
C764 a_n100_74693# a_100_74790# 0.133664f
C765 a_n158_n146354# a_100_n146354# 0.328443f
C766 a_n100_n146451# a_n100_n147887# 0.205388f
C767 w_n358_n183987# a_n158_129358# 0.352467f
C768 a_n158_n30038# a_n158_n31474# 0.010536f
C769 w_n358_n183987# a_n158_n136302# 0.352467f
C770 a_n158_119306# a_100_119306# 0.328443f
C771 a_n100_119209# a_n100_117773# 0.205388f
C772 a_n100_47409# a_100_47506# 0.133664f
C773 a_n158_178182# a_100_178182# 0.328443f
C774 w_n358_n183987# a_100_n47270# 0.352467f
C775 a_n100_178085# a_n100_176649# 0.205388f
C776 w_n358_n183987# a_n100_163725# 0.269531f
C777 a_n158_n173638# a_100_n173638# 0.328443f
C778 a_n100_n173735# a_n100_n175171# 0.205388f
C779 w_n358_n183987# a_n158_74790# 0.352467f
C780 a_n158_n57322# a_n158_n58758# 0.010536f
C781 a_n158_92022# a_100_92022# 0.328443f
C782 a_n100_91925# a_n100_90489# 0.205388f
C783 a_n100_20125# a_100_20222# 0.133664f
C784 w_n358_n183987# a_100_n101838# 0.352467f
C785 a_n158_64738# a_100_64738# 0.328443f
C786 a_n100_64641# a_n100_63205# 0.205388f
C787 w_n358_n183987# a_n158_20222# 0.352467f
C788 a_n158_n84606# a_n158_n86042# 0.010536f
C789 w_n358_n183987# a_n100_n14339# 0.269531f
C790 w_n358_n183987# a_100_109254# 0.352467f
C791 w_n358_n183987# a_100_n156406# 0.352467f
C792 a_n158_37454# a_100_37454# 0.328443f
C793 a_n100_37357# a_n100_35921# 0.205388f
C794 a_n158_165258# a_n158_166694# 0.010536f
C795 a_n158_n111890# a_n158_n113326# 0.010536f
C796 a_n158_153770# a_n158_152334# 0.010536f
C797 w_n358_n183987# a_n100_n68907# 0.269531f
C798 w_n358_n183987# a_n158_7298# 0.352467f
C799 w_n358_n183987# a_100_54686# 0.352467f
C800 a_n100_7201# a_100_7298# 0.133664f
C801 w_n358_n183987# a_100_175310# 0.352467f
C802 a_n158_126486# a_n158_125050# 0.010536f
C803 a_n158_10170# a_100_10170# 0.328443f
C804 a_n100_10073# a_n100_8637# 0.205388f
C805 a_n158_n139174# a_n158_n140610# 0.010536f
C806 w_n358_n183987# a_n100_142185# 0.269531f
C807 a_100_n22858# a_100_n24294# 0.010536f
C808 a_n100_n24391# a_n158_n24294# 0.133664f
C809 w_n358_n183987# a_n100_n123475# 0.269531f
C810 w_n358_n183987# a_n158_n34346# 0.352467f
C811 a_n158_n166458# a_n158_n167894# 0.010536f
C812 w_n358_n183987# a_100_168130# 0.352467f
C813 a_n158_99202# a_n158_97766# 0.010536f
C814 w_n358_n183987# a_n100_87617# 0.269531f
C815 a_100_n50142# a_100_n51578# 0.010536f
C816 a_n100_n51675# a_n158_n51578# 0.133664f
C817 a_n158_160950# a_100_160950# 0.328443f
C818 a_n100_160853# a_n100_159417# 0.205388f
C819 a_n158_156642# a_n158_155206# 0.010536f
C820 w_n358_n183987# a_n100_n178043# 0.269531f
C821 w_n358_n183987# a_n158_n88914# 0.352467f
C822 a_n100_n7159# a_100_n7062# 0.133664f
C823 a_n158_71918# a_n158_70482# 0.010536f
C824 w_n358_n183987# a_n100_33049# 0.269531f
C825 a_100_n77426# a_100_n78862# 0.010536f
C826 a_n100_n78959# a_n158_n78862# 0.133664f
C827 w_n358_n183987# a_n158_122178# 0.352467f
C828 a_n158_1554# a_n158_118# 0.010536f
C829 w_n358_n183987# a_n158_n143482# 0.352467f
C830 a_n100_n34443# a_100_n34346# 0.133664f
C831 a_n158_44634# a_n158_43198# 0.010536f
C832 a_100_n104710# a_100_n106146# 0.010536f
C833 a_n100_n106243# a_n158_n106146# 0.133664f
C834 w_n358_n183987# a_100_n54450# 0.352467f
C835 w_n358_n183987# a_n158_67610# 0.352467f
C836 a_n100_n61727# a_100_n61630# 0.133664f
C837 a_100_n131994# a_100_n133430# 0.010536f
C838 a_n100_n133527# a_n158_n133430# 0.133664f
C839 a_100_133666# a_100_132230# 0.010536f
C840 a_n100_132133# a_n158_132230# 0.133664f
C841 a_n158_17350# a_n158_15914# 0.010536f
C842 w_n358_n183987# a_100_2990# 0.352467f
C843 a_n158_n17114# a_100_n17114# 0.328443f
C844 a_n100_n17211# a_n100_n18647# 0.205388f
C845 w_n358_n183987# a_100_n109018# 0.352467f
C846 w_n358_n183987# a_n158_13042# 0.352467f
C847 w_n358_n183987# a_n100_n21519# 0.269531f
C848 a_n100_n89011# a_100_n88914# 0.133664f
C849 a_100_n159278# a_100_n160714# 0.010536f
C850 a_n100_n160811# a_n158_n160714# 0.133664f
C851 a_100_106382# a_100_104946# 0.010536f
C852 a_n100_104849# a_n158_104946# 0.133664f
C853 w_n358_n183987# a_100_102074# 0.352467f
C854 a_n158_n44398# a_100_n44398# 0.328443f
C855 a_n100_n44495# a_n100_n45931# 0.205388f
C856 w_n358_n183987# a_100_n163586# 0.352467f
C857 a_n100_n116295# a_100_n116198# 0.133664f
C858 a_n100_149365# a_100_149462# 0.133664f
C859 w_n358_n183987# a_n100_n76087# 0.269531f
C860 a_100_79098# a_100_77662# 0.010536f
C861 a_n100_77565# a_n158_77662# 0.133664f
C862 w_n358_n183987# a_100_47506# 0.352467f
C863 a_n158_n71682# a_100_n71682# 0.328443f
C864 a_n100_n71779# a_n100_n73215# 0.205388f
C865 a_n100_n143579# a_100_n143482# 0.133664f
C866 a_n100_122081# a_100_122178# 0.133664f
C867 w_n358_n183987# a_n100_135005# 0.269531f
C868 w_n358_n183987# a_n100_n130655# 0.269531f
C869 a_n100_179521# a_100_179618# 0.133664f
C870 a_n158_n98966# a_100_n98966# 0.328443f
C871 a_n100_n99063# a_n100_n100499# 0.205388f
C872 a_100_51814# a_100_50378# 0.010536f
C873 a_n100_50281# a_n158_50378# 0.133664f
C874 w_n358_n183987# a_n158_n41526# 0.352467f
C875 a_n100_n170863# a_100_n170766# 0.133664f
C876 a_n100_94797# a_100_94894# 0.133664f
C877 w_n358_n183987# a_n100_80437# 0.269531f
C878 a_n158_n126250# a_100_n126250# 0.328443f
C879 a_n100_n126347# a_n100_n127783# 0.205388f
C880 a_n158_139410# a_100_139410# 0.328443f
C881 a_n100_139313# a_n100_137877# 0.205388f
C882 a_100_24530# a_100_23094# 0.010536f
C883 a_n100_22997# a_n158_23094# 0.133664f
C884 a_n158_n9934# a_n158_n11370# 0.010536f
C885 w_n358_n183987# a_n158_n96094# 0.352467f
C886 a_n100_67513# a_100_67610# 0.133664f
C887 w_n358_n183987# a_n100_25869# 0.269531f
C888 w_n358_n183987# a_100_n7062# 0.352467f
C889 a_n158_n153534# a_100_n153534# 0.328443f
C890 a_n100_n153631# a_n100_n155067# 0.205388f
C891 a_n158_112126# a_100_112126# 0.328443f
C892 a_n100_112029# a_n100_110593# 0.205388f
C893 w_n358_n183987# a_n158_n150662# 0.352467f
C894 w_n358_n183987# a_n158_114998# 0.352467f
C895 a_n158_n37218# a_n158_n38654# 0.010536f
C896 a_n158_175310# a_n158_173874# 0.010536f
C897 a_n100_40229# a_100_40326# 0.133664f
C898 w_n358_n183987# a_100_n61630# 0.352467f
C899 a_n158_n180818# a_100_n180818# 0.328443f
C900 a_n100_n180915# a_n100_n182351# 0.205388f
C901 a_n158_84842# a_100_84842# 0.328443f
C902 a_n100_84745# a_n100_83309# 0.205388f
C903 a_n158_n64502# a_n158_n65938# 0.010536f
C904 w_n358_n183987# a_n158_60430# 0.352467f
C905 a_n100_170905# a_100_171002# 0.133664f
C906 a_n100_12945# a_100_13042# 0.133664f
C907 w_n358_n183987# a_100_n116198# 0.352467f
C908 w_n358_n183987# a_100_149462# 0.352467f
C909 a_n158_n91786# a_n158_n93222# 0.010536f
C910 a_n158_57558# a_100_57558# 0.328443f
C911 a_n100_57461# a_n100_56025# 0.205388f
C912 w_n358_n183987# a_100_179618# 0.352467f
C913 a_n100_155109# a_n100_153673# 0.205388f
C914 w_n358_n183987# a_n100_n28699# 0.269531f
C915 w_n358_n183987# a_100_n170766# 0.352467f
C916 w_n358_n183987# a_100_94894# 0.352467f
C917 a_n100_163725# a_100_163822# 0.133664f
C918 a_n158_n119070# a_n158_n120506# 0.010536f
C919 a_n158_146590# a_n158_145154# 0.010536f
C920 a_n158_30274# a_100_30274# 0.328443f
C921 a_n100_30177# a_n100_28741# 0.205388f
C922 w_n358_n183987# a_n100_n83267# 0.269531f
C923 a_100_n2754# a_100_n4190# 0.010536f
C924 a_n100_n4287# a_n158_n4190# 0.133664f
C925 w_n358_n183987# a_100_40326# 0.352467f
C926 a_n158_n146354# a_n158_n147790# 0.010536f
C927 a_n158_119306# a_n158_117870# 0.010536f
C928 a_100_n30038# a_100_n31474# 0.010536f
C929 a_n100_n31571# a_n158_n31474# 0.133664f
C930 w_n358_n183987# a_n100_n137835# 0.269531f
C931 w_n358_n183987# a_n100_127825# 0.269531f
C932 w_n358_n183987# a_n158_n48706# 0.352467f
C933 w_n358_n183987# a_100_163822# 0.352467f
C934 a_n158_178182# a_n158_176746# 0.010536f
C935 a_n158_n173638# a_n158_n175074# 0.010536f
C936 a_n158_92022# a_n158_90586# 0.010536f
C937 w_n358_n183987# a_n100_73257# 0.269531f
C938 a_100_n57322# a_100_n58758# 0.010536f
C939 a_n100_n58855# a_n158_n58758# 0.133664f
C940 a_n100_2893# a_n100_1457# 0.205388f
C941 w_n358_n183987# a_n158_n103274# 0.352467f
C942 a_n100_n14339# a_100_n14242# 0.133664f
C943 a_n158_64738# a_n158_63302# 0.010536f
C944 w_n358_n183987# a_n100_18689# 0.269531f
C945 a_100_n84606# a_100_n86042# 0.010536f
C946 a_n100_n86139# a_n158_n86042# 0.133664f
C947 w_n358_n183987# a_100_n14242# 0.352467f
C948 w_n358_n183987# a_n158_107818# 0.352467f
C949 w_n358_n183987# a_n158_n157842# 0.352467f
C950 a_n100_n41623# a_100_n41526# 0.133664f
C951 a_n158_37454# a_n158_36018# 0.010536f
C952 a_100_165258# a_100_166694# 0.010536f
C953 a_100_n111890# a_100_n113326# 0.010536f
C954 a_n100_n113423# a_n158_n113326# 0.133664f
C955 a_100_153770# a_100_152334# 0.010536f
C956 a_n100_152237# a_n158_152334# 0.133664f
C957 w_n358_n183987# a_100_n68810# 0.352467f
C958 w_n358_n183987# a_n158_53250# 0.352467f
C959 a_n100_n68907# a_100_n68810# 0.133664f
C960 a_n158_10170# a_n158_8734# 0.010536f
C961 a_100_n139174# a_100_n140610# 0.010536f
C962 a_n100_n140707# a_n158_n140610# 0.133664f
C963 a_100_126486# a_100_125050# 0.010536f
C964 a_n100_124953# a_n158_125050# 0.133664f
C965 w_n358_n183987# a_100_142282# 0.352467f
C966 a_n158_n24294# a_100_n24294# 0.328443f
C967 a_n100_n24391# a_n100_n25827# 0.205388f
C968 w_n358_n183987# a_100_n123378# 0.352467f
C969 w_n358_n183987# a_n100_n35879# 0.269531f
C970 a_n100_n96191# a_100_n96094# 0.133664f
C971 a_100_118# a_100_n1318# 0.010536f
C972 a_100_99202# a_100_97766# 0.010536f
C973 a_n100_97669# a_n158_97766# 0.133664f
C974 w_n358_n183987# a_n158_166694# 0.352467f
C975 a_100_n166458# a_100_n167894# 0.010536f
C976 a_n100_n167991# a_n158_n167894# 0.133664f
C977 w_n358_n183987# a_100_87714# 0.352467f
C978 a_n158_n51578# a_100_n51578# 0.328443f
C979 a_n100_n51675# a_n100_n53111# 0.205388f
C980 a_n158_160950# a_n158_159514# 0.010536f
C981 w_n358_n183987# a_100_n177946# 0.352467f
C982 w_n358_n183987# a_n100_n90447# 0.269531f
C983 a_n100_n123475# a_100_n123378# 0.133664f
C984 a_n100_142185# a_100_142282# 0.133664f
C985 a_100_71918# a_100_70482# 0.010536f
C986 a_n100_70385# a_n158_70482# 0.133664f
C987 w_n358_n183987# a_n158_n1318# 0.352467f
C988 w_n358_n183987# a_100_33146# 0.352467f
C989 a_n158_n78862# a_100_n78862# 0.328443f
C990 a_n100_n78959# a_n100_n80395# 0.205388f
C991 a_n100_114901# a_100_114998# 0.133664f
C992 w_n358_n183987# a_n100_120645# 0.269531f
C993 w_n358_n183987# a_n100_n145015# 0.269531f
C994 a_n100_n150759# a_100_n150662# 0.133664f
C995 a_100_44634# a_100_43198# 0.010536f
C996 a_n100_43101# a_n158_43198# 0.133664f
C997 a_n158_n106146# a_100_n106146# 0.328443f
C998 a_n100_n106243# a_n100_n107679# 0.205388f
C999 w_n358_n183987# a_n158_n55886# 0.352467f
C1000 a_n100_n178043# a_100_n177946# 0.133664f
C1001 a_n100_87617# a_100_87714# 0.133664f
C1002 w_n358_n183987# a_n100_66077# 0.269531f
C1003 a_n158_132230# a_100_132230# 0.328443f
C1004 a_n100_132133# a_n100_130697# 0.205388f
C1005 a_100_17350# a_100_15914# 0.010536f
C1006 a_n100_15817# a_n158_15914# 0.133664f
C1007 a_n158_n133430# a_100_n133430# 0.328443f
C1008 a_n100_n133527# a_n100_n134963# 0.205388f
C1009 w_n358_n183987# a_n158_155206# 0.352467f
C1010 a_n158_n17114# a_n158_n18550# 0.010536f
C1011 w_n358_n183987# a_n158_n110454# 0.352467f
C1012 a_n100_60333# a_100_60430# 0.133664f
C1013 w_n358_n183987# a_n100_11509# 0.269531f
C1014 w_n358_n183987# a_100_n21422# 0.352467f
C1015 a_n100_7201# a_n100_5765# 0.205388f
C1016 a_n158_n160714# a_100_n160714# 0.328443f
C1017 a_n100_n160811# a_n100_n162247# 0.205388f
C1018 a_n158_104946# a_100_104946# 0.328443f
C1019 a_n100_104849# a_n100_103413# 0.205388f
C1020 w_n358_n183987# a_n158_100638# 0.352467f
C1021 a_n158_n44398# a_n158_n45834# 0.010536f
C1022 w_n358_n183987# a_n158_n165022# 0.352467f
C1023 a_n100_33049# a_100_33146# 0.133664f
C1024 w_n358_n183987# a_100_n75990# 0.352467f
C1025 a_n158_77662# a_100_77662# 0.328443f
C1026 a_n100_77565# a_n100_76129# 0.205388f
C1027 w_n358_n183987# a_n158_46070# 0.352467f
C1028 a_n158_n71682# a_n158_n73118# 0.010536f
C1029 w_n358_n183987# a_100_135102# 0.352467f
C1030 w_n358_n183987# a_100_n130558# 0.352467f
C1031 a_n158_50378# a_100_50378# 0.328443f
C1032 a_n100_50281# a_n100_48845# 0.205388f
C1033 w_n358_n183987# a_n100_n43059# 0.269531f
C1034 a_n158_n98966# a_n158_n100402# 0.010536f
C1035 w_n358_n183987# a_100_80534# 0.352467f
C1036 a_n158_23094# a_100_23094# 0.328443f
C1037 a_n100_22997# a_n100_21561# 0.205388f
C1038 a_n158_n126250# a_n158_n127686# 0.010536f
C1039 a_n158_139410# a_n158_137974# 0.010536f
C1040 w_n358_n183987# a_100_173874# 0.352467f
C1041 a_100_n9934# a_100_n11370# 0.010536f
C1042 a_n100_n11467# a_n158_n11370# 0.133664f
C1043 w_n358_n183987# a_n100_n97627# 0.269531f
C1044 w_n358_n183987# a_100_25966# 0.352467f
C1045 w_n358_n183987# a_n158_n8498# 0.352467f
C1046 a_n158_n153534# a_n158_n154970# 0.010536f
C1047 a_n158_112126# a_n158_110690# 0.010536f
C1048 w_n358_n183987# a_n100_1457# 0.269531f
C1049 w_n358_n183987# a_n100_113465# 0.269531f
C1050 a_100_n37218# a_100_n38654# 0.010536f
C1051 a_n100_n38751# a_n158_n38654# 0.133664f
C1052 w_n358_n183987# a_n100_n152195# 0.269531f
C1053 a_100_175310# a_100_173874# 0.010536f
C1054 a_n100_173777# a_n158_173874# 0.133664f
C1055 a_n100_4329# a_n158_4426# 0.133664f
C1056 w_n358_n183987# a_n158_n63066# 0.352467f
C1057 a_n158_n180818# a_n158_n182254# 0.010536f
C1058 a_n158_84842# a_n158_83406# 0.010536f
C1059 w_n358_n183987# a_n100_58897# 0.269531f
C1060 a_100_n64502# a_100_n65938# 0.010536f
C1061 a_n100_n66035# a_n158_n65938# 0.133664f
C1062 w_n358_n183987# a_n158_148026# 0.352467f
C1063 w_n358_n183987# a_n158_n117634# 0.352467f
C1064 a_n158_57558# a_n158_56122# 0.010536f
C1065 a_n100_n21519# a_100_n21422# 0.133664f
C1066 a_100_n91786# a_100_n93222# 0.010536f
C1067 a_n100_n93319# a_n158_n93222# 0.133664f
C1068 w_n358_n183987# a_100_n28602# 0.352467f
C1069 w_n358_n183987# a_n158_n172202# 0.352467f
C1070 w_n358_n183987# a_n158_93458# 0.352467f
C1071 a_n158_30274# a_n158_28838# 0.010536f
C1072 a_n100_n48803# a_100_n48706# 0.133664f
C1073 a_100_n119070# a_100_n120506# 0.010536f
C1074 a_n100_n120603# a_n158_n120506# 0.133664f
C1075 a_100_146590# a_100_145154# 0.010536f
C1076 a_n100_145057# a_n158_145154# 0.133664f
C1077 w_n358_n183987# a_100_n83170# 0.352467f
C1078 a_n158_n4190# a_100_n4190# 0.328443f
C1079 a_n100_n4287# a_n100_n5723# 0.205388f
C1080 w_n358_n183987# a_n158_38890# 0.352467f
C1081 a_n100_n76087# a_100_n75990# 0.133664f
C1082 a_100_n146354# a_100_n147790# 0.010536f
C1083 a_n100_n147887# a_n158_n147790# 0.133664f
C1084 a_100_119306# a_100_117870# 0.010536f
C1085 a_n100_117773# a_n158_117870# 0.133664f
C1086 w_n358_n183987# a_100_n137738# 0.352467f
C1087 w_n358_n183987# a_100_127922# 0.352467f
C1088 a_n158_n31474# a_100_n31474# 0.328443f
C1089 a_n100_n31571# a_n100_n33007# 0.205388f
C1090 w_n358_n183987# a_n158_162386# 0.352467f
C1091 a_n100_n103371# a_100_n103274# 0.133664f
C1092 a_n100_176649# a_n158_176746# 0.133664f
C1093 w_n358_n183987# a_n100_n50239# 0.269531f
C1094 a_100_n173638# a_100_n175074# 0.010536f
C1095 a_n100_n175171# a_n158_n175074# 0.133664f
C1096 a_100_92022# a_100_90586# 0.010536f
C1097 a_n100_90489# a_n158_90586# 0.133664f
C1098 a_n158_n58758# a_100_n58758# 0.328443f
C1099 a_n100_n58855# a_n100_n60291# 0.205388f
C1100 w_n358_n183987# a_100_73354# 0.352467f
C1101 w_n358_n183987# a_n100_n104807# 0.269531f
C1102 a_n100_n130655# a_100_n130558# 0.133664f
C1103 a_n100_135005# a_100_135102# 0.133664f
C1104 a_n158_2990# a_n158_1554# 0.010536f
C1105 a_100_64738# a_100_63302# 0.010536f
C1106 a_n100_63205# a_n158_63302# 0.133664f
C1107 w_n358_n183987# a_n158_n15678# 0.352467f
C1108 w_n358_n183987# a_100_18786# 0.352467f
C1109 a_n158_n86042# a_100_n86042# 0.328443f
C1110 a_n100_n86139# a_n100_n87575# 0.205388f
C1111 w_n358_n183987# a_n100_n159375# 0.269531f
C1112 a_n100_n157939# a_100_n157842# 0.133664f
C1113 a_n100_107721# a_100_107818# 0.133664f
C1114 w_n358_n183987# a_n100_106285# 0.269531f
C1115 a_100_37454# a_100_36018# 0.010536f
C1116 a_n100_35921# a_n158_36018# 0.133664f
C1117 w_n358_n183987# a_n158_n70246# 0.352467f
C1118 a_n158_n113326# a_100_n113326# 0.328443f
C1119 a_n100_n113423# a_n100_n114859# 0.205388f
C1120 a_n158_152334# a_100_152334# 0.328443f
C1121 a_n100_152237# a_n100_150801# 0.205388f
C1122 w_n358_n183987# a_n100_51717# 0.269531f
C1123 a_n100_80437# a_100_80534# 0.133664f
C1124 a_100_10170# a_100_8734# 0.010536f
C1125 a_n100_8637# a_n158_8734# 0.133664f
C1126 w_n358_n183987# a_n158_n124814# 0.352467f
C1127 a_n158_n140610# a_100_n140610# 0.328443f
C1128 a_n100_n140707# a_n100_n142143# 0.205388f
C1129 a_100_182490# a_n158_182490# 0.328443f
C1130 a_n158_125050# a_100_125050# 0.328443f
C1131 a_n100_124953# a_n100_123517# 0.205388f
C1132 a_n158_n24294# a_n158_n25730# 0.010536f
C1133 w_n358_n183987# a_n158_140846# 0.352467f
C1134 a_n100_53153# a_100_53250# 0.133664f
C1135 w_n358_n183987# a_100_n35782# 0.352467f
C1136 a_n158_n167894# a_100_n167894# 0.328443f
C1137 a_n100_n167991# a_n100_n169427# 0.205388f
C1138 a_n158_97766# a_100_97766# 0.328443f
C1139 a_n100_97669# a_n100_96233# 0.205388f
C1140 w_n358_n183987# a_n158_86278# 0.352467f
C1141 a_n158_n51578# a_n158_n53014# 0.010536f
C1142 a_100_160950# a_100_159514# 0.010536f
C1143 a_n100_159417# a_n158_159514# 0.133664f
C1144 w_n358_n183987# a_n158_n179382# 0.352467f
C1145 a_n100_25869# a_100_25966# 0.133664f
C1146 w_n358_n183987# a_100_n90350# 0.352467f
C1147 a_n158_70482# a_100_70482# 0.328443f
C1148 a_n100_70385# a_n100_68949# 0.205388f
C1149 w_n358_n183987# a_n100_n2851# 0.269531f
C1150 w_n358_n183987# a_n158_31710# 0.352467f
C1151 a_n158_n78862# a_n158_n80298# 0.010536f
C1152 w_n358_n183987# a_100_120742# 0.352467f
C1153 w_n358_n183987# a_100_n144918# 0.352467f
C1154 a_n158_43198# a_100_43198# 0.328443f
C1155 a_n100_43101# a_n100_41665# 0.205388f
C1156 w_n358_n183987# a_n100_n57419# 0.269531f
C1157 a_n158_n106146# a_n158_n107582# 0.010536f
C1158 a_n100_166597# a_100_166694# 0.133664f
C1159 w_n358_n183987# a_100_66174# 0.352467f
C1160 a_n158_15914# a_100_15914# 0.328443f
C1161 a_n100_15817# a_n100_14381# 0.205388f
C1162 a_100_176746# a_100_178182# 0.010536f
C1163 w_n358_n183987# a_n100_n111987# 0.269531f
C1164 a_n158_n133430# a_n158_n134866# 0.010536f
C1165 a_n158_132230# a_n158_130794# 0.010536f
C1166 w_n358_n183987# a_n100_153673# 0.269531f
C1167 a_100_n17114# a_100_n18550# 0.010536f
C1168 a_n100_n18647# a_n158_n18550# 0.133664f
C1169 w_n358_n183987# a_n158_5862# 0.352467f
C1170 w_n358_n183987# a_100_11606# 0.352467f
C1171 w_n358_n183987# a_n158_n22858# 0.352467f
C1172 a_n158_7298# a_n158_5862# 0.010536f
C1173 a_n158_104946# a_n158_103510# 0.010536f
C1174 w_n358_n183987# a_n100_n166555# 0.269531f
C1175 a_n158_n160714# a_n158_n162150# 0.010536f
C1176 w_n358_n183987# a_n100_99105# 0.269531f
C1177 a_100_n44398# a_100_n45834# 0.010536f
C1178 a_n100_n45931# a_n158_n45834# 0.133664f
C1179 a_n100_n1415# a_100_n1318# 0.133664f
C1180 w_n358_n183987# a_n158_n77426# 0.352467f
C1181 a_n158_77662# a_n158_76226# 0.010536f
C1182 w_n358_n183987# a_n100_44537# 0.269531f
C1183 a_100_n71682# a_100_n73118# 0.010536f
C1184 a_n100_n73215# a_n158_n73118# 0.133664f
C1185 w_n358_n183987# a_n158_133666# 0.352467f
C1186 a_n100_n28699# a_100_n28602# 0.133664f
C1187 w_n358_n183987# a_n158_n131994# 0.352467f
C1188 a_n158_50378# a_n158_48942# 0.010536f
C1189 w_n358_n183987# a_100_n42962# 0.352467f
C1190 a_100_n98966# a_100_n100402# 0.010536f
C1191 a_n100_n100499# a_n158_n100402# 0.133664f
C1192 w_n358_n183987# a_n158_79098# 0.352467f
C1193 a_n158_23094# a_n158_21658# 0.010536f
C1194 a_n100_n55983# a_100_n55886# 0.133664f
C1195 a_100_139410# a_100_137974# 0.010536f
C1196 a_n100_137877# a_n158_137974# 0.133664f
C1197 w_n358_n183987# a_100_n97530# 0.352467f
C1198 a_100_n126250# a_100_n127686# 0.010536f
C1199 a_n100_n127783# a_n158_n127686# 0.133664f
C1200 w_n358_n183987# a_n158_172438# 0.352467f
C1201 a_n158_n11370# a_100_n11370# 0.328443f
C1202 a_n100_n11467# a_n100_n12903# 0.205388f
C1203 w_n358_n183987# a_n158_24530# 0.352467f
C1204 w_n358_n183987# a_n100_n10031# 0.269531f
C1205 a_n100_n83267# a_100_n83170# 0.133664f
C1206 a_100_n153534# a_100_n154970# 0.010536f
C1207 a_n100_n155067# a_n158_n154970# 0.133664f
C1208 a_100_112126# a_100_110690# 0.010536f
C1209 a_n100_110593# a_n158_110690# 0.133664f
C1210 w_n358_n183987# a_100_n152098# 0.352467f
C1211 w_n358_n183987# a_100_1554# 0.352467f
C1212 w_n358_n183987# a_100_113562# 0.352467f
C1213 a_n158_n38654# a_100_n38654# 0.328443f
C1214 a_n100_n38751# a_n100_n40187# 0.205388f
C1215 a_n100_173777# a_n100_172341# 0.205388f
C1216 a_n158_4426# a_100_4426# 0.328443f
C1217 w_n358_n183987# a_n100_n64599# 0.269531f
C1218 a_n100_n110551# a_100_n110454# 0.133664f
C1219 a_100_n180818# a_100_n182254# 0.010536f
C1220 a_n100_n182351# a_n158_n182254# 0.133664f
C1221 a_100_84842# a_100_83406# 0.010536f
C1222 a_n100_83309# a_n158_83406# 0.133664f
C1223 w_n358_n183987# a_100_58994# 0.352467f
C1224 a_n158_n65938# a_100_n65938# 0.328443f
C1225 a_n100_n66035# a_n100_n67471# 0.205388f
C1226 a_n100_n137835# a_100_n137738# 0.133664f
C1227 a_n100_127825# a_100_127922# 0.133664f
C1228 w_n358_n183987# a_n100_146493# 0.269531f
C1229 w_n358_n183987# a_n100_n119167# 0.269531f
C1230 a_100_57558# a_100_56122# 0.010536f
C1231 a_n100_56025# a_n158_56122# 0.133664f
C1232 w_n358_n183987# a_n158_n30038# 0.352467f
C1233 a_n158_n93222# a_100_n93222# 0.328443f
C1234 a_n100_n93319# a_n100_n94755# 0.205388f
C1235 a_n100_n165119# a_100_n165022# 0.133664f
C1236 a_n100_100541# a_100_100638# 0.133664f
C1237 w_n358_n183987# a_n100_91925# 0.269531f
C1238 w_n358_n183987# a_n100_n173735# 0.269531f
C1239 a_100_30274# a_100_28838# 0.010536f
C1240 a_n100_28741# a_n158_28838# 0.133664f
C1241 a_n158_n120506# a_100_n120506# 0.328443f
C1242 a_n100_n120603# a_n100_n122039# 0.205388f
C1243 a_n158_145154# a_100_145154# 0.328443f
C1244 a_n100_145057# a_n100_143621# 0.205388f
C1245 w_n358_n183987# a_n158_n84606# 0.352467f
C1246 a_n158_n4190# a_n158_n5626# 0.010536f
C1247 a_n100_73257# a_100_73354# 0.133664f
C1248 w_n358_n183987# a_n100_37357# 0.269531f
C1249 a_n158_n147790# a_100_n147790# 0.328443f
C1250 a_n100_n147887# a_n100_n149323# 0.205388f
C1251 a_n158_117870# a_100_117870# 0.328443f
C1252 a_n100_117773# a_n100_116337# 0.205388f
C1253 w_n358_n183987# a_n158_n139174# 0.352467f
C1254 w_n358_n183987# a_n158_126486# 0.352467f
C1255 a_n158_n31474# a_n158_n32910# 0.010536f
C1256 a_n100_45973# a_100_46070# 0.133664f
C1257 a_100_171002# a_100_169566# 0.010536f
C1258 a_n100_169469# a_n158_169566# 0.133664f
C1259 w_n358_n183987# a_100_n50142# 0.352467f
C1260 w_n358_n183987# a_n100_160853# 0.269531f
C1261 a_n158_n175074# a_100_n175074# 0.328443f
C1262 a_n100_n175171# a_n100_n176607# 0.205388f
C1263 a_n158_90586# a_100_90586# 0.328443f
C1264 a_n100_90489# a_n100_89053# 0.205388f
C1265 w_n358_n183987# a_n158_71918# 0.352467f
C1266 a_n158_n58758# a_n158_n60194# 0.010536f
C1267 a_n100_18689# a_100_18786# 0.133664f
C1268 a_100_2990# a_100_1554# 0.010536f
C1269 w_n358_n183987# a_100_n104710# 0.352467f
C1270 a_n158_63302# a_100_63302# 0.328443f
C1271 a_n100_63205# a_n100_61769# 0.205388f
C1272 a_n158_n86042# a_n158_n87478# 0.010536f
C1273 w_n358_n183987# a_n100_n17211# 0.269531f
C1274 w_n358_n183987# a_n158_17350# 0.352467f
C1275 w_n358_n183987# a_100_n159278# 0.352467f
C1276 w_n358_n183987# a_100_106382# 0.352467f
C1277 a_n158_36018# a_100_36018# 0.328443f
C1278 a_n100_35921# a_n100_34485# 0.205388f
C1279 w_n358_n183987# a_n100_n71779# 0.269531f
C1280 a_n158_n113326# a_n158_n114762# 0.010536f
C1281 a_n158_152334# a_n158_150898# 0.010536f
C1282 w_n358_n183987# a_100_51814# 0.352467f
C1283 a_n158_181054# a_n158_182490# 0.010536f
C1284 a_n158_8734# a_100_8734# 0.328443f
C1285 w_n358_n183987# a_n100_n126347# 0.269531f
C1286 a_n158_n140610# a_n158_n142046# 0.010536f
C1287 a_n158_125050# a_n158_123614# 0.010536f
C1288 w_n358_n183987# a_n100_139313# 0.269531f
C1289 a_100_n24294# a_100_n25730# 0.010536f
C1290 a_n100_n25827# a_n158_n25730# 0.133664f
C1291 w_n358_n183987# a_n158_n37218# 0.352467f
C1292 w_n358_n183987# a_n100_n180915# 0.269531f
C1293 a_n158_n167894# a_n158_n169330# 0.010536f
C1294 a_n158_97766# a_n158_96330# 0.010536f
C1295 a_100_n51578# a_100_n53014# 0.010536f
C1296 a_n100_n53111# a_n158_n53014# 0.133664f
C1297 a_n158_159514# a_100_159514# 0.328443f
C1298 w_n358_n183987# a_n100_84745# 0.269531f
C1299 w_n358_n183987# a_n158_n91786# 0.352467f
C1300 a_n100_n8595# a_100_n8498# 0.133664f
C1301 a_n158_70482# a_n158_69046# 0.010536f
C1302 w_n358_n183987# a_100_n2754# 0.352467f
C1303 w_n358_n183987# a_n100_30177# 0.269531f
C1304 a_100_n78862# a_100_n80298# 0.010536f
C1305 a_n100_n80395# a_n158_n80298# 0.133664f
C1306 a_n100_n35879# a_100_n35782# 0.133664f
C1307 w_n358_n183987# a_n158_n146354# 0.352467f
C1308 w_n358_n183987# a_n158_119306# 0.352467f
C1309 a_n158_43198# a_n158_41762# 0.010536f
C1310 w_n358_n183987# a_n158_178182# 0.352467f
C1311 w_n358_n183987# a_100_n57322# 0.352467f
C1312 a_100_n106146# a_100_n107582# 0.010536f
C1313 a_n100_n107679# a_n158_n107582# 0.133664f
C1314 w_n358_n183987# a_n158_64738# 0.352467f
C1315 a_n100_n63163# a_100_n63066# 0.133664f
C1316 a_n158_15914# a_n158_14478# 0.010536f
C1317 a_100_176746# a_n158_176746# 0.328443f
C1318 a_n100_175213# a_n100_176649# 0.205388f
C1319 w_n358_n183987# a_100_n111890# 0.352467f
C1320 a_100_n133430# a_100_n134866# 0.010536f
C1321 a_n100_n134963# a_n158_n134866# 0.133664f
C1322 a_100_132230# a_100_130794# 0.010536f
C1323 a_n100_130697# a_n158_130794# 0.133664f
C1324 a_n158_n18550# a_100_n18550# 0.328443f
C1325 a_n100_n18647# a_n100_n20083# 0.205388f
C1326 w_n358_n183987# a_100_153770# 0.352467f
C1327 w_n358_n183987# a_n158_10170# 0.352467f
C1328 a_n100_n90447# a_100_n90350# 0.133664f
C1329 w_n358_n183987# a_n100_n24391# 0.269531f
C1330 a_100_7298# a_100_5862# 0.010536f
C1331 w_n358_n183987# a_100_n166458# 0.352467f
C1332 a_100_n160714# a_100_n162150# 0.010536f
C1333 a_n100_n162247# a_n158_n162150# 0.133664f
C1334 a_100_104946# a_100_103510# 0.010536f
C1335 a_n100_103413# a_n158_103510# 0.133664f
C1336 w_n358_n183987# a_100_99202# 0.352467f
C1337 a_n158_n45834# a_100_n45834# 0.328443f
C1338 a_n100_n45931# a_n100_n47367# 0.205388f
C1339 w_n358_n183987# a_n100_n78959# 0.269531f
C1340 a_n100_n117731# a_100_n117634# 0.133664f
C1341 a_n100_147929# a_100_148026# 0.133664f
C1342 a_n100_180957# a_n158_181054# 0.133664f
C1343 a_100_77662# a_100_76226# 0.010536f
C1344 a_n100_76129# a_n158_76226# 0.133664f
C1345 w_n358_n183987# a_100_44634# 0.352467f
C1346 a_n158_n73118# a_100_n73118# 0.328443f
C1347 a_n100_n73215# a_n100_n74651# 0.205388f
C1348 w_n358_n183987# a_n100_132133# 0.269531f
C1349 w_n358_n183987# a_n100_n133527# 0.269531f
C1350 a_n100_n145015# a_100_n144918# 0.133664f
C1351 a_n100_120645# a_100_120742# 0.133664f
C1352 a_100_50378# a_100_48942# 0.010536f
C1353 a_n100_48845# a_n158_48942# 0.133664f
C1354 w_n358_n183987# a_n158_n44398# 0.352467f
C1355 a_n158_n100402# a_100_n100402# 0.328443f
C1356 a_n100_n100499# a_n100_n101935# 0.205388f
C1357 a_n100_93361# a_100_93458# 0.133664f
C1358 w_n358_n183987# a_n100_77565# 0.269531f
C1359 a_n100_n172299# a_100_n172202# 0.133664f
C1360 a_100_23094# a_100_21658# 0.010536f
C1361 a_n100_21561# a_n158_21658# 0.133664f
C1362 w_n358_n183987# a_n158_n98966# 0.352467f
C1363 a_n158_n127686# a_100_n127686# 0.328443f
C1364 a_n100_n127783# a_n100_n129219# 0.205388f
C1365 a_n158_137974# a_100_137974# 0.328443f
C1366 a_n100_137877# a_n100_136441# 0.205388f
C1367 w_n358_n183987# a_n100_170905# 0.269531f
C1368 a_n158_n11370# a_n158_n12806# 0.010536f
C1369 a_n100_66077# a_100_66174# 0.133664f
C1370 w_n358_n183987# a_n100_22997# 0.269531f
C1371 w_n358_n183987# a_100_n9934# 0.352467f
C1372 a_n158_110690# a_100_110690# 0.328443f
C1373 a_n100_110593# a_n100_109157# 0.205388f
C1374 w_n358_n183987# a_n158_n153534# 0.352467f
C1375 a_n158_n154970# a_100_n154970# 0.328443f
C1376 a_n100_n155067# a_n100_n156503# 0.205388f
C1377 w_n358_n183987# a_n158_112126# 0.352467f
C1378 a_n158_n38654# a_n158_n40090# 0.010536f
C1379 a_n100_38793# a_100_38890# 0.133664f
C1380 w_n358_n183987# a_100_n64502# 0.352467f
C1381 a_n158_n182254# a_100_n182254# 0.328443f
C1382 a_n100_n182351# a_n100_n183787# 0.205388f
C1383 a_n158_83406# a_100_83406# 0.328443f
C1384 a_n100_83309# a_n100_81873# 0.205388f
C1385 w_n358_n183987# a_n158_57558# 0.352467f
C1386 a_n158_n65938# a_n158_n67374# 0.010536f
C1387 a_n100_11509# a_100_11606# 0.133664f
C1388 w_n358_n183987# a_100_146590# 0.352467f
C1389 w_n358_n183987# a_100_n119070# 0.352467f
C1390 a_n158_56122# a_100_56122# 0.328443f
C1391 a_n100_56025# a_n100_54589# 0.205388f
C1392 w_n358_n183987# a_n100_n31571# 0.269531f
C1393 a_n158_n93222# a_n158_n94658# 0.010536f
C1394 w_n358_n183987# a_100_92022# 0.352467f
C1395 w_n358_n183987# a_100_n173638# 0.352467f
C1396 a_n158_28838# a_100_28838# 0.328443f
C1397 a_n100_28741# a_n100_27305# 0.205388f
C1398 a_n100_162289# a_100_162386# 0.133664f
C1399 a_n158_145154# a_n158_143718# 0.010536f
C1400 w_n358_n183987# a_n100_n86139# 0.269531f
C1401 a_n158_n120506# a_n158_n121942# 0.010536f
C1402 a_100_n4190# a_100_n5626# 0.010536f
C1403 a_n100_n5723# a_n158_n5626# 0.133664f
C1404 w_n358_n183987# a_100_37454# 0.352467f
C1405 a_n158_n147790# a_n158_n149226# 0.010536f
C1406 a_n158_117870# a_n158_116434# 0.010536f
C1407 w_n358_n183987# a_n100_124953# 0.269531f
C1408 w_n358_n183987# a_n100_n140707# 0.269531f
C1409 a_100_n31474# a_100_n32910# 0.010536f
C1410 a_n100_n33007# a_n158_n32910# 0.133664f
C1411 a_100_182490# a_n100_182393# 0.133664f
C1412 a_n158_169566# a_100_169566# 0.328443f
C1413 a_n100_169469# a_n100_168033# 0.205388f
C1414 w_n358_n183987# a_n158_n51578# 0.352467f
C1415 w_n358_n183987# a_100_160950# 0.352467f
C1416 a_n158_n175074# a_n158_n176510# 0.010536f
C1417 a_n158_90586# a_n158_89150# 0.010536f
C1418 w_n358_n183987# a_n100_70385# 0.269531f
C1419 a_100_n58758# a_100_n60194# 0.010536f
C1420 a_n100_n60291# a_n158_n60194# 0.133664f
C1421 w_n358_n183987# a_n100_21# 0.269531f
C1422 a_n100_n15775# a_100_n15678# 0.133664f
C1423 w_n358_n183987# a_n158_n106146# 0.352467f
C1424 a_n158_63302# a_n158_61866# 0.010536f
C1425 w_n358_n183987# a_100_n17114# 0.352467f
C1426 w_n358_n183987# a_n100_15817# 0.269531f
C1427 a_100_n86042# a_100_n87478# 0.010536f
C1428 a_n100_n87575# a_n158_n87478# 0.133664f
C1429 w_n358_n183987# a_n158_104946# 0.352467f
C1430 a_n100_n43059# a_100_n42962# 0.133664f
C1431 w_n358_n183987# a_n158_n160714# 0.352467f
C1432 a_n158_36018# a_n158_34582# 0.010536f
C1433 a_100_n113326# a_100_n114762# 0.010536f
C1434 a_n100_n114859# a_n158_n114762# 0.133664f
C1435 a_100_152334# a_100_150898# 0.010536f
C1436 a_n100_150801# a_n158_150898# 0.133664f
C1437 w_n358_n183987# a_100_n71682# 0.352467f
C1438 w_n358_n183987# a_n158_50378# 0.352467f
C1439 a_n100_n70343# a_100_n70246# 0.133664f
C1440 w_n358_n183987# a_100_n126250# 0.352467f
C1441 a_100_n140610# a_100_n142046# 0.010536f
C1442 a_n100_n142143# a_n158_n142046# 0.133664f
C1443 a_100_125050# a_100_123614# 0.010536f
C1444 a_n100_123517# a_n158_123614# 0.133664f
C1445 w_n358_n183987# a_100_139410# 0.352467f
C1446 a_n158_n25730# a_100_n25730# 0.328443f
C1447 a_n100_n25827# a_n100_n27263# 0.205388f
C1448 a_n100_n97627# a_100_n97530# 0.133664f
C1449 w_n358_n183987# a_n100_n38751# 0.269531f
C1450 w_n358_n183987# a_100_n180818# 0.352467f
C1451 a_100_n167894# a_100_n169330# 0.010536f
C1452 a_n100_n169427# a_n158_n169330# 0.133664f
C1453 a_100_97766# a_100_96330# 0.010536f
C1454 a_n100_96233# a_n158_96330# 0.133664f
C1455 w_n358_n183987# a_100_84842# 0.352467f
C1456 a_n158_n53014# a_100_n53014# 0.328443f
C1457 a_n100_n53111# a_n100_n54547# 0.205388f
C1458 a_n100_n124911# a_100_n124814# 0.133664f
C1459 w_n358_n183987# a_n100_n93319# 0.269531f
C1460 a_n100_140749# a_100_140846# 0.133664f
C1461 a_100_70482# a_100_69046# 0.010536f
C1462 a_n100_68949# a_n158_69046# 0.133664f
C1463 a_n158_n80298# a_100_n80298# 0.328443f
C1464 a_n100_n80395# a_n100_n81831# 0.205388f
C1465 w_n358_n183987# a_n158_n4190# 0.352467f
C1466 w_n358_n183987# a_100_30274# 0.352467f
C1467 a_n100_n152195# a_100_n152098# 0.133664f
C1468 w_n358_n183987# a_n100_n147887# 0.269531f
C1469 a_n100_1457# a_100_1554# 0.133664f
C1470 a_n100_113465# a_100_113562# 0.133664f
C1471 w_n358_n183987# a_n100_117773# 0.269531f
C1472 a_100_43198# a_100_41762# 0.010536f
C1473 a_n100_41665# a_n158_41762# 0.133664f
C1474 w_n358_n183987# a_n100_176649# 0.269531f
C1475 w_n358_n183987# a_n158_n58758# 0.352467f
C1476 a_n158_n107582# a_100_n107582# 0.328443f
C1477 a_n100_n107679# a_n100_n109115# 0.205388f
C1478 a_n100_180957# a_100_181054# 0.133664f
C1479 a_n100_n179479# a_100_n179382# 0.133664f
C1480 a_n100_86181# a_100_86278# 0.133664f
C1481 w_n358_n183987# a_n100_63205# 0.269531f
C1482 a_100_15914# a_100_14478# 0.010536f
C1483 a_n100_14381# a_n158_14478# 0.133664f
C1484 a_n158_159514# a_n158_158078# 0.010536f
C1485 w_n358_n183987# a_n158_n113326# 0.352467f
C1486 a_n158_n134866# a_100_n134866# 0.328443f
C1487 a_n100_n134963# a_n100_n136399# 0.205388f
C1488 a_n158_130794# a_100_130794# 0.328443f
C1489 a_n100_130697# a_n100_129261# 0.205388f
C1490 w_n358_n183987# a_n158_152334# 0.352467f
C1491 a_n158_175310# a_n158_176746# 0.010536f
C1492 a_n158_n18550# a_n158_n19986# 0.010536f
C1493 w_n358_n183987# a_n100_8637# 0.269531f
C1494 a_n100_58897# a_100_58994# 0.133664f
C1495 w_n358_n183987# a_100_n24294# 0.352467f
C1496 w_n358_n183987# a_n158_n167894# 0.352467f
C1497 a_n158_n162150# a_100_n162150# 0.328443f
C1498 a_n100_n162247# a_n100_n163683# 0.205388f
C1499 a_n158_103510# a_100_103510# 0.328443f
C1500 a_n100_103413# a_n100_101977# 0.205388f
C1501 w_n358_n183987# a_n158_97766# 0.352467f
C1502 a_n158_n45834# a_n158_n47270# 0.010536f
C1503 a_n100_165161# a_n158_165258# 0.133664f
C1504 a_n100_31613# a_100_31710# 0.133664f
C1505 w_n358_n183987# a_100_n78862# 0.352467f
C1506 w_n358_n183987# a_n158_43198# 0.352467f
C1507 a_n158_76226# a_100_76226# 0.328443f
C1508 a_n100_76129# a_n100_74693# 0.205388f
C1509 a_n158_n73118# a_n158_n74554# 0.010536f
C1510 w_n358_n183987# a_100_n133430# 0.352467f
C1511 w_n358_n183987# a_100_132230# 0.352467f
C1512 a_n158_48942# a_100_48942# 0.328443f
C1513 a_n100_48845# a_n100_47409# 0.205388f
C1514 w_n358_n183987# a_n100_n45931# 0.269531f
C1515 a_n158_n100402# a_n158_n101838# 0.010536f
C1516 w_n358_n183987# a_100_182490# 0.35701f
C1517 w_n358_n183987# a_100_77662# 0.352467f
C1518 a_n158_21658# a_100_21658# 0.328443f
C1519 a_n100_21561# a_n100_20125# 0.205388f
C1520 w_n358_n183987# a_n100_n100499# 0.269531f
C1521 a_n158_n127686# a_n158_n129122# 0.010536f
C1522 a_n158_137974# a_n158_136538# 0.010536f
C1523 a_100_n11370# a_100_n12806# 0.010536f
C1524 a_n100_n12903# a_n158_n12806# 0.133664f
C1525 w_n358_n183987# a_100_23094# 0.352467f
C1526 w_n358_n183987# a_n158_n11370# 0.352467f
C1527 w_n358_n183987# a_n100_110593# 0.269531f
C1528 w_n358_n183987# a_n100_n155067# 0.269531f
C1529 a_n158_n154970# a_n158_n156406# 0.010536f
C1530 a_n158_110690# a_n158_109254# 0.010536f
C1531 a_100_n38654# a_100_n40090# 0.010536f
C1532 a_n100_n40187# a_n158_n40090# 0.133664f
C1533 w_n358_n183987# a_n158_4426# 0.352467f
C1534 w_n358_n183987# a_n158_n65938# 0.352467f
C1535 a_n158_83406# a_n158_81970# 0.010536f
C1536 w_n358_n183987# a_n100_56025# 0.269531f
C1537 a_n100_5765# a_100_5862# 0.133664f
C1538 a_n158_n182254# a_n158_n183690# 0.010536f
C1539 a_100_n65938# a_100_n67374# 0.010536f
C1540 a_n100_n67471# a_n158_n67374# 0.133664f
C1541 w_n358_n183987# a_n158_145154# 0.352467f
C1542 a_n100_n22955# a_100_n22858# 0.133664f
C1543 w_n358_n183987# a_n158_n120506# 0.352467f
C1544 a_n158_56122# a_n158_54686# 0.010536f
C1545 w_n358_n183987# a_100_n31474# 0.352467f
C1546 a_100_n93222# a_100_n94658# 0.010536f
C1547 a_n100_n94755# a_n158_n94658# 0.133664f
C1548 w_n358_n183987# a_n100_169469# 0.269531f
C1549 w_n358_n183987# a_n158_90586# 0.352467f
C1550 a_n100_n50239# a_100_n50142# 0.133664f
C1551 w_n358_n183987# a_n158_n175074# 0.352467f
C1552 a_n158_28838# a_n158_27402# 0.010536f
C1553 w_n358_n183987# a_100_n86042# 0.352467f
C1554 a_100_n120506# a_100_n121942# 0.010536f
C1555 a_n100_n122039# a_n158_n121942# 0.133664f
C1556 a_100_145154# a_100_143718# 0.010536f
C1557 a_n100_143621# a_n158_143718# 0.133664f
C1558 a_n158_n5626# a_100_n5626# 0.328443f
C1559 a_n100_n5723# a_n100_n7159# 0.205388f
C1560 w_n358_n183987# a_n158_36018# 0.352467f
C1561 a_n100_n77523# a_100_n77426# 0.133664f
C1562 a_100_117870# a_100_116434# 0.010536f
C1563 a_n100_116337# a_n158_116434# 0.133664f
C1564 w_n358_n183987# a_100_125050# 0.352467f
C1565 w_n358_n183987# a_100_n140610# 0.352467f
C1566 a_100_n147790# a_100_n149226# 0.010536f
C1567 a_n100_n149323# a_n158_n149226# 0.133664f
C1568 a_n158_n32910# a_100_n32910# 0.328443f
C1569 a_n100_n33007# a_n100_n34443# 0.205388f
C1570 a_n100_n104807# a_100_n104710# 0.133664f
C1571 a_n158_169566# a_n158_168130# 0.010536f
C1572 w_n358_n183987# a_n100_n53111# 0.269531f
C1573 w_n358_n183987# a_n158_159514# 0.352467f
C1574 a_100_n175074# a_100_n176510# 0.010536f
C1575 a_n100_n176607# a_n158_n176510# 0.133664f
C1576 a_100_90586# a_100_89150# 0.010536f
C1577 a_n100_89053# a_n158_89150# 0.133664f
C1578 w_n358_n183987# a_100_70482# 0.352467f
C1579 a_n158_n60194# a_100_n60194# 0.328443f
C1580 a_n100_n60291# a_n100_n61727# 0.205388f
C1581 a_n100_n132091# a_100_n131994# 0.133664f
C1582 a_n100_133569# a_100_133666# 0.133664f
C1583 w_n358_n183987# a_n100_n107679# 0.269531f
C1584 a_100_63302# a_100_61866# 0.010536f
C1585 a_n100_61769# a_n158_61866# 0.133664f
C1586 w_n358_n183987# a_100_15914# 0.352467f
C1587 w_n358_n183987# a_n158_n18550# 0.352467f
C1588 a_n158_n87478# a_100_n87478# 0.328443f
C1589 a_n100_n87575# a_n100_n89011# 0.205388f
C1590 a_n100_n159375# a_100_n159278# 0.133664f
C1591 a_n100_106285# a_100_106382# 0.133664f
C1592 w_n358_n183987# a_n100_103413# 0.269531f
C1593 w_n358_n183987# a_n100_n162247# 0.269531f
C1594 a_100_36018# a_100_34582# 0.010536f
C1595 a_n100_34485# a_n158_34582# 0.133664f
C1596 a_n158_150898# a_100_150898# 0.328443f
C1597 a_n100_150801# a_n100_149365# 0.205388f
C1598 w_n358_n183987# a_n158_n73118# 0.352467f
C1599 a_n158_n114762# a_100_n114762# 0.328443f
C1600 a_n100_n114859# a_n100_n116295# 0.205388f
C1601 a_n100_79001# a_100_79098# 0.133664f
C1602 w_n358_n183987# a_n100_48845# 0.269531f
C1603 a_n158_n142046# a_100_n142046# 0.328443f
C1604 a_n100_n142143# a_n100_n143579# 0.205388f
C1605 a_n158_123614# a_100_123614# 0.328443f
C1606 a_n100_123517# a_n100_122081# 0.205388f
C1607 w_n358_n183987# a_n158_137974# 0.352467f
C1608 w_n358_n183987# a_n158_n127686# 0.352467f
C1609 a_n158_n25730# a_n158_n27166# 0.010536f
C1610 a_n100_51717# a_100_51814# 0.133664f
C1611 a_n100_172341# a_100_172438# 0.133664f
C1612 w_n358_n183987# a_100_n38654# 0.352467f
C1613 w_n358_n183987# a_n158_n182254# 0.352467f
C1614 a_n158_n169330# a_100_n169330# 0.328443f
C1615 a_n100_n169427# a_n100_n170863# 0.205388f
C1616 a_n158_96330# a_100_96330# 0.328443f
C1617 a_n100_96233# a_n100_94797# 0.205388f
C1618 w_n358_n183987# a_n158_83406# 0.352467f
C1619 a_n158_n53014# a_n158_n54450# 0.010536f
C1620 a_n100_24433# a_100_24530# 0.133664f
C1621 w_n358_n183987# a_100_n93222# 0.352467f
C1622 a_n158_69046# a_100_69046# 0.328443f
C1623 a_n100_68949# a_n100_67513# 0.205388f
C1624 w_n358_n183987# a_n158_28838# 0.352467f
C1625 w_n358_n183987# a_n100_n5723# 0.269531f
C1626 a_n158_n80298# a_n158_n81734# 0.010536f
C1627 w_n358_n183987# a_n158_118# 0.352467f
C1628 w_n358_n183987# a_100_n147790# 0.352467f
C1629 w_n358_n183987# a_100_117870# 0.352467f
C1630 a_n158_41762# a_100_41762# 0.328443f
C1631 a_n100_41665# a_n100_40229# 0.205388f
C1632 a_n158_n107582# a_n158_n109018# 0.010536f
C1633 w_n358_n183987# a_n100_n60291# 0.269531f
C1634 w_n358_n183987# a_100_63302# 0.352467f
C1635 a_n158_14478# a_100_14478# 0.328443f
C1636 a_n100_14381# a_n100_12945# 0.205388f
C1637 w_n358_n183987# a_n100_n114859# 0.269531f
C1638 a_n158_n134866# a_n158_n136302# 0.010536f
C1639 a_n158_130794# a_n158_129358# 0.010536f
C1640 w_n358_n183987# a_n100_150801# 0.269531f
C1641 a_100_n18550# a_100_n19986# 0.010536f
C1642 a_n100_n20083# a_n158_n19986# 0.133664f
C1643 w_n358_n183987# a_100_8734# 0.352467f
C1644 w_n358_n183987# a_n158_n25730# 0.352467f
C1645 w_n358_n183987# a_n100_n169427# 0.269531f
C1646 a_n158_n162150# a_n158_n163586# 0.010536f
C1647 a_n158_103510# a_n158_102074# 0.010536f
C1648 w_n358_n183987# a_n100_96233# 0.269531f
C1649 a_100_n45834# a_100_n47270# 0.010536f
C1650 a_n100_n47367# a_n158_n47270# 0.133664f
C1651 a_n158_165258# a_100_165258# 0.328443f
C1652 a_n100_165161# a_n100_163725# 0.205388f
C1653 w_n358_n183987# a_n158_n80298# 0.352467f
C1654 a_n100_n2851# a_100_n2754# 0.133664f
C1655 a_n158_76226# a_n158_74790# 0.010536f
C1656 w_n358_n183987# a_n100_41665# 0.269531f
C1657 a_100_n73118# a_100_n74554# 0.010536f
C1658 a_n100_n74651# a_n158_n74554# 0.133664f
C1659 a_n100_n30135# a_100_n30038# 0.133664f
C1660 w_n358_n183987# a_n158_n134866# 0.352467f
C1661 w_n358_n183987# a_n158_130794# 0.352467f
C1662 a_n158_48942# a_n158_47506# 0.010536f
C1663 w_n358_n183987# a_100_n45834# 0.352467f
C1664 a_100_n100402# a_100_n101838# 0.010536f
C1665 a_n100_n101935# a_n158_n101838# 0.133664f
C1666 w_n358_n183987# a_n100_165161# 0.269531f
C1667 w_n358_n183987# a_n158_181054# 0.352467f
C1668 a_n100_n57419# a_100_n57322# 0.133664f
C1669 w_n358_n183987# a_n158_76226# 0.352467f
C1670 a_n158_21658# a_n158_20222# 0.010536f
C1671 a_n100_1457# a_n100_21# 0.205388f
C1672 w_n358_n183987# a_100_n100402# 0.352467f
C1673 a_100_n127686# a_100_n129122# 0.010536f
C1674 a_n100_n129219# a_n158_n129122# 0.133664f
C1675 a_100_137974# a_100_136538# 0.010536f
C1676 a_n100_136441# a_n158_136538# 0.133664f
C1677 a_n158_n12806# a_100_n12806# 0.328443f
C1678 a_n100_n12903# a_n100_n14339# 0.205388f
C1679 w_n358_n183987# a_n158_21658# 0.352467f
C1680 a_n100_n84703# a_100_n84606# 0.133664f
C1681 w_n358_n183987# a_n100_n12903# 0.269531f
C1682 a_n158_171002# a_100_171002# 0.328443f
C1683 w_n358_n183987# a_100_n154970# 0.352467f
C1684 a_100_n154970# a_100_n156406# 0.010536f
C1685 a_n100_n156503# a_n158_n156406# 0.133664f
C1686 a_100_110690# a_100_109254# 0.010536f
C1687 a_n100_109157# a_n158_109254# 0.133664f
C1688 w_n358_n183987# a_100_110690# 0.352467f
C1689 a_n158_n40090# a_100_n40090# 0.328443f
C1690 a_n100_n40187# a_n100_n41623# 0.205388f
C1691 a_n100_n111987# a_100_n111890# 0.133664f
C1692 w_n358_n183987# a_n100_n67471# 0.269531f
C1693 a_n100_153673# a_100_153770# 0.133664f
C1694 w_n358_n183987# a_100_56122# 0.352467f
C1695 a_100_n182254# a_100_n183690# 0.010536f
C1696 a_n100_n183787# a_n158_n183690# 0.133664f
C1697 a_100_83406# a_100_81970# 0.010536f
C1698 a_n100_81873# a_n158_81970# 0.133664f
C1699 a_n158_n67374# a_100_n67374# 0.328443f
C1700 a_n100_n67471# a_n100_n68907# 0.205388f
C1701 w_n358_n183987# a_100_176746# 0.352467f
C1702 a_n100_n139271# a_100_n139174# 0.133664f
C1703 w_n358_n183987# a_n100_n122039# 0.269531f
C1704 a_n100_126389# a_100_126486# 0.133664f
C1705 w_n358_n183987# a_n100_143621# 0.269531f
C1706 a_100_56122# a_100_54686# 0.010536f
C1707 a_n100_54589# a_n158_54686# 0.133664f
C1708 w_n358_n183987# a_n158_n32910# 0.352467f
C1709 a_n158_n94658# a_100_n94658# 0.328443f
C1710 a_n100_n94755# a_n100_n96191# 0.205388f
C1711 w_n358_n183987# a_100_169566# 0.352467f
C1712 a_n100_175213# a_n158_175310# 0.133664f
C1713 a_n100_n166555# a_100_n166458# 0.133664f
C1714 a_100_176746# a_100_175310# 0.010536f
C1715 w_n358_n183987# a_n100_89053# 0.269531f
C1716 w_n358_n183987# a_n100_n176607# 0.269531f
C1717 a_n100_99105# a_100_99202# 0.133664f
C1718 a_100_28838# a_100_27402# 0.010536f
C1719 a_n100_27305# a_n158_27402# 0.133664f
C1720 w_n358_n183987# a_n158_n87478# 0.352467f
C1721 a_n158_n121942# a_100_n121942# 0.328443f
C1722 a_n100_n122039# a_n100_n123475# 0.205388f
C1723 a_n158_143718# a_100_143718# 0.328443f
C1724 a_n100_143621# a_n100_142185# 0.205388f
C1725 a_n158_n5626# a_n158_n7062# 0.010536f
C1726 a_n100_71821# a_100_71918# 0.133664f
C1727 w_n358_n183987# a_n100_34485# 0.269531f
C1728 w_n358_n183987# a_n158_123614# 0.352467f
C1729 w_n358_n183987# a_n158_n142046# 0.352467f
C1730 a_n158_n149226# a_100_n149226# 0.328443f
C1731 a_n100_n149323# a_n100_n150759# 0.205388f
C1732 a_n158_116434# a_100_116434# 0.328443f
C1733 a_n100_116337# a_n100_114901# 0.205388f
C1734 a_n158_n32910# a_n158_n34346# 0.010536f
C1735 a_n100_44537# a_100_44634# 0.133664f
C1736 w_n358_n183987# a_100_n53014# 0.352467f
C1737 a_100_169566# a_100_168130# 0.010536f
C1738 a_n100_168033# a_n158_168130# 0.133664f
C1739 a_n158_89150# a_100_89150# 0.328443f
C1740 a_n100_89053# a_n100_87617# 0.205388f
C1741 w_n358_n183987# a_n158_69046# 0.352467f
C1742 a_n158_n176510# a_100_n176510# 0.328443f
C1743 a_n100_n176607# a_n100_n178043# 0.205388f
C1744 a_n158_n60194# a_n158_n61630# 0.010536f
C1745 a_n100_17253# a_100_17350# 0.133664f
C1746 w_n358_n183987# a_100_n107582# 0.352467f
C1747 a_n100_5765# a_n100_4329# 0.205388f
C1748 a_n158_61866# a_100_61866# 0.328443f
C1749 a_n100_61769# a_n100_60333# 0.205388f
C1750 w_n358_n183987# a_n158_14478# 0.352467f
C1751 w_n358_n183987# a_n100_n20083# 0.269531f
C1752 a_n158_n87478# a_n158_n88914# 0.010536f
C1753 w_n358_n183987# a_100_103510# 0.352467f
C1754 w_n358_n183987# a_100_n162150# 0.352467f
C1755 a_n158_34582# a_100_34582# 0.328443f
C1756 a_n100_34485# a_n100_33049# 0.205388f
C1757 w_n358_n183987# a_n100_n74651# 0.269531f
C1758 a_n158_n114762# a_n158_n116198# 0.010536f
C1759 a_n158_150898# a_n158_149462# 0.010536f
C1760 w_n358_n183987# a_100_48942# 0.352467f
C1761 a_n158_123614# a_n158_122178# 0.010536f
C1762 w_n358_n183987# a_n100_136441# 0.269531f
C1763 w_n358_n183987# a_n100_n129219# 0.269531f
C1764 a_n158_n142046# a_n158_n143482# 0.010536f
C1765 a_100_n25730# a_100_n27166# 0.010536f
C1766 a_n100_n27263# a_n158_n27166# 0.133664f
C1767 w_n358_n183987# a_n158_n40090# 0.352467f
C1768 a_n158_n169330# a_n158_n170766# 0.010536f
C1769 a_n158_96330# a_n158_94894# 0.010536f
C1770 w_n358_n183987# a_n100_81873# 0.269531f
C1771 w_n358_n183987# a_n100_n183787# 0.349164f
C1772 a_100_n53014# a_100_n54450# 0.010536f
C1773 a_n100_n54547# a_n158_n54450# 0.133664f
C1774 a_n100_n10031# a_100_n9934# 0.133664f
C1775 w_n358_n183987# a_n158_n94658# 0.352467f
C1776 a_n158_69046# a_n158_67610# 0.010536f
C1777 w_n358_n183987# a_n100_27305# 0.269531f
C1778 w_n358_n183987# a_100_n5626# 0.352467f
C1779 a_100_n80298# a_100_n81734# 0.010536f
C1780 a_n100_n81831# a_n158_n81734# 0.133664f
C1781 w_n358_n183987# a_n158_116434# 0.352467f
C1782 a_n100_n37315# a_100_n37218# 0.133664f
C1783 w_n358_n183987# a_n158_n149226# 0.352467f
C1784 a_n100_2893# a_n158_2990# 0.133664f
C1785 a_n158_41762# a_n158_40326# 0.010536f
C1786 w_n358_n183987# a_100_n60194# 0.352467f
C1787 a_100_n107582# a_100_n109018# 0.010536f
C1788 a_n100_n109115# a_n158_n109018# 0.133664f
C1789 w_n358_n183987# a_n158_61866# 0.352467f
C1790 a_n100_n64599# a_100_n64502# 0.133664f
C1791 a_n158_14478# a_n158_13042# 0.010536f
C1792 a_100_n134866# a_100_n136302# 0.010536f
C1793 a_n100_n136399# a_n158_n136302# 0.133664f
C1794 a_100_130794# a_100_129358# 0.010536f
C1795 a_n100_129261# a_n158_129358# 0.133664f
C1796 w_n358_n183987# a_100_150898# 0.352467f
C1797 w_n358_n183987# a_100_n114762# 0.352467f
C1798 a_n158_n19986# a_100_n19986# 0.328443f
C1799 a_n100_n20083# a_n100_n21519# 0.205388f
C1800 a_n100_n91883# a_100_n91786# 0.133664f
C1801 w_n358_n183987# a_n100_n27263# 0.269531f
C1802 w_n358_n183987# a_100_n169330# 0.352467f
C1803 a_100_n162150# a_100_n163586# 0.010536f
C1804 a_n100_n163683# a_n158_n163586# 0.133664f
C1805 a_100_103510# a_100_102074# 0.010536f
C1806 a_n100_101977# a_n158_102074# 0.133664f
C1807 w_n358_n183987# a_100_181054# 0.352467f
C1808 w_n358_n183987# a_100_96330# 0.352467f
C1809 a_n158_165258# a_n158_163822# 0.010536f
C1810 a_n158_n47270# a_100_n47270# 0.328443f
C1811 a_n100_n47367# a_n100_n48803# 0.205388f
C1812 a_n100_n119167# a_100_n119070# 0.133664f
C1813 a_n100_146493# a_100_146590# 0.133664f
C1814 w_n358_n183987# a_n100_n81831# 0.269531f
C1815 a_n158_118# a_n158_n1318# 0.010536f
C1816 a_100_76226# a_100_74790# 0.010536f
C1817 a_n100_74693# a_n158_74790# 0.133664f
C1818 w_n358_n183987# a_100_41762# 0.352467f
C1819 a_n158_n74554# a_100_n74554# 0.328443f
C1820 a_n100_n74651# a_n100_n76087# 0.205388f
C1821 a_n100_n146451# a_100_n146354# 0.133664f
C1822 w_n358_n183987# a_n100_n136399# 0.269531f
C1823 a_n100_119209# a_100_119306# 0.133664f
C1824 w_n358_n183987# a_n100_129261# 0.269531f
C1825 a_100_48942# a_100_47506# 0.010536f
C1826 a_n100_47409# a_n158_47506# 0.133664f
C1827 a_n158_n101838# a_100_n101838# 0.328443f
C1828 a_n100_n101935# a_n100_n103371# 0.205388f
C1829 w_n358_n183987# a_100_165258# 0.352467f
C1830 a_n100_178085# a_100_178182# 0.133664f
C1831 w_n358_n183987# a_n158_n47270# 0.352467f
C1832 a_n100_n173735# a_100_n173638# 0.133664f
C1833 w_n358_n183987# a_100_118# 0.352467f
C1834 a_n100_91925# a_100_92022# 0.133664f
C1835 w_n358_n183987# a_n100_74693# 0.269531f
C1836 a_100_21658# a_100_20222# 0.010536f
C1837 a_n100_20125# a_n158_20222# 0.133664f
C1838 w_n358_n183987# a_n158_n101838# 0.352467f
C1839 a_n158_n129122# a_100_n129122# 0.328443f
C1840 a_n100_n129219# a_n100_n130655# 0.205388f
C1841 a_n158_136538# a_100_136538# 0.328443f
C1842 a_n100_136441# a_n100_135005# 0.205388f
C1843 a_n158_n12806# a_n158_n14242# 0.010536f
C1844 a_n100_64641# a_100_64738# 0.133664f
C1845 w_n358_n183987# a_n100_20125# 0.269531f
C1846 a_n158_171002# a_n158_169566# 0.010536f
C1847 w_n358_n183987# a_100_n12806# 0.352467f
C1848 w_n358_n183987# a_n158_n156406# 0.352467f
C1849 a_n158_n156406# a_100_n156406# 0.328443f
C1850 a_n100_n156503# a_n100_n157939# 0.205388f
C1851 a_n158_109254# a_100_109254# 0.328443f
C1852 a_n100_109157# a_n100_107721# 0.205388f
C1853 w_n358_n183987# a_n158_109254# 0.352467f
C1854 a_n158_n40090# a_n158_n41526# 0.010536f
C1855 a_n100_37357# a_100_37454# 0.133664f
C1856 w_n358_n183987# a_100_n67374# 0.352467f
C1857 w_n358_n183987# a_n100_7201# 0.269531f
C1858 a_n158_n183690# a_100_n183690# 0.328443f
C1859 a_n158_81970# a_100_81970# 0.328443f
C1860 a_n100_81873# a_n100_80437# 0.205388f
C1861 w_n358_n183987# a_n158_54686# 0.352467f
C1862 a_n158_n67374# a_n158_n68810# 0.010536f
C1863 w_n358_n183987# a_n158_175310# 0.352467f
C1864 a_n100_7201# a_n158_7298# 0.133664f
C1865 a_n100_10073# a_100_10170# 0.133664f
C1866 w_n358_n183987# a_100_n121942# 0.352467f
C1867 w_n358_n183987# a_100_143718# 0.352467f
C1868 a_n158_54686# a_100_54686# 0.328443f
C1869 a_n100_54589# a_n100_53153# 0.205388f
C1870 w_n358_n183987# a_n100_n34443# 0.269531f
C1871 a_n158_n94658# a_n158_n96094# 0.010536f
C1872 w_n358_n183987# a_n158_168130# 0.352467f
C1873 a_n100_175213# a_n100_173777# 0.205388f
C1874 a_n158_175310# a_100_175310# 0.328443f
C1875 a_n100_160853# a_100_160950# 0.133664f
C1876 w_n358_n183987# a_100_n176510# 0.352467f
C1877 w_n358_n183987# a_100_89150# 0.352467f
C1878 a_n158_27402# a_100_27402# 0.328443f
C1879 a_n100_27305# a_n100_25869# 0.205388f
C1880 w_n358_n183987# a_n100_n89011# 0.269531f
C1881 a_n158_n121942# a_n158_n123378# 0.010536f
C1882 a_n158_143718# a_n158_142282# 0.010536f
C1883 a_100_n5626# a_100_n7062# 0.010536f
C1884 a_n100_n7159# a_n158_n7062# 0.133664f
C1885 w_n358_n183987# a_100_34582# 0.352467f
C1886 w_n358_n183987# a_n100_n143579# 0.269531f
C1887 a_n158_n149226# a_n158_n150662# 0.010536f
C1888 a_n158_116434# a_n158_114998# 0.010536f
C1889 w_n358_n183987# a_n100_122081# 0.269531f
C1890 a_100_n32910# a_100_n34346# 0.010536f
C1891 a_n100_n34443# a_n158_n34346# 0.133664f
C1892 a_n100_168033# a_n100_166597# 0.205388f
C1893 a_n158_168130# a_100_168130# 0.328443f
C1894 w_n358_n183987# a_n158_n54450# 0.352467f
C1895 w_n358_n183987# a_n100_67513# 0.269531f
C1896 a_n158_n176510# a_n158_n177946# 0.010536f
C1897 a_n158_89150# a_n158_87714# 0.010536f
C1898 a_100_n60194# a_100_n61630# 0.010536f
C1899 a_n100_n61727# a_n158_n61630# 0.133664f
C1900 w_n358_n183987# a_n158_2990# 0.352467f
C1901 a_n100_n17211# a_100_n17114# 0.133664f
C1902 w_n358_n183987# a_n158_n109018# 0.352467f
C1903 a_n158_61866# a_n158_60430# 0.010536f
C1904 w_n358_n183987# a_n100_12945# 0.269531f
C1905 a_n158_5862# a_n158_4426# 0.010536f
C1906 w_n358_n183987# a_100_n19986# 0.352467f
C1907 a_100_n87478# a_100_n88914# 0.010536f
C1908 a_n100_n89011# a_n158_n88914# 0.133664f
C1909 w_n358_n183987# a_n158_102074# 0.352467f
C1910 a_n100_n44495# a_100_n44398# 0.133664f
C1911 w_n358_n183987# a_n158_n163586# 0.352467f
C1912 a_n158_34582# a_n158_33146# 0.010536f
C1913 w_n358_n183987# a_100_n74554# 0.352467f
C1914 a_100_n114762# a_100_n116198# 0.010536f
C1915 a_n100_n116295# a_n158_n116198# 0.133664f
C1916 a_100_150898# a_100_149462# 0.010536f
C1917 a_n100_149365# a_n158_149462# 0.133664f
C1918 w_n358_n183987# a_n158_47506# 0.352467f
C1919 a_n100_n71779# a_100_n71682# 0.133664f
C1920 w_n358_n183987# a_100_136538# 0.352467f
C1921 w_n358_n183987# a_100_n129122# 0.352467f
C1922 a_100_n142046# a_100_n143482# 0.010536f
C1923 a_n100_n143579# a_n158_n143482# 0.133664f
C1924 a_100_123614# a_100_122178# 0.010536f
C1925 a_n100_122081# a_n158_122178# 0.133664f
C1926 a_n158_n27166# a_100_n27166# 0.328443f
C1927 a_n100_n27263# a_n100_n28699# 0.205388f
C1928 a_100_181054# a_100_179618# 0.010536f
C1929 a_n100_179521# a_n158_179618# 0.133664f
C1930 a_n100_n99063# a_100_n98966# 0.133664f
C1931 w_n358_n183987# a_n100_n41623# 0.269531f
C1932 a_100_96330# a_100_94894# 0.010536f
C1933 a_n100_94797# a_n158_94894# 0.133664f
C1934 w_n358_n183987# a_100_81970# 0.352467f
C1935 w_n358_n183987# a_100_n183690# 0.35701f
C1936 a_100_n169330# a_100_n170766# 0.010536f
C1937 a_n100_n170863# a_n158_n170766# 0.133664f
C1938 a_n158_n54450# a_100_n54450# 0.328443f
C1939 a_n100_n54547# a_n100_n55983# 0.205388f
C1940 a_n100_n126347# a_100_n126250# 0.133664f
C1941 a_n100_139313# a_100_139410# 0.133664f
C1942 w_n358_n183987# a_n100_n96191# 0.269531f
C1943 a_100_69046# a_100_67610# 0.010536f
C1944 a_n100_67513# a_n158_67610# 0.133664f
C1945 w_n358_n183987# a_100_27402# 0.352467f
C1946 w_n358_n183987# a_n158_n7062# 0.352467f
C1947 a_n158_n81734# a_100_n81734# 0.328443f
C1948 a_n100_n81831# a_n100_n83267# 0.205388f
C1949 a_n100_n153631# a_100_n153534# 0.133664f
C1950 a_n100_112029# a_100_112126# 0.133664f
C1951 w_n358_n183987# a_n100_114901# 0.269531f
C1952 w_n358_n183987# a_n100_n150759# 0.269531f
C1953 a_n158_2990# a_100_2990# 0.328443f
C1954 a_100_41762# a_100_40326# 0.010536f
C1955 a_n100_40229# a_n158_40326# 0.133664f
C1956 w_n358_n183987# a_n158_n61630# 0.352467f
C1957 a_n158_n109018# a_100_n109018# 0.328443f
C1958 a_n100_n109115# a_n100_n110551# 0.205388f
C1959 a_n100_n180915# a_100_n180818# 0.133664f
C1960 a_n100_84745# a_100_84842# 0.133664f
C1961 w_n358_n183987# a_n100_60333# 0.269531f
C1962 a_100_172438# a_100_171002# 0.010536f
C1963 a_100_14478# a_100_13042# 0.010536f
C1964 a_n100_12945# a_n158_13042# 0.133664f
C1965 a_n158_129358# a_100_129358# 0.328443f
C1966 a_n100_129261# a_n100_127825# 0.205388f
C1967 w_n358_n183987# a_n158_149462# 0.352467f
C1968 w_n358_n183987# a_n158_n116198# 0.352467f
C1969 a_n158_n136302# a_100_n136302# 0.328443f
C1970 a_n100_n136399# a_n100_n137835# 0.205388f
C1971 a_n158_n19986# a_n158_n21422# 0.010536f
C1972 a_n100_57461# a_100_57558# 0.133664f
C1973 a_n100_155109# a_100_155206# 0.133664f
C1974 w_n358_n183987# a_100_n27166# 0.352467f
C1975 w_n358_n183987# a_n158_179618# 0.352467f
C1976 a_n158_n163586# a_100_n163586# 0.328443f
C1977 a_n100_n163683# a_n100_n165119# 0.205388f
C1978 a_n158_102074# a_100_102074# 0.328443f
C1979 a_n100_101977# a_n100_100541# 0.205388f
C1980 w_n358_n183987# a_n158_94894# 0.352467f
C1981 w_n358_n183987# a_n158_n170766# 0.352467f
C1982 a_100_165258# a_100_163822# 0.010536f
C1983 a_n158_n47270# a_n158_n48706# 0.010536f
C1984 a_n100_163725# a_n158_163822# 0.133664f
C1985 a_n100_30177# a_100_30274# 0.133664f
C1986 w_n358_n183987# a_100_n81734# 0.352467f
C1987 a_n158_74790# a_100_74790# 0.328443f
C1988 a_n100_74693# a_n100_73257# 0.205388f
C1989 w_n358_n183987# a_n158_40326# 0.352467f
C1990 a_n158_n74554# a_n158_n75990# 0.010536f
C1991 w_n358_n183987# a_100_129358# 0.352467f
C1992 w_n358_n183987# a_100_n136302# 0.352467f
C1993 a_n158_47506# a_100_47506# 0.328443f
C1994 a_n100_47409# a_n100_45973# 0.205388f
C1995 a_n158_n101838# a_n158_n103274# 0.010536f
C1996 w_n358_n183987# a_n158_163822# 0.352467f
C1997 w_n358_n183987# a_n100_n48803# 0.269531f
C1998 w_n358_n183987# a_100_74790# 0.352467f
C1999 a_n158_20222# a_100_20222# 0.328443f
C2000 a_n100_20125# a_n100_18689# 0.205388f
C2001 a_n158_n129122# a_n158_n130558# 0.010536f
C2002 a_n158_136538# a_n158_135102# 0.010536f
C2003 a_100_156642# a_100_155206# 0.010536f
C2004 w_n358_n183987# a_n100_n103371# 0.269531f
C2005 a_100_n12806# a_100_n14242# 0.010536f
C2006 a_n100_n14339# a_n158_n14242# 0.133664f
C2007 w_n358_n183987# a_100_20222# 0.352467f
C2008 w_n358_n183987# a_n158_n14242# 0.352467f
C2009 w_n358_n183987# a_n100_n157939# 0.269531f
C2010 a_n158_n156406# a_n158_n157842# 0.010536f
C2011 a_n158_109254# a_n158_107818# 0.010536f
C2012 w_n358_n183987# a_n100_107721# 0.269531f
C2013 a_100_n40090# a_100_n41526# 0.010536f
C2014 a_n100_n41623# a_n158_n41526# 0.133664f
C2015 w_n358_n183987# a_100_7298# 0.352467f
C2016 w_n358_n183987# a_n158_n68810# 0.352467f
C2017 a_n158_81970# a_n158_80534# 0.010536f
C2018 w_n358_n183987# a_n100_53153# 0.269531f
C2019 a_100_n67374# a_100_n68810# 0.010536f
C2020 a_n100_n68907# a_n158_n68810# 0.133664f
C2021 w_n358_n183987# a_n100_173777# 0.269531f
C2022 a_n158_7298# a_100_7298# 0.328443f
C2023 w_n358_n183987# a_n158_n123378# 0.352467f
C2024 w_n358_n183987# a_n158_142282# 0.352467f
C2025 a_n100_n24391# a_100_n24294# 0.133664f
C2026 a_n158_54686# a_n158_53250# 0.010536f
C2027 a_100_n94658# a_100_n96094# 0.010536f
C2028 a_n100_n96191# a_n158_n96094# 0.133664f
C2029 w_n358_n183987# a_100_n34346# 0.352467f
C2030 w_n358_n183987# a_n100_166597# 0.269531f
C2031 a_n100_n51675# a_100_n51578# 0.133664f
C2032 w_n358_n183987# a_n158_n177946# 0.352467f
C2033 w_n358_n183987# a_n158_87714# 0.352467f
C2034 a_n158_27402# a_n158_25966# 0.010536f
C2035 w_n358_n183987# a_100_n88914# 0.352467f
C2036 a_100_n121942# a_100_n123378# 0.010536f
C2037 a_n100_n123475# a_n158_n123378# 0.133664f
C2038 a_100_143718# a_100_142282# 0.010536f
C2039 a_n100_142185# a_n158_142282# 0.133664f
C2040 a_n158_n7062# a_100_n7062# 0.328443f
C2041 a_n100_n7159# a_n100_n8595# 0.205388f
C2042 a_n100_n78959# a_100_n78862# 0.133664f
C2043 w_n358_n183987# a_n158_33146# 0.352467f
C2044 w_n358_n183987# a_n100_n1415# 0.269531f
C2045 w_n358_n183987# a_100_n143482# 0.352467f
C2046 a_100_n149226# a_100_n150662# 0.010536f
C2047 a_n100_n150759# a_n158_n150662# 0.133664f
C2048 a_100_116434# a_100_114998# 0.010536f
C2049 a_n100_114901# a_n158_114998# 0.133664f
C2050 w_n358_n183987# a_100_122178# 0.352467f
C2051 a_n158_n34346# a_100_n34346# 0.328443f
C2052 a_n100_n34443# a_n100_n35879# 0.205388f
C2053 a_n100_n106243# a_100_n106146# 0.133664f
C2054 a_n158_168130# a_n158_166694# 0.010536f
C2055 w_n358_n183987# a_n100_n55983# 0.269531f
C2056 a_100_n176510# a_100_n177946# 0.010536f
C2057 a_n100_n178043# a_n158_n177946# 0.133664f
C2058 a_100_89150# a_100_87714# 0.010536f
C2059 a_n100_87617# a_n158_87714# 0.133664f
C2060 w_n358_n183987# a_100_67610# 0.352467f
C2061 a_n158_n61630# a_100_n61630# 0.328443f
C2062 a_n100_n61727# a_n100_n63163# 0.205388f
C2063 a_n100_n133527# a_100_n133430# 0.133664f
C2064 a_n100_132133# a_100_132230# 0.133664f
C2065 w_n358_n183987# a_n100_n110551# 0.269531f
C2066 w_n358_n183987# a_100_13042# 0.352467f
C2067 a_100_5862# a_100_4426# 0.010536f
C2068 a_100_61866# a_100_60430# 0.010536f
C2069 a_n100_60333# a_n158_60430# 0.133664f
C2070 w_n358_n183987# a_n158_n21422# 0.352467f
C2071 a_n158_n88914# a_100_n88914# 0.328443f
C2072 a_n100_n89011# a_n100_n90447# 0.205388f
C2073 a_n100_n160811# a_100_n160714# 0.133664f
C2074 a_n100_104849# a_100_104946# 0.133664f
C2075 w_n358_n183987# a_n100_n165119# 0.269531f
C2076 w_n358_n183987# a_n100_100541# 0.269531f
C2077 a_100_34582# a_100_33146# 0.010536f
C2078 a_n100_33049# a_n158_33146# 0.133664f
C2079 w_n358_n183987# a_n158_n75990# 0.352467f
C2080 a_n158_n116198# a_100_n116198# 0.328443f
C2081 a_n100_n116295# a_n100_n117731# 0.205388f
C2082 a_n158_149462# a_100_149462# 0.328443f
C2083 a_n100_149365# a_n100_147929# 0.205388f
C2084 a_n100_77565# a_100_77662# 0.133664f
C2085 w_n358_n183987# a_n100_45973# 0.269531f
C2086 w_n358_n183987# a_n158_n130558# 0.352467f
C2087 a_n158_n143482# a_100_n143482# 0.328443f
C2088 a_n100_n143579# a_n100_n145015# 0.205388f
C2089 a_n158_122178# a_100_122178# 0.328443f
C2090 a_n100_122081# a_n100_120645# 0.205388f
C2091 w_n358_n183987# a_n158_135102# 0.352467f
C2092 a_n158_n27166# a_n158_n28602# 0.010536f
C2093 a_n100_50281# a_100_50378# 0.133664f
C2094 a_n158_179618# a_100_179618# 0.328443f
C2095 w_n358_n183987# a_100_n41526# 0.352467f
C2096 w_n358_n183987# a_n158_80534# 0.352467f
C2097 a_n158_n170766# a_100_n170766# 0.328443f
C2098 a_n100_n170863# a_n100_n172299# 0.205388f
C2099 a_n158_94894# a_100_94894# 0.328443f
C2100 a_n100_94797# a_n100_93361# 0.205388f
C2101 a_n158_n54450# a_n158_n55886# 0.010536f
C2102 a_n100_22997# a_100_23094# 0.133664f
C2103 w_n358_n183987# a_100_n96094# 0.352467f
C2104 w_n358_n183987# a_n158_173874# 0.352467f
C2105 a_n158_67610# a_100_67610# 0.328443f
C2106 a_n100_67513# a_n100_66077# 0.205388f
C2107 w_n358_n183987# a_n158_25966# 0.352467f
C2108 w_n358_n183987# a_n100_n8595# 0.269531f
C2109 a_n158_n81734# a_n158_n83170# 0.010536f
C2110 w_n358_n183987# a_100_114998# 0.352467f
C2111 w_n358_n183987# a_100_n150662# 0.352467f
C2112 a_n158_40326# a_100_40326# 0.328443f
C2113 a_n100_40229# a_n100_38793# 0.205388f
C2114 w_n358_n183987# a_n100_n63163# 0.269531f
C2115 a_n158_n109018# a_n158_n110454# 0.010536f
C2116 w_n358_n183987# a_100_60430# 0.352467f
C2117 a_n100_170905# a_n100_169469# 0.205388f
C2118 a_n158_13042# a_100_13042# 0.328443f
C2119 a_n100_12945# a_n100_11509# 0.205388f
C2120 w_n358_n183987# a_n100_147929# 0.269531f
C2121 w_n358_n183987# a_n100_n117731# 0.269531f
C2122 a_n158_n136302# a_n158_n137738# 0.010536f
C2123 a_n158_129358# a_n158_127922# 0.010536f
C2124 a_100_n19986# a_100_n21422# 0.010536f
C2125 a_n100_n21519# a_n158_n21422# 0.133664f
C2126 w_n358_n183987# a_n158_n28602# 0.352467f
C2127 a_n158_102074# a_n158_100638# 0.010536f
C2128 w_n358_n183987# a_n100_93361# 0.269531f
C2129 w_n358_n183987# a_n100_n172299# 0.269531f
C2130 a_n158_n163586# a_n158_n165022# 0.010536f
C2131 a_n158_163822# a_100_163822# 0.328443f
C2132 a_n100_163725# a_n100_162289# 0.205388f
C2133 a_100_n47270# a_100_n48706# 0.010536f
C2134 a_n100_n48803# a_n158_n48706# 0.133664f
C2135 a_n100_n4287# a_100_n4190# 0.133664f
C2136 w_n358_n183987# a_n158_n83170# 0.352467f
C2137 a_n158_74790# a_n158_73354# 0.010536f
C2138 w_n358_n183987# a_n100_38793# 0.269531f
C2139 a_100_n74554# a_100_n75990# 0.010536f
C2140 a_n100_n76087# a_n158_n75990# 0.133664f
C2141 w_n358_n183987# a_n158_171002# 0.352467f
C2142 w_n358_n183987# a_n158_127922# 0.352467f
C2143 a_n100_n31571# a_100_n31474# 0.133664f
C2144 w_n358_n183987# a_n158_n137738# 0.352467f
C2145 a_n158_47506# a_n158_46070# 0.010536f
C2146 w_n358_n183987# a_100_n48706# 0.352467f
C2147 w_n358_n183987# a_n100_162289# 0.269531f
C2148 a_100_n101838# a_100_n103274# 0.010536f
C2149 a_n100_n103371# a_n158_n103274# 0.133664f
C2150 w_n358_n183987# a_n158_73354# 0.352467f
C2151 a_n100_n58855# a_100_n58758# 0.133664f
C2152 a_n158_20222# a_n158_18786# 0.010536f
C2153 a_100_n129122# a_100_n130558# 0.010536f
C2154 a_n100_n130655# a_n158_n130558# 0.133664f
C2155 a_100_136538# a_100_135102# 0.010536f
C2156 a_n100_135005# a_n158_135102# 0.133664f
C2157 w_n358_n183987# a_100_n103274# 0.352467f
C2158 a_n158_n14242# a_100_n14242# 0.328443f
C2159 a_n100_n14339# a_n100_n15775# 0.205388f
C2160 w_n358_n183987# a_n100_n15775# 0.269531f
C2161 w_n358_n183987# a_n158_18786# 0.352467f
C2162 a_n100_n86139# a_100_n86042# 0.133664f
C2163 a_100_n156406# a_100_n157842# 0.010536f
C2164 a_n100_n157939# a_n158_n157842# 0.133664f
C2165 a_100_109254# a_100_107818# 0.010536f
C2166 a_n100_107721# a_n158_107818# 0.133664f
C2167 w_n358_n183987# a_100_107818# 0.352467f
C2168 w_n358_n183987# a_100_n157842# 0.352467f
C2169 a_n158_n41526# a_100_n41526# 0.328443f
C2170 a_n100_n41623# a_n100_n43059# 0.205388f
C2171 a_n100_n113423# a_100_n113326# 0.133664f
C2172 a_n100_152237# a_100_152334# 0.133664f
C2173 w_n358_n183987# a_n100_n70343# 0.269531f
C2174 a_100_81970# a_100_80534# 0.010536f
C2175 a_n100_80437# a_n158_80534# 0.133664f
C2176 w_n358_n183987# a_100_53250# 0.352467f
C2177 a_n158_n68810# a_100_n68810# 0.328443f
C2178 a_n100_n68907# a_n100_n70343# 0.205388f
C2179 a_n100_n140707# a_100_n140610# 0.133664f
C2180 a_n100_124953# a_100_125050# 0.133664f
C2181 w_n358_n183987# a_n100_140749# 0.269531f
C2182 w_n358_n183987# a_n100_n124911# 0.269531f
C2183 a_100_54686# a_100_53250# 0.010536f
C2184 a_n100_53153# a_n158_53250# 0.133664f
C2185 a_n158_n96094# a_100_n96094# 0.328443f
C2186 a_n100_n96191# a_n100_n97627# 0.205388f
C2187 w_n358_n183987# a_n158_n35782# 0.352467f
C2188 w_n358_n183987# a_100_166694# 0.352467f
C2189 a_n100_n167991# a_100_n167894# 0.133664f
C2190 a_n100_97669# a_100_97766# 0.133664f
C2191 w_n358_n183987# a_n100_n179479# 0.269531f
C2192 w_n358_n183987# a_n100_86181# 0.269531f
C2193 a_100_27402# a_100_25966# 0.010536f
C2194 a_n100_25869# a_n158_25966# 0.133664f
C2195 a_n158_n123378# a_100_n123378# 0.328443f
C2196 a_n100_n123475# a_n100_n124911# 0.205388f
C2197 a_n158_142282# a_100_142282# 0.328443f
C2198 a_n100_142185# a_n100_140749# 0.205388f
C2199 w_n358_n183987# a_n158_n90350# 0.352467f
C2200 a_n100_70385# a_100_70482# 0.133664f
C2201 a_n158_n7062# a_n158_n8498# 0.010536f
C2202 w_n358_n183987# a_100_n1318# 0.352467f
C2203 w_n358_n183987# a_n100_31613# 0.269531f
C2204 w_n358_n183987# a_n158_n144918# 0.352467f
C2205 a_n158_n150662# a_100_n150662# 0.328443f
C2206 a_n100_n150759# a_n100_n152195# 0.205388f
C2207 a_n158_114998# a_100_114998# 0.328443f
C2208 a_n100_114901# a_n100_113465# 0.205388f
C2209 w_n358_n183987# a_n158_120742# 0.352467f
C2210 a_n100_43101# a_100_43198# 0.133664f
C2211 a_n158_n34346# a_n158_n35782# 0.010536f
C2212 a_n100_166597# a_n158_166694# 0.133664f
C2213 a_100_168130# a_100_166694# 0.010536f
C2214 w_n358_n183987# a_100_n55886# 0.352467f
C2215 a_n158_n177946# a_100_n177946# 0.328443f
C2216 a_n100_n178043# a_n100_n179479# 0.205388f
C2217 a_n158_87714# a_100_87714# 0.328443f
C2218 a_n100_87617# a_n100_86181# 0.205388f
C2219 w_n358_n183987# a_n158_66174# 0.352467f
C2220 a_n158_n61630# a_n158_n63066# 0.010536f
C2221 a_n100_15817# a_100_15914# 0.133664f
C2222 w_n358_n183987# a_100_n110454# 0.352467f
C2223 w_n358_n183987# a_n100_5765# 0.269531f
C2224 w_n358_n183987# a_100_155206# 0.352467f
C2225 a_n158_60430# a_100_60430# 0.328443f
C2226 a_n100_60333# a_n100_58897# 0.205388f
C2227 w_n358_n183987# a_n158_11606# 0.352467f
C2228 a_n158_n88914# a_n158_n90350# 0.010536f
C2229 w_n358_n183987# a_n100_n22955# 0.269531f
C2230 w_n358_n183987# a_100_n165022# 0.352467f
C2231 w_n358_n183987# a_100_100638# 0.352467f
C2232 a_n158_33146# a_100_33146# 0.328443f
C2233 a_n100_33049# a_n100_31613# 0.205388f
C2234 w_n358_n183987# a_n100_n77523# 0.269531f
C2235 a_n158_n116198# a_n158_n117634# 0.010536f
C2236 a_n158_149462# a_n158_148026# 0.010536f
C2237 a_n100_n1415# a_n158_n1318# 0.133664f
C2238 w_n358_n183987# a_100_46070# 0.352467f
C2239 w_n358_n183987# a_n100_n132091# 0.269531f
C2240 a_n158_n143482# a_n158_n144918# 0.010536f
C2241 a_n158_122178# a_n158_120742# 0.010536f
C2242 w_n358_n183987# a_n100_133569# 0.269531f
C2243 a_100_n27166# a_100_n28602# 0.010536f
C2244 a_n100_n28699# a_n158_n28602# 0.133664f
C2245 w_n358_n183987# a_n158_n42962# 0.352467f
C2246 a_100_1554# a_100_118# 0.010536f
C2247 a_n100_21# a_n158_118# 0.133664f
C2248 a_n158_n170766# a_n158_n172202# 0.010536f
C2249 a_n158_94894# a_n158_93458# 0.010536f
C2250 w_n358_n183987# a_n100_79001# 0.269531f
C2251 a_100_n54450# a_100_n55886# 0.010536f
C2252 a_n100_n55983# a_n158_n55886# 0.133664f
C2253 w_n358_n183987# a_n158_n97530# 0.352467f
C2254 a_n100_n11467# a_100_n11370# 0.133664f
C2255 w_n358_n183987# a_n100_172341# 0.269531f
C2256 w_n358_n183987# a_n100_24433# 0.269531f
C2257 a_n158_67610# a_n158_66174# 0.010536f
C2258 w_n358_n183987# a_100_n8498# 0.352467f
C2259 a_100_n81734# a_100_n83170# 0.010536f
C2260 a_n100_n83267# a_n158_n83170# 0.133664f
C2261 a_n100_n38751# a_100_n38654# 0.133664f
C2262 w_n358_n183987# a_n158_n152098# 0.352467f
C2263 w_n358_n183987# a_n158_1554# 0.352467f
C2264 w_n358_n183987# a_n158_113562# 0.352467f
C2265 a_n158_40326# a_n158_38890# 0.010536f
C2266 a_n100_173777# a_100_173874# 0.133664f
C2267 a_n100_4329# a_100_4426# 0.133664f
C2268 w_n358_n183987# a_100_n63066# 0.352467f
C2269 a_100_n109018# a_100_n110454# 0.010536f
C2270 a_n100_n110551# a_n158_n110454# 0.133664f
C2271 w_n358_n183987# a_n158_58994# 0.352467f
C2272 a_n100_n66035# a_100_n65938# 0.133664f
C2273 a_n158_13042# a_n158_11606# 0.010536f
C2274 a_n158_n21422# a_100_n21422# 0.328443f
C2275 a_n100_n21519# a_n100_n22955# 0.205388f
C2276 w_n358_n183987# a_100_n117634# 0.352467f
C2277 a_100_n136302# a_100_n137738# 0.010536f
C2278 a_n100_n137835# a_n158_n137738# 0.133664f
C2279 a_100_129358# a_100_127922# 0.010536f
C2280 a_n100_127825# a_n158_127922# 0.133664f
C2281 w_n358_n183987# a_100_148026# 0.352467f
C2282 w_n358_n183987# a_n100_n30135# 0.269531f
C2283 a_n100_n93319# a_100_n93222# 0.133664f
C2284 w_n358_n183987# a_100_93458# 0.352467f
C2285 w_n358_n183987# a_100_n172202# 0.352467f
C2286 a_100_n163586# a_100_n165022# 0.010536f
C2287 a_n100_n165119# a_n158_n165022# 0.133664f
C2288 a_100_102074# a_100_100638# 0.010536f
C2289 a_n100_100541# a_n158_100638# 0.133664f
C2290 a_n158_163822# a_n158_162386# 0.010536f
C2291 a_n158_n48706# a_100_n48706# 0.328443f
C2292 a_n100_n48803# a_n100_n50239# 0.205388f
C2293 w_n358_n183987# a_n100_n84703# 0.269531f
C2294 a_n100_n120603# a_100_n120506# 0.133664f
C2295 a_n100_145057# a_100_145154# 0.133664f
C2296 a_100_74790# a_100_73354# 0.010536f
C2297 a_n100_73257# a_n158_73354# 0.133664f
C2298 w_n358_n183987# a_100_38890# 0.352467f
C2299 a_n158_n75990# a_100_n75990# 0.328443f
C2300 a_n100_n76087# a_n100_n77523# 0.205388f
C2301 a_100_n183690# VSUBS 0.292592f
C2302 a_n158_n183690# VSUBS 0.292592f
C2303 a_n100_n183787# VSUBS 0.265338f
C2304 a_100_n182254# VSUBS 0.287142f
C2305 a_n158_n182254# VSUBS 0.287142f
C2306 a_n100_n182351# VSUBS 0.221608f
C2307 a_100_n180818# VSUBS 0.287142f
C2308 a_n158_n180818# VSUBS 0.287142f
C2309 a_n100_n180915# VSUBS 0.221608f
C2310 a_100_n179382# VSUBS 0.287142f
C2311 a_n158_n179382# VSUBS 0.287142f
C2312 a_n100_n179479# VSUBS 0.221608f
C2313 a_100_n177946# VSUBS 0.287142f
C2314 a_n158_n177946# VSUBS 0.287142f
C2315 a_n100_n178043# VSUBS 0.221608f
C2316 a_100_n176510# VSUBS 0.287142f
C2317 a_n158_n176510# VSUBS 0.287142f
C2318 a_n100_n176607# VSUBS 0.221608f
C2319 a_100_n175074# VSUBS 0.287142f
C2320 a_n158_n175074# VSUBS 0.287142f
C2321 a_n100_n175171# VSUBS 0.221608f
C2322 a_100_n173638# VSUBS 0.287142f
C2323 a_n158_n173638# VSUBS 0.287142f
C2324 a_n100_n173735# VSUBS 0.221608f
C2325 a_100_n172202# VSUBS 0.287142f
C2326 a_n158_n172202# VSUBS 0.287142f
C2327 a_n100_n172299# VSUBS 0.221608f
C2328 a_100_n170766# VSUBS 0.287142f
C2329 a_n158_n170766# VSUBS 0.287142f
C2330 a_n100_n170863# VSUBS 0.221608f
C2331 a_100_n169330# VSUBS 0.287142f
C2332 a_n158_n169330# VSUBS 0.287142f
C2333 a_n100_n169427# VSUBS 0.221608f
C2334 a_100_n167894# VSUBS 0.287142f
C2335 a_n158_n167894# VSUBS 0.287142f
C2336 a_n100_n167991# VSUBS 0.221608f
C2337 a_100_n166458# VSUBS 0.287142f
C2338 a_n158_n166458# VSUBS 0.287142f
C2339 a_n100_n166555# VSUBS 0.221608f
C2340 a_100_n165022# VSUBS 0.287142f
C2341 a_n158_n165022# VSUBS 0.287142f
C2342 a_n100_n165119# VSUBS 0.221608f
C2343 a_100_n163586# VSUBS 0.287142f
C2344 a_n158_n163586# VSUBS 0.287142f
C2345 a_n100_n163683# VSUBS 0.221608f
C2346 a_100_n162150# VSUBS 0.287142f
C2347 a_n158_n162150# VSUBS 0.287142f
C2348 a_n100_n162247# VSUBS 0.221608f
C2349 a_100_n160714# VSUBS 0.287142f
C2350 a_n158_n160714# VSUBS 0.287142f
C2351 a_n100_n160811# VSUBS 0.221608f
C2352 a_100_n159278# VSUBS 0.287142f
C2353 a_n158_n159278# VSUBS 0.287142f
C2354 a_n100_n159375# VSUBS 0.221608f
C2355 a_100_n157842# VSUBS 0.287142f
C2356 a_n158_n157842# VSUBS 0.287142f
C2357 a_n100_n157939# VSUBS 0.221608f
C2358 a_100_n156406# VSUBS 0.287142f
C2359 a_n158_n156406# VSUBS 0.287142f
C2360 a_n100_n156503# VSUBS 0.221608f
C2361 a_100_n154970# VSUBS 0.287142f
C2362 a_n158_n154970# VSUBS 0.287142f
C2363 a_n100_n155067# VSUBS 0.221608f
C2364 a_100_n153534# VSUBS 0.287142f
C2365 a_n158_n153534# VSUBS 0.287142f
C2366 a_n100_n153631# VSUBS 0.221608f
C2367 a_100_n152098# VSUBS 0.287142f
C2368 a_n158_n152098# VSUBS 0.287142f
C2369 a_n100_n152195# VSUBS 0.221608f
C2370 a_100_n150662# VSUBS 0.287142f
C2371 a_n158_n150662# VSUBS 0.287142f
C2372 a_n100_n150759# VSUBS 0.221608f
C2373 a_100_n149226# VSUBS 0.287142f
C2374 a_n158_n149226# VSUBS 0.287142f
C2375 a_n100_n149323# VSUBS 0.221608f
C2376 a_100_n147790# VSUBS 0.287142f
C2377 a_n158_n147790# VSUBS 0.287142f
C2378 a_n100_n147887# VSUBS 0.221608f
C2379 a_100_n146354# VSUBS 0.287142f
C2380 a_n158_n146354# VSUBS 0.287142f
C2381 a_n100_n146451# VSUBS 0.221608f
C2382 a_100_n144918# VSUBS 0.287142f
C2383 a_n158_n144918# VSUBS 0.287142f
C2384 a_n100_n145015# VSUBS 0.221608f
C2385 a_100_n143482# VSUBS 0.287142f
C2386 a_n158_n143482# VSUBS 0.287142f
C2387 a_n100_n143579# VSUBS 0.221608f
C2388 a_100_n142046# VSUBS 0.287142f
C2389 a_n158_n142046# VSUBS 0.287142f
C2390 a_n100_n142143# VSUBS 0.221608f
C2391 a_100_n140610# VSUBS 0.287142f
C2392 a_n158_n140610# VSUBS 0.287142f
C2393 a_n100_n140707# VSUBS 0.221608f
C2394 a_100_n139174# VSUBS 0.287142f
C2395 a_n158_n139174# VSUBS 0.287142f
C2396 a_n100_n139271# VSUBS 0.221608f
C2397 a_100_n137738# VSUBS 0.287142f
C2398 a_n158_n137738# VSUBS 0.287142f
C2399 a_n100_n137835# VSUBS 0.221608f
C2400 a_100_n136302# VSUBS 0.287142f
C2401 a_n158_n136302# VSUBS 0.287142f
C2402 a_n100_n136399# VSUBS 0.221608f
C2403 a_100_n134866# VSUBS 0.287142f
C2404 a_n158_n134866# VSUBS 0.287142f
C2405 a_n100_n134963# VSUBS 0.221608f
C2406 a_100_n133430# VSUBS 0.287142f
C2407 a_n158_n133430# VSUBS 0.287142f
C2408 a_n100_n133527# VSUBS 0.221608f
C2409 a_100_n131994# VSUBS 0.287142f
C2410 a_n158_n131994# VSUBS 0.287142f
C2411 a_n100_n132091# VSUBS 0.221608f
C2412 a_100_n130558# VSUBS 0.287142f
C2413 a_n158_n130558# VSUBS 0.287142f
C2414 a_n100_n130655# VSUBS 0.221608f
C2415 a_100_n129122# VSUBS 0.287142f
C2416 a_n158_n129122# VSUBS 0.287142f
C2417 a_n100_n129219# VSUBS 0.221608f
C2418 a_100_n127686# VSUBS 0.287142f
C2419 a_n158_n127686# VSUBS 0.287142f
C2420 a_n100_n127783# VSUBS 0.221608f
C2421 a_100_n126250# VSUBS 0.287142f
C2422 a_n158_n126250# VSUBS 0.287142f
C2423 a_n100_n126347# VSUBS 0.221608f
C2424 a_100_n124814# VSUBS 0.287142f
C2425 a_n158_n124814# VSUBS 0.287142f
C2426 a_n100_n124911# VSUBS 0.221608f
C2427 a_100_n123378# VSUBS 0.287142f
C2428 a_n158_n123378# VSUBS 0.287142f
C2429 a_n100_n123475# VSUBS 0.221608f
C2430 a_100_n121942# VSUBS 0.287142f
C2431 a_n158_n121942# VSUBS 0.287142f
C2432 a_n100_n122039# VSUBS 0.221608f
C2433 a_100_n120506# VSUBS 0.287142f
C2434 a_n158_n120506# VSUBS 0.287142f
C2435 a_n100_n120603# VSUBS 0.221608f
C2436 a_100_n119070# VSUBS 0.287142f
C2437 a_n158_n119070# VSUBS 0.287142f
C2438 a_n100_n119167# VSUBS 0.221608f
C2439 a_100_n117634# VSUBS 0.287142f
C2440 a_n158_n117634# VSUBS 0.287142f
C2441 a_n100_n117731# VSUBS 0.221608f
C2442 a_100_n116198# VSUBS 0.287142f
C2443 a_n158_n116198# VSUBS 0.287142f
C2444 a_n100_n116295# VSUBS 0.221608f
C2445 a_100_n114762# VSUBS 0.287142f
C2446 a_n158_n114762# VSUBS 0.287142f
C2447 a_n100_n114859# VSUBS 0.221608f
C2448 a_100_n113326# VSUBS 0.287142f
C2449 a_n158_n113326# VSUBS 0.287142f
C2450 a_n100_n113423# VSUBS 0.221608f
C2451 a_100_n111890# VSUBS 0.287142f
C2452 a_n158_n111890# VSUBS 0.287142f
C2453 a_n100_n111987# VSUBS 0.221608f
C2454 a_100_n110454# VSUBS 0.287142f
C2455 a_n158_n110454# VSUBS 0.287142f
C2456 a_n100_n110551# VSUBS 0.221608f
C2457 a_100_n109018# VSUBS 0.287142f
C2458 a_n158_n109018# VSUBS 0.287142f
C2459 a_n100_n109115# VSUBS 0.221608f
C2460 a_100_n107582# VSUBS 0.287142f
C2461 a_n158_n107582# VSUBS 0.287142f
C2462 a_n100_n107679# VSUBS 0.221608f
C2463 a_100_n106146# VSUBS 0.287142f
C2464 a_n158_n106146# VSUBS 0.287142f
C2465 a_n100_n106243# VSUBS 0.221608f
C2466 a_100_n104710# VSUBS 0.287142f
C2467 a_n158_n104710# VSUBS 0.287142f
C2468 a_n100_n104807# VSUBS 0.221608f
C2469 a_100_n103274# VSUBS 0.287142f
C2470 a_n158_n103274# VSUBS 0.287142f
C2471 a_n100_n103371# VSUBS 0.221608f
C2472 a_100_n101838# VSUBS 0.287142f
C2473 a_n158_n101838# VSUBS 0.287142f
C2474 a_n100_n101935# VSUBS 0.221608f
C2475 a_100_n100402# VSUBS 0.287142f
C2476 a_n158_n100402# VSUBS 0.287142f
C2477 a_n100_n100499# VSUBS 0.221608f
C2478 a_100_n98966# VSUBS 0.287142f
C2479 a_n158_n98966# VSUBS 0.287142f
C2480 a_n100_n99063# VSUBS 0.221608f
C2481 a_100_n97530# VSUBS 0.287142f
C2482 a_n158_n97530# VSUBS 0.287142f
C2483 a_n100_n97627# VSUBS 0.221608f
C2484 a_100_n96094# VSUBS 0.287142f
C2485 a_n158_n96094# VSUBS 0.287142f
C2486 a_n100_n96191# VSUBS 0.221608f
C2487 a_100_n94658# VSUBS 0.287142f
C2488 a_n158_n94658# VSUBS 0.287142f
C2489 a_n100_n94755# VSUBS 0.221608f
C2490 a_100_n93222# VSUBS 0.287142f
C2491 a_n158_n93222# VSUBS 0.287142f
C2492 a_n100_n93319# VSUBS 0.221608f
C2493 a_100_n91786# VSUBS 0.287142f
C2494 a_n158_n91786# VSUBS 0.287142f
C2495 a_n100_n91883# VSUBS 0.221608f
C2496 a_100_n90350# VSUBS 0.287142f
C2497 a_n158_n90350# VSUBS 0.287142f
C2498 a_n100_n90447# VSUBS 0.221608f
C2499 a_100_n88914# VSUBS 0.287142f
C2500 a_n158_n88914# VSUBS 0.287142f
C2501 a_n100_n89011# VSUBS 0.221608f
C2502 a_100_n87478# VSUBS 0.287142f
C2503 a_n158_n87478# VSUBS 0.287142f
C2504 a_n100_n87575# VSUBS 0.221608f
C2505 a_100_n86042# VSUBS 0.287142f
C2506 a_n158_n86042# VSUBS 0.287142f
C2507 a_n100_n86139# VSUBS 0.221608f
C2508 a_100_n84606# VSUBS 0.287142f
C2509 a_n158_n84606# VSUBS 0.287142f
C2510 a_n100_n84703# VSUBS 0.221608f
C2511 a_100_n83170# VSUBS 0.287142f
C2512 a_n158_n83170# VSUBS 0.287142f
C2513 a_n100_n83267# VSUBS 0.221608f
C2514 a_100_n81734# VSUBS 0.287142f
C2515 a_n158_n81734# VSUBS 0.287142f
C2516 a_n100_n81831# VSUBS 0.221608f
C2517 a_100_n80298# VSUBS 0.287142f
C2518 a_n158_n80298# VSUBS 0.287142f
C2519 a_n100_n80395# VSUBS 0.221608f
C2520 a_100_n78862# VSUBS 0.287142f
C2521 a_n158_n78862# VSUBS 0.287142f
C2522 a_n100_n78959# VSUBS 0.221608f
C2523 a_100_n77426# VSUBS 0.287142f
C2524 a_n158_n77426# VSUBS 0.287142f
C2525 a_n100_n77523# VSUBS 0.221608f
C2526 a_100_n75990# VSUBS 0.287142f
C2527 a_n158_n75990# VSUBS 0.287142f
C2528 a_n100_n76087# VSUBS 0.221608f
C2529 a_100_n74554# VSUBS 0.287142f
C2530 a_n158_n74554# VSUBS 0.287142f
C2531 a_n100_n74651# VSUBS 0.221608f
C2532 a_100_n73118# VSUBS 0.287142f
C2533 a_n158_n73118# VSUBS 0.287142f
C2534 a_n100_n73215# VSUBS 0.221608f
C2535 a_100_n71682# VSUBS 0.287142f
C2536 a_n158_n71682# VSUBS 0.287142f
C2537 a_n100_n71779# VSUBS 0.221608f
C2538 a_100_n70246# VSUBS 0.287142f
C2539 a_n158_n70246# VSUBS 0.287142f
C2540 a_n100_n70343# VSUBS 0.221608f
C2541 a_100_n68810# VSUBS 0.287142f
C2542 a_n158_n68810# VSUBS 0.287142f
C2543 a_n100_n68907# VSUBS 0.221608f
C2544 a_100_n67374# VSUBS 0.287142f
C2545 a_n158_n67374# VSUBS 0.287142f
C2546 a_n100_n67471# VSUBS 0.221608f
C2547 a_100_n65938# VSUBS 0.287142f
C2548 a_n158_n65938# VSUBS 0.287142f
C2549 a_n100_n66035# VSUBS 0.221608f
C2550 a_100_n64502# VSUBS 0.287142f
C2551 a_n158_n64502# VSUBS 0.287142f
C2552 a_n100_n64599# VSUBS 0.221608f
C2553 a_100_n63066# VSUBS 0.287142f
C2554 a_n158_n63066# VSUBS 0.287142f
C2555 a_n100_n63163# VSUBS 0.221608f
C2556 a_100_n61630# VSUBS 0.287142f
C2557 a_n158_n61630# VSUBS 0.287142f
C2558 a_n100_n61727# VSUBS 0.221608f
C2559 a_100_n60194# VSUBS 0.287142f
C2560 a_n158_n60194# VSUBS 0.287142f
C2561 a_n100_n60291# VSUBS 0.221608f
C2562 a_100_n58758# VSUBS 0.287142f
C2563 a_n158_n58758# VSUBS 0.287142f
C2564 a_n100_n58855# VSUBS 0.221608f
C2565 a_100_n57322# VSUBS 0.287142f
C2566 a_n158_n57322# VSUBS 0.287142f
C2567 a_n100_n57419# VSUBS 0.221608f
C2568 a_100_n55886# VSUBS 0.287142f
C2569 a_n158_n55886# VSUBS 0.287142f
C2570 a_n100_n55983# VSUBS 0.221608f
C2571 a_100_n54450# VSUBS 0.287142f
C2572 a_n158_n54450# VSUBS 0.287142f
C2573 a_n100_n54547# VSUBS 0.221608f
C2574 a_100_n53014# VSUBS 0.287142f
C2575 a_n158_n53014# VSUBS 0.287142f
C2576 a_n100_n53111# VSUBS 0.221608f
C2577 a_100_n51578# VSUBS 0.287142f
C2578 a_n158_n51578# VSUBS 0.287142f
C2579 a_n100_n51675# VSUBS 0.221608f
C2580 a_100_n50142# VSUBS 0.287142f
C2581 a_n158_n50142# VSUBS 0.287142f
C2582 a_n100_n50239# VSUBS 0.221608f
C2583 a_100_n48706# VSUBS 0.287142f
C2584 a_n158_n48706# VSUBS 0.287142f
C2585 a_n100_n48803# VSUBS 0.221608f
C2586 a_100_n47270# VSUBS 0.287142f
C2587 a_n158_n47270# VSUBS 0.287142f
C2588 a_n100_n47367# VSUBS 0.221608f
C2589 a_100_n45834# VSUBS 0.287142f
C2590 a_n158_n45834# VSUBS 0.287142f
C2591 a_n100_n45931# VSUBS 0.221608f
C2592 a_100_n44398# VSUBS 0.287142f
C2593 a_n158_n44398# VSUBS 0.287142f
C2594 a_n100_n44495# VSUBS 0.221608f
C2595 a_100_n42962# VSUBS 0.287142f
C2596 a_n158_n42962# VSUBS 0.287142f
C2597 a_n100_n43059# VSUBS 0.221608f
C2598 a_100_n41526# VSUBS 0.287142f
C2599 a_n158_n41526# VSUBS 0.287142f
C2600 a_n100_n41623# VSUBS 0.221608f
C2601 a_100_n40090# VSUBS 0.287142f
C2602 a_n158_n40090# VSUBS 0.287142f
C2603 a_n100_n40187# VSUBS 0.221608f
C2604 a_100_n38654# VSUBS 0.287142f
C2605 a_n158_n38654# VSUBS 0.287142f
C2606 a_n100_n38751# VSUBS 0.221608f
C2607 a_100_n37218# VSUBS 0.287142f
C2608 a_n158_n37218# VSUBS 0.287142f
C2609 a_n100_n37315# VSUBS 0.221608f
C2610 a_100_n35782# VSUBS 0.287142f
C2611 a_n158_n35782# VSUBS 0.287142f
C2612 a_n100_n35879# VSUBS 0.221608f
C2613 a_100_n34346# VSUBS 0.287142f
C2614 a_n158_n34346# VSUBS 0.287142f
C2615 a_n100_n34443# VSUBS 0.221608f
C2616 a_100_n32910# VSUBS 0.287142f
C2617 a_n158_n32910# VSUBS 0.287142f
C2618 a_n100_n33007# VSUBS 0.221608f
C2619 a_100_n31474# VSUBS 0.287142f
C2620 a_n158_n31474# VSUBS 0.287142f
C2621 a_n100_n31571# VSUBS 0.221608f
C2622 a_100_n30038# VSUBS 0.287142f
C2623 a_n158_n30038# VSUBS 0.287142f
C2624 a_n100_n30135# VSUBS 0.221608f
C2625 a_100_n28602# VSUBS 0.287142f
C2626 a_n158_n28602# VSUBS 0.287142f
C2627 a_n100_n28699# VSUBS 0.221608f
C2628 a_100_n27166# VSUBS 0.287142f
C2629 a_n158_n27166# VSUBS 0.287142f
C2630 a_n100_n27263# VSUBS 0.221608f
C2631 a_100_n25730# VSUBS 0.287142f
C2632 a_n158_n25730# VSUBS 0.287142f
C2633 a_n100_n25827# VSUBS 0.221608f
C2634 a_100_n24294# VSUBS 0.287142f
C2635 a_n158_n24294# VSUBS 0.287142f
C2636 a_n100_n24391# VSUBS 0.221608f
C2637 a_100_n22858# VSUBS 0.287142f
C2638 a_n158_n22858# VSUBS 0.287142f
C2639 a_n100_n22955# VSUBS 0.221608f
C2640 a_100_n21422# VSUBS 0.287142f
C2641 a_n158_n21422# VSUBS 0.287142f
C2642 a_n100_n21519# VSUBS 0.221608f
C2643 a_100_n19986# VSUBS 0.287142f
C2644 a_n158_n19986# VSUBS 0.287142f
C2645 a_n100_n20083# VSUBS 0.221608f
C2646 a_100_n18550# VSUBS 0.287142f
C2647 a_n158_n18550# VSUBS 0.287142f
C2648 a_n100_n18647# VSUBS 0.221608f
C2649 a_100_n17114# VSUBS 0.287142f
C2650 a_n158_n17114# VSUBS 0.287142f
C2651 a_n100_n17211# VSUBS 0.221608f
C2652 a_100_n15678# VSUBS 0.287142f
C2653 a_n158_n15678# VSUBS 0.287142f
C2654 a_n100_n15775# VSUBS 0.221608f
C2655 a_100_n14242# VSUBS 0.287142f
C2656 a_n158_n14242# VSUBS 0.287142f
C2657 a_n100_n14339# VSUBS 0.221608f
C2658 a_100_n12806# VSUBS 0.287142f
C2659 a_n158_n12806# VSUBS 0.287142f
C2660 a_n100_n12903# VSUBS 0.221608f
C2661 a_100_n11370# VSUBS 0.287142f
C2662 a_n158_n11370# VSUBS 0.287142f
C2663 a_n100_n11467# VSUBS 0.221608f
C2664 a_100_n9934# VSUBS 0.287142f
C2665 a_n158_n9934# VSUBS 0.287142f
C2666 a_n100_n10031# VSUBS 0.221608f
C2667 a_100_n8498# VSUBS 0.287142f
C2668 a_n158_n8498# VSUBS 0.287142f
C2669 a_n100_n8595# VSUBS 0.221608f
C2670 a_100_n7062# VSUBS 0.287142f
C2671 a_n158_n7062# VSUBS 0.287142f
C2672 a_n100_n7159# VSUBS 0.221608f
C2673 a_100_n5626# VSUBS 0.287142f
C2674 a_n158_n5626# VSUBS 0.287142f
C2675 a_n100_n5723# VSUBS 0.221608f
C2676 a_100_n4190# VSUBS 0.287142f
C2677 a_n158_n4190# VSUBS 0.287142f
C2678 a_n100_n4287# VSUBS 0.221608f
C2679 a_100_n2754# VSUBS 0.287142f
C2680 a_n158_n2754# VSUBS 0.287142f
C2681 a_n100_n2851# VSUBS 0.221608f
C2682 a_100_n1318# VSUBS 0.287142f
C2683 a_n158_n1318# VSUBS 0.287142f
C2684 a_n100_n1415# VSUBS 0.221608f
C2685 a_100_118# VSUBS 0.287142f
C2686 a_n158_118# VSUBS 0.287142f
C2687 a_n100_21# VSUBS 0.221608f
C2688 a_100_1554# VSUBS 0.287142f
C2689 a_n158_1554# VSUBS 0.287142f
C2690 a_n100_1457# VSUBS 0.221608f
C2691 a_100_2990# VSUBS 0.287142f
C2692 a_n158_2990# VSUBS 0.287142f
C2693 a_n100_2893# VSUBS 0.221608f
C2694 a_100_4426# VSUBS 0.287142f
C2695 a_n158_4426# VSUBS 0.287142f
C2696 a_n100_4329# VSUBS 0.221608f
C2697 a_100_5862# VSUBS 0.287142f
C2698 a_n158_5862# VSUBS 0.287142f
C2699 a_n100_5765# VSUBS 0.221608f
C2700 a_100_7298# VSUBS 0.287142f
C2701 a_n158_7298# VSUBS 0.287142f
C2702 a_n100_7201# VSUBS 0.221608f
C2703 a_100_8734# VSUBS 0.287142f
C2704 a_n158_8734# VSUBS 0.287142f
C2705 a_n100_8637# VSUBS 0.221608f
C2706 a_100_10170# VSUBS 0.287142f
C2707 a_n158_10170# VSUBS 0.287142f
C2708 a_n100_10073# VSUBS 0.221608f
C2709 a_100_11606# VSUBS 0.287142f
C2710 a_n158_11606# VSUBS 0.287142f
C2711 a_n100_11509# VSUBS 0.221608f
C2712 a_100_13042# VSUBS 0.287142f
C2713 a_n158_13042# VSUBS 0.287142f
C2714 a_n100_12945# VSUBS 0.221608f
C2715 a_100_14478# VSUBS 0.287142f
C2716 a_n158_14478# VSUBS 0.287142f
C2717 a_n100_14381# VSUBS 0.221608f
C2718 a_100_15914# VSUBS 0.287142f
C2719 a_n158_15914# VSUBS 0.287142f
C2720 a_n100_15817# VSUBS 0.221608f
C2721 a_100_17350# VSUBS 0.287142f
C2722 a_n158_17350# VSUBS 0.287142f
C2723 a_n100_17253# VSUBS 0.221608f
C2724 a_100_18786# VSUBS 0.287142f
C2725 a_n158_18786# VSUBS 0.287142f
C2726 a_n100_18689# VSUBS 0.221608f
C2727 a_100_20222# VSUBS 0.287142f
C2728 a_n158_20222# VSUBS 0.287142f
C2729 a_n100_20125# VSUBS 0.221608f
C2730 a_100_21658# VSUBS 0.287142f
C2731 a_n158_21658# VSUBS 0.287142f
C2732 a_n100_21561# VSUBS 0.221608f
C2733 a_100_23094# VSUBS 0.287142f
C2734 a_n158_23094# VSUBS 0.287142f
C2735 a_n100_22997# VSUBS 0.221608f
C2736 a_100_24530# VSUBS 0.287142f
C2737 a_n158_24530# VSUBS 0.287142f
C2738 a_n100_24433# VSUBS 0.221608f
C2739 a_100_25966# VSUBS 0.287142f
C2740 a_n158_25966# VSUBS 0.287142f
C2741 a_n100_25869# VSUBS 0.221608f
C2742 a_100_27402# VSUBS 0.287142f
C2743 a_n158_27402# VSUBS 0.287142f
C2744 a_n100_27305# VSUBS 0.221608f
C2745 a_100_28838# VSUBS 0.287142f
C2746 a_n158_28838# VSUBS 0.287142f
C2747 a_n100_28741# VSUBS 0.221608f
C2748 a_100_30274# VSUBS 0.287142f
C2749 a_n158_30274# VSUBS 0.287142f
C2750 a_n100_30177# VSUBS 0.221608f
C2751 a_100_31710# VSUBS 0.287142f
C2752 a_n158_31710# VSUBS 0.287142f
C2753 a_n100_31613# VSUBS 0.221608f
C2754 a_100_33146# VSUBS 0.287142f
C2755 a_n158_33146# VSUBS 0.287142f
C2756 a_n100_33049# VSUBS 0.221608f
C2757 a_100_34582# VSUBS 0.287142f
C2758 a_n158_34582# VSUBS 0.287142f
C2759 a_n100_34485# VSUBS 0.221608f
C2760 a_100_36018# VSUBS 0.287142f
C2761 a_n158_36018# VSUBS 0.287142f
C2762 a_n100_35921# VSUBS 0.221608f
C2763 a_100_37454# VSUBS 0.287142f
C2764 a_n158_37454# VSUBS 0.287142f
C2765 a_n100_37357# VSUBS 0.221608f
C2766 a_100_38890# VSUBS 0.287142f
C2767 a_n158_38890# VSUBS 0.287142f
C2768 a_n100_38793# VSUBS 0.221608f
C2769 a_100_40326# VSUBS 0.287142f
C2770 a_n158_40326# VSUBS 0.287142f
C2771 a_n100_40229# VSUBS 0.221608f
C2772 a_100_41762# VSUBS 0.287142f
C2773 a_n158_41762# VSUBS 0.287142f
C2774 a_n100_41665# VSUBS 0.221608f
C2775 a_100_43198# VSUBS 0.287142f
C2776 a_n158_43198# VSUBS 0.287142f
C2777 a_n100_43101# VSUBS 0.221608f
C2778 a_100_44634# VSUBS 0.287142f
C2779 a_n158_44634# VSUBS 0.287142f
C2780 a_n100_44537# VSUBS 0.221608f
C2781 a_100_46070# VSUBS 0.287142f
C2782 a_n158_46070# VSUBS 0.287142f
C2783 a_n100_45973# VSUBS 0.221608f
C2784 a_100_47506# VSUBS 0.287142f
C2785 a_n158_47506# VSUBS 0.287142f
C2786 a_n100_47409# VSUBS 0.221608f
C2787 a_100_48942# VSUBS 0.287142f
C2788 a_n158_48942# VSUBS 0.287142f
C2789 a_n100_48845# VSUBS 0.221608f
C2790 a_100_50378# VSUBS 0.287142f
C2791 a_n158_50378# VSUBS 0.287142f
C2792 a_n100_50281# VSUBS 0.221608f
C2793 a_100_51814# VSUBS 0.287142f
C2794 a_n158_51814# VSUBS 0.287142f
C2795 a_n100_51717# VSUBS 0.221608f
C2796 a_100_53250# VSUBS 0.287142f
C2797 a_n158_53250# VSUBS 0.287142f
C2798 a_n100_53153# VSUBS 0.221608f
C2799 a_100_54686# VSUBS 0.287142f
C2800 a_n158_54686# VSUBS 0.287142f
C2801 a_n100_54589# VSUBS 0.221608f
C2802 a_100_56122# VSUBS 0.287142f
C2803 a_n158_56122# VSUBS 0.287142f
C2804 a_n100_56025# VSUBS 0.221608f
C2805 a_100_57558# VSUBS 0.287142f
C2806 a_n158_57558# VSUBS 0.287142f
C2807 a_n100_57461# VSUBS 0.221608f
C2808 a_100_58994# VSUBS 0.287142f
C2809 a_n158_58994# VSUBS 0.287142f
C2810 a_n100_58897# VSUBS 0.221608f
C2811 a_100_60430# VSUBS 0.287142f
C2812 a_n158_60430# VSUBS 0.287142f
C2813 a_n100_60333# VSUBS 0.221608f
C2814 a_100_61866# VSUBS 0.287142f
C2815 a_n158_61866# VSUBS 0.287142f
C2816 a_n100_61769# VSUBS 0.221608f
C2817 a_100_63302# VSUBS 0.287142f
C2818 a_n158_63302# VSUBS 0.287142f
C2819 a_n100_63205# VSUBS 0.221608f
C2820 a_100_64738# VSUBS 0.287142f
C2821 a_n158_64738# VSUBS 0.287142f
C2822 a_n100_64641# VSUBS 0.221608f
C2823 a_100_66174# VSUBS 0.287142f
C2824 a_n158_66174# VSUBS 0.287142f
C2825 a_n100_66077# VSUBS 0.221608f
C2826 a_100_67610# VSUBS 0.287142f
C2827 a_n158_67610# VSUBS 0.287142f
C2828 a_n100_67513# VSUBS 0.221608f
C2829 a_100_69046# VSUBS 0.287142f
C2830 a_n158_69046# VSUBS 0.287142f
C2831 a_n100_68949# VSUBS 0.221608f
C2832 a_100_70482# VSUBS 0.287142f
C2833 a_n158_70482# VSUBS 0.287142f
C2834 a_n100_70385# VSUBS 0.221608f
C2835 a_100_71918# VSUBS 0.287142f
C2836 a_n158_71918# VSUBS 0.287142f
C2837 a_n100_71821# VSUBS 0.221608f
C2838 a_100_73354# VSUBS 0.287142f
C2839 a_n158_73354# VSUBS 0.287142f
C2840 a_n100_73257# VSUBS 0.221608f
C2841 a_100_74790# VSUBS 0.287142f
C2842 a_n158_74790# VSUBS 0.287142f
C2843 a_n100_74693# VSUBS 0.221608f
C2844 a_100_76226# VSUBS 0.287142f
C2845 a_n158_76226# VSUBS 0.287142f
C2846 a_n100_76129# VSUBS 0.221608f
C2847 a_100_77662# VSUBS 0.287142f
C2848 a_n158_77662# VSUBS 0.287142f
C2849 a_n100_77565# VSUBS 0.221608f
C2850 a_100_79098# VSUBS 0.287142f
C2851 a_n158_79098# VSUBS 0.287142f
C2852 a_n100_79001# VSUBS 0.221608f
C2853 a_100_80534# VSUBS 0.287142f
C2854 a_n158_80534# VSUBS 0.287142f
C2855 a_n100_80437# VSUBS 0.221608f
C2856 a_100_81970# VSUBS 0.287142f
C2857 a_n158_81970# VSUBS 0.287142f
C2858 a_n100_81873# VSUBS 0.221608f
C2859 a_100_83406# VSUBS 0.287142f
C2860 a_n158_83406# VSUBS 0.287142f
C2861 a_n100_83309# VSUBS 0.221608f
C2862 a_100_84842# VSUBS 0.287142f
C2863 a_n158_84842# VSUBS 0.287142f
C2864 a_n100_84745# VSUBS 0.221608f
C2865 a_100_86278# VSUBS 0.287142f
C2866 a_n158_86278# VSUBS 0.287142f
C2867 a_n100_86181# VSUBS 0.221608f
C2868 a_100_87714# VSUBS 0.287142f
C2869 a_n158_87714# VSUBS 0.287142f
C2870 a_n100_87617# VSUBS 0.221608f
C2871 a_100_89150# VSUBS 0.287142f
C2872 a_n158_89150# VSUBS 0.287142f
C2873 a_n100_89053# VSUBS 0.221608f
C2874 a_100_90586# VSUBS 0.287142f
C2875 a_n158_90586# VSUBS 0.287142f
C2876 a_n100_90489# VSUBS 0.221608f
C2877 a_100_92022# VSUBS 0.287142f
C2878 a_n158_92022# VSUBS 0.287142f
C2879 a_n100_91925# VSUBS 0.221608f
C2880 a_100_93458# VSUBS 0.287142f
C2881 a_n158_93458# VSUBS 0.287142f
C2882 a_n100_93361# VSUBS 0.221608f
C2883 a_100_94894# VSUBS 0.287142f
C2884 a_n158_94894# VSUBS 0.287142f
C2885 a_n100_94797# VSUBS 0.221608f
C2886 a_100_96330# VSUBS 0.287142f
C2887 a_n158_96330# VSUBS 0.287142f
C2888 a_n100_96233# VSUBS 0.221608f
C2889 a_100_97766# VSUBS 0.287142f
C2890 a_n158_97766# VSUBS 0.287142f
C2891 a_n100_97669# VSUBS 0.221608f
C2892 a_100_99202# VSUBS 0.287142f
C2893 a_n158_99202# VSUBS 0.287142f
C2894 a_n100_99105# VSUBS 0.221608f
C2895 a_100_100638# VSUBS 0.287142f
C2896 a_n158_100638# VSUBS 0.287142f
C2897 a_n100_100541# VSUBS 0.221608f
C2898 a_100_102074# VSUBS 0.287142f
C2899 a_n158_102074# VSUBS 0.287142f
C2900 a_n100_101977# VSUBS 0.221608f
C2901 a_100_103510# VSUBS 0.287142f
C2902 a_n158_103510# VSUBS 0.287142f
C2903 a_n100_103413# VSUBS 0.221608f
C2904 a_100_104946# VSUBS 0.287142f
C2905 a_n158_104946# VSUBS 0.287142f
C2906 a_n100_104849# VSUBS 0.221608f
C2907 a_100_106382# VSUBS 0.287142f
C2908 a_n158_106382# VSUBS 0.287142f
C2909 a_n100_106285# VSUBS 0.221608f
C2910 a_100_107818# VSUBS 0.287142f
C2911 a_n158_107818# VSUBS 0.287142f
C2912 a_n100_107721# VSUBS 0.221608f
C2913 a_100_109254# VSUBS 0.287142f
C2914 a_n158_109254# VSUBS 0.287142f
C2915 a_n100_109157# VSUBS 0.221608f
C2916 a_100_110690# VSUBS 0.287142f
C2917 a_n158_110690# VSUBS 0.287142f
C2918 a_n100_110593# VSUBS 0.221608f
C2919 a_100_112126# VSUBS 0.287142f
C2920 a_n158_112126# VSUBS 0.287142f
C2921 a_n100_112029# VSUBS 0.221608f
C2922 a_100_113562# VSUBS 0.287142f
C2923 a_n158_113562# VSUBS 0.287142f
C2924 a_n100_113465# VSUBS 0.221608f
C2925 a_100_114998# VSUBS 0.287142f
C2926 a_n158_114998# VSUBS 0.287142f
C2927 a_n100_114901# VSUBS 0.221608f
C2928 a_100_116434# VSUBS 0.287142f
C2929 a_n158_116434# VSUBS 0.287142f
C2930 a_n100_116337# VSUBS 0.221608f
C2931 a_100_117870# VSUBS 0.287142f
C2932 a_n158_117870# VSUBS 0.287142f
C2933 a_n100_117773# VSUBS 0.221608f
C2934 a_100_119306# VSUBS 0.287142f
C2935 a_n158_119306# VSUBS 0.287142f
C2936 a_n100_119209# VSUBS 0.221608f
C2937 a_100_120742# VSUBS 0.287142f
C2938 a_n158_120742# VSUBS 0.287142f
C2939 a_n100_120645# VSUBS 0.221608f
C2940 a_100_122178# VSUBS 0.287142f
C2941 a_n158_122178# VSUBS 0.287142f
C2942 a_n100_122081# VSUBS 0.221608f
C2943 a_100_123614# VSUBS 0.287142f
C2944 a_n158_123614# VSUBS 0.287142f
C2945 a_n100_123517# VSUBS 0.221608f
C2946 a_100_125050# VSUBS 0.287142f
C2947 a_n158_125050# VSUBS 0.287142f
C2948 a_n100_124953# VSUBS 0.221608f
C2949 a_100_126486# VSUBS 0.287142f
C2950 a_n158_126486# VSUBS 0.287142f
C2951 a_n100_126389# VSUBS 0.221608f
C2952 a_100_127922# VSUBS 0.287142f
C2953 a_n158_127922# VSUBS 0.287142f
C2954 a_n100_127825# VSUBS 0.221608f
C2955 a_100_129358# VSUBS 0.287142f
C2956 a_n158_129358# VSUBS 0.287142f
C2957 a_n100_129261# VSUBS 0.221608f
C2958 a_100_130794# VSUBS 0.287142f
C2959 a_n158_130794# VSUBS 0.287142f
C2960 a_n100_130697# VSUBS 0.221608f
C2961 a_100_132230# VSUBS 0.287142f
C2962 a_n158_132230# VSUBS 0.287142f
C2963 a_n100_132133# VSUBS 0.221608f
C2964 a_100_133666# VSUBS 0.287142f
C2965 a_n158_133666# VSUBS 0.287142f
C2966 a_n100_133569# VSUBS 0.221608f
C2967 a_100_135102# VSUBS 0.287142f
C2968 a_n158_135102# VSUBS 0.287142f
C2969 a_n100_135005# VSUBS 0.221608f
C2970 a_100_136538# VSUBS 0.287142f
C2971 a_n158_136538# VSUBS 0.287142f
C2972 a_n100_136441# VSUBS 0.221608f
C2973 a_100_137974# VSUBS 0.287142f
C2974 a_n158_137974# VSUBS 0.287142f
C2975 a_n100_137877# VSUBS 0.221608f
C2976 a_100_139410# VSUBS 0.287142f
C2977 a_n158_139410# VSUBS 0.287142f
C2978 a_n100_139313# VSUBS 0.221608f
C2979 a_100_140846# VSUBS 0.287142f
C2980 a_n158_140846# VSUBS 0.287142f
C2981 a_n100_140749# VSUBS 0.221608f
C2982 a_100_142282# VSUBS 0.287142f
C2983 a_n158_142282# VSUBS 0.287142f
C2984 a_n100_142185# VSUBS 0.221608f
C2985 a_100_143718# VSUBS 0.287142f
C2986 a_n158_143718# VSUBS 0.287142f
C2987 a_n100_143621# VSUBS 0.221608f
C2988 a_100_145154# VSUBS 0.287142f
C2989 a_n158_145154# VSUBS 0.287142f
C2990 a_n100_145057# VSUBS 0.221608f
C2991 a_100_146590# VSUBS 0.287142f
C2992 a_n158_146590# VSUBS 0.287142f
C2993 a_n100_146493# VSUBS 0.221608f
C2994 a_100_148026# VSUBS 0.287142f
C2995 a_n158_148026# VSUBS 0.287142f
C2996 a_n100_147929# VSUBS 0.221608f
C2997 a_100_149462# VSUBS 0.287142f
C2998 a_n158_149462# VSUBS 0.287142f
C2999 a_n100_149365# VSUBS 0.221608f
C3000 a_100_150898# VSUBS 0.287142f
C3001 a_n158_150898# VSUBS 0.287142f
C3002 a_n100_150801# VSUBS 0.221608f
C3003 a_100_152334# VSUBS 0.287142f
C3004 a_n158_152334# VSUBS 0.287142f
C3005 a_n100_152237# VSUBS 0.221608f
C3006 a_100_153770# VSUBS 0.287142f
C3007 a_n158_153770# VSUBS 0.287142f
C3008 a_n100_153673# VSUBS 0.221608f
C3009 a_100_155206# VSUBS 0.287142f
C3010 a_n158_155206# VSUBS 0.287142f
C3011 a_n100_155109# VSUBS 0.221608f
C3012 a_100_156642# VSUBS 0.287142f
C3013 a_n158_156642# VSUBS 0.287142f
C3014 a_n100_156545# VSUBS 0.221608f
C3015 a_100_158078# VSUBS 0.287142f
C3016 a_n158_158078# VSUBS 0.287142f
C3017 a_n100_157981# VSUBS 0.221608f
C3018 a_100_159514# VSUBS 0.287142f
C3019 a_n158_159514# VSUBS 0.287142f
C3020 a_n100_159417# VSUBS 0.221608f
C3021 a_100_160950# VSUBS 0.287142f
C3022 a_n158_160950# VSUBS 0.287142f
C3023 a_n100_160853# VSUBS 0.221608f
C3024 a_100_162386# VSUBS 0.287142f
C3025 a_n158_162386# VSUBS 0.287142f
C3026 a_n100_162289# VSUBS 0.221608f
C3027 a_100_163822# VSUBS 0.287142f
C3028 a_n158_163822# VSUBS 0.287142f
C3029 a_n100_163725# VSUBS 0.221608f
C3030 a_100_165258# VSUBS 0.287142f
C3031 a_n158_165258# VSUBS 0.287142f
C3032 a_n100_165161# VSUBS 0.221608f
C3033 a_100_166694# VSUBS 0.287142f
C3034 a_n158_166694# VSUBS 0.287142f
C3035 a_n100_166597# VSUBS 0.221608f
C3036 a_100_168130# VSUBS 0.287142f
C3037 a_n158_168130# VSUBS 0.287142f
C3038 a_n100_168033# VSUBS 0.221608f
C3039 a_100_169566# VSUBS 0.287142f
C3040 a_n158_169566# VSUBS 0.287142f
C3041 a_n100_169469# VSUBS 0.221608f
C3042 a_100_171002# VSUBS 0.287142f
C3043 a_n158_171002# VSUBS 0.287142f
C3044 a_n100_170905# VSUBS 0.221608f
C3045 a_100_172438# VSUBS 0.287142f
C3046 a_n158_172438# VSUBS 0.287142f
C3047 a_n100_172341# VSUBS 0.221608f
C3048 a_100_173874# VSUBS 0.287142f
C3049 a_n158_173874# VSUBS 0.287142f
C3050 a_n100_173777# VSUBS 0.221608f
C3051 a_100_175310# VSUBS 0.287142f
C3052 a_n158_175310# VSUBS 0.287142f
C3053 a_n100_175213# VSUBS 0.221608f
C3054 a_100_176746# VSUBS 0.287142f
C3055 a_n158_176746# VSUBS 0.287142f
C3056 a_n100_176649# VSUBS 0.221608f
C3057 a_100_178182# VSUBS 0.287142f
C3058 a_n158_178182# VSUBS 0.287142f
C3059 a_n100_178085# VSUBS 0.221608f
C3060 a_100_179618# VSUBS 0.287142f
C3061 a_n158_179618# VSUBS 0.287142f
C3062 a_n100_179521# VSUBS 0.221608f
C3063 a_100_181054# VSUBS 0.287142f
C3064 a_n158_181054# VSUBS 0.287142f
C3065 a_n100_180957# VSUBS 0.221608f
C3066 a_100_182490# VSUBS 0.292592f
C3067 a_n158_182490# VSUBS 0.292592f
C3068 a_n100_182393# VSUBS 0.265338f
C3069 w_n358_n183987# VSUBS 0.982325p
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_AJ8KYZ a_n100_n42155# a_100_n252938# a_n158_26478#
+ a_n100_n226675# a_n158_n268754# a_n100_n181863# a_n100_n21067# a_n100_n205587# a_n158_n247666#
+ a_n100_n160775# a_n158_n5154# a_n100_n324207# a_100_n334654# a_n100_n308391# a_n100_10565#
+ a_n158_n226578# a_n158_n181766# a_100_n47330# a_n100_n303119# a_100_n107958# a_100_n313566#
+ a_n158_n78962# a_n158_n329382# a_n100_n242491# a_n158_n284570# a_100_13298# a_n158_n160678#
+ a_100_n26242# a_n100_n155503# a_100_n165950# a_n158_n308294# a_n158_n57874# a_n158_n263482#
+ a_n100_n134415# a_100_29114# a_n158_n36786# a_100_n144862# a_n158_n242394# a_n100_n184499#
+ a_n100_n113327# a_n158_n15698# a_100_n123774# a_n158_n155406# a_n158_n139590# a_n100_n57971#
+ a_n100_n216131# a_n158_n258210# a_n158_n134318# a_n158_n73690# a_100_n102686# a_100_n292478#
+ a_n100_n36883# a_100_n221306# a_100_n205490# a_n158_n237122# a_n100_n150231# a_n100_n179227#
+ a_100_n189674# a_n158_n192310# a_n100_n7887# a_n100_n15795# a_100_n118502# a_100_n324110#
+ a_100_n200218# a_n158_n216034# a_n100_29017# a_n100_n158139# a_n158_n171222# a_100_n168586#
+ a_n100_7929# a_n100_n318935# a_100_n303022# a_100_n287206# a_n158_n150134# a_100_n147498#
+ a_n158_n310930# a_n158_n47330# a_100_n266118# a_n100_n195043# a_n158_n26242# a_n158_n318838#
+ a_n158_2754# a_100_n7790# a_n100_n231947# a_100_n2518# a_100_n113230# a_n100_n334751#
+ a_n100_n210859# a_n158_n252938# a_n100_2657# a_n100_n313663# a_n100_n297847# a_100_n52602#
+ a_n100_n92239# a_100_n179130# a_n158_n334654# a_n100_n276759# a_100_n31514# a_n158_n107958#
+ a_100_n158042# a_n158_n313566# a_100_n81598# a_100_n10426# a_100_18570# a_n100_n123871#
+ a_n158_n165950# a_100_n97414# a_n100_n102783# a_n158_n144862# a_n100_n337387# a_n100_n292575#
+ a_100_n76326# a_n100_n221403# a_n158_21206# a_100_n231850# a_n100_n316299# a_n158_n123774#
+ a_n100_n189771# a_n100_n271487# a_100_n55238# a_n100_n200315# a_100_n210762# a_100_n239758#
+ a_n158_n102686# a_n100_n168683# a_100_n194946# a_n100_n250399# a_n158_n292478# a_100_5390#
+ a_n158_118# a_n158_n221306# a_n158_n205490# a_100_n297750# a_n100_n287303# a_n100_18473#
+ a_100_n173858# a_n100_n147595# a_n158_n189674# a_n100_21# a_n158_n118502# a_n158_n324110#
+ a_100_n92142# a_n158_n200218# a_n100_n266215# a_100_n276662# a_n158_n168586# a_n100_n86967#
+ a_n158_n52602# a_n158_n303022# a_100_n71054# a_n100_n245127# a_n158_n287206# a_100_n255574#
+ a_n158_n147498# a_n100_n65879# a_n158_n31514# a_n100_n224039# a_n158_n266118# a_100_n234486#
+ a_n158_n81598# a_n158_n10426# a_100_n337290# a_100_n213398# a_n100_n282031# a_100_n332018#
+ a_n158_n97414# a_n158_n113230# a_n100_n31611# a_100_n271390# a_n100_n81695# a_100_n229214#
+ a_n158_15934# a_n158_n76326# a_100_n184402# a_n100_n2615# a_n100_n10523# a_n100_n39519#
+ a_100_n279298# a_100_n20970# a_100_n49966# a_100_n208126# a_100_n163314# a_n158_n55238#
+ a_n100_n137051# a_n158_n179130# a_n100_n97511# a_100_n28878# a_100_n142226# a_100_23842#
+ a_n158_n158042# a_n100_n76423# a_100_n86870# a_100_n245030# a_100_n121138# a_n158_n92142#
+ a_n100_n55335# a_n158_10662# a_100_n65782# a_n100_n239855# a_n158_n71054# a_n100_n34247#
+ a_100_n44694# a_n100_n218767# a_n158_n231850# a_n100_n173955# a_100_n187038# a_n100_n13159#
+ a_n158_n210762# a_n158_n239758# a_n100_23745# a_n100_n152867# a_n158_n194946# a_n100_n71151#
+ a_100_n326746# a_100_n281934# a_n158_n297750# a_n100_n255671# a_100_26478# a_n100_n131779#
+ a_n158_n173858# w_n358_n337587# a_n100_n50063# a_n100_n79059# a_100_n39422# a_100_n305658#
+ a_n158_5390# a_100_n260846# a_n100_n234583# a_n158_n276662# a_100_n18334# a_100_n5154#
+ a_n158_n20970# a_n158_n49966# a_n158_13298# a_n100_n213495# a_n158_n255574# a_n100_n197679#
+ a_n100_n126507# a_n100_n332115# a_n158_n28878# a_100_n136954# a_n100_5293# a_n158_n234486#
+ a_n158_29114# a_n100_n229311# a_n100_n105419# a_n100_n311027# a_100_n115866# a_100_n321474#
+ a_n158_n86870# a_n158_n213398# a_n158_n337290# a_n100_n279395# a_100_n34150# a_n100_n208223#
+ a_n100_n163411# a_100_n218670# a_n158_n332018# a_100_n300386# a_n158_n65782# a_n100_n28975#
+ a_n158_n271390# a_100_n13062# a_n158_n229214# a_n100_13201# a_n100_n142323# a_n158_n44694#
+ a_100_n152770# a_n158_n184402# a_100_8026# a_n158_n279298# a_100_n316202# a_n158_n208126#
+ a_n100_n121235# a_n158_n163314# a_100_n131682# a_100_n250302# a_n100_n100147# a_100_n110594#
+ a_n158_n142226# a_n100_n60607# a_n100_n44791# a_n158_n39422# a_n158_n245030# a_n158_n121138#
+ a_n100_n187135# a_100_n197582# a_n158_n18334# a_100_n126410# a_n100_n166047# a_100_n176494#
+ a_n158_n7790# a_100_n105322# a_n100_n326843# a_100_n295114# a_n158_n187038# a_n158_n2518#
+ a_n100_n305755# a_100_n274026# a_n100_n260943# a_n100_n18431# a_n100_n289939# a_n158_n34150#
+ a_n158_n326746# a_100_n94778# a_n158_n281934# a_100_n23606# a_n158_n13062# a_n158_n305658#
+ a_n158_n260846# a_100_n100050# a_n100_n115963# a_100_n129046# a_n100_n321571# a_100_n60510#
+ a_100_n89506# a_n158_18570# a_n100_n300483# a_n158_n136954# a_n100_n329479# a_n100_n284667#
+ a_n100_n5251# a_100_n68418# a_100_n223942# a_n158_n115866# a_n158_n321474# a_n100_n263579#
+ a_100_n202854# a_n158_n218670# a_n158_n300386# a_100_n289842# a_100_21206# a_n100_n110691#
+ a_n100_n139687# a_n158_n152770# a_n158_n316202# a_100_n84234# a_100_n268754# a_n100_n258307#
+ a_n100_n118599# a_n158_n131682# a_n158_8026# a_100_n63146# a_n100_n237219# a_n158_n250302#
+ a_100_n247666# a_n100_n192407# a_n158_n94778# a_n158_n110594# a_n100_n176591# a_n158_n23606#
+ a_100_n42058# a_100_n226578# a_n100_n295211# a_n100_26381# a_n100_n171319# a_100_n181766#
+ a_n158_n197582# a_n158_n126410# a_100_n329382# a_n100_n274123# a_n100_21109# a_100_n284570#
+ a_100_n160678# a_100_118# a_n158_n176494# a_n100_n94875# a_n158_n60510# a_n158_n89506#
+ a_n158_n105322# a_100_n308294# a_n100_n253035# a_n158_n295114# a_n100_n23703# a_100_n263482#
+ a_n100_n73787# a_n158_n68418# a_n158_n274026# a_100_n242394# a_n100_n52699# a_100_n155406#
+ a_n100_n129143# a_100_n139590# a_n100_n89603# a_100_n258210# a_100_n134318# a_100_15934#
+ a_n100_n108055# a_n100_n68515# a_n158_23842# a_100_n78962# a_100_n237122# a_100_n192310#
+ a_n158_n84234# a_n158_n100050# a_n158_n129046# a_n100_n47427# a_100_n57874# a_n100_n202951#
+ a_100_n216034# a_100_n171222# a_n158_n63146# a_n100_n26339# a_100_n36786# a_n158_n223942#
+ a_n158_n42058# a_100_n150134# a_100_2754# a_n100_n84331# a_100_n310930# a_100_n15698#
+ a_n158_n202854# a_n100_n268851# a_100_10662# a_n100_15837# a_n100_n144959# a_n100_n63243#
+ VSUBS a_100_n318838# a_100_n73690# a_n100_n247763# a_n158_n289842#
X0 a_100_213634# a_n100_213537# a_n158_213634# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X1 a_100_42294# a_n100_42197# a_n158_42294# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X2 a_100_n115866# a_n100_n115963# a_n158_n115866# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X3 a_100_n184402# a_n100_n184499# a_n158_n184402# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X4 a_100_253174# a_n100_253077# a_n158_253174# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X5 a_100_n36786# a_n100_n36883# a_n158_n36786# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X6 a_100_305894# a_n100_305797# a_n158_305894# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X7 a_100_15934# a_n100_15837# a_n158_15934# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X8 a_100_n7790# a_n100_n7887# a_n158_n7790# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X9 a_100_n276662# a_n100_n276759# a_n158_n276662# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X10 a_100_105558# a_n100_105461# a_n158_105558# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X11 a_100_226814# a_n100_226717# a_n158_226814# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X12 a_100_n324110# a_n100_n324207# a_n158_n324110# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X13 a_100_n321474# a_n100_n321571# a_n158_n321474# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X14 a_100_n237122# a_n100_n237219# a_n158_n237122# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X15 a_100_n160678# a_n100_n160775# a_n158_n160678# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X16 a_100_55474# a_n100_55377# a_n158_55474# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X17 a_100_n281934# a_n100_n282031# a_n158_n281934# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X18 a_100_145098# a_n100_145001# a_n158_145098# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X19 a_100_n81598# a_n100_n81695# a_n158_n81598# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X20 a_100_n121138# a_n100_n121235# a_n158_n121138# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X21 a_100_266354# a_n100_266257# a_n158_266354# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X22 a_100_n49966# a_n100_n50063# a_n158_n49966# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X23 a_100_60746# a_n100_60649# a_n158_60746# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X24 a_100_n42058# a_n100_n42155# a_n158_n42058# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X25 a_100_n329382# a_n100_n329479# a_n158_n329382# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X26 a_100_n168586# a_n100_n168683# a_n158_n168586# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X27 a_100_n289842# a_n100_n289939# a_n158_n289842# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X28 a_100_311166# a_n100_311069# a_n158_311166# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X29 a_100_21206# a_n100_21109# a_n158_21206# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X30 a_100_n213398# a_n100_n213495# a_n158_n213398# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X31 a_100_271626# a_n100_271529# a_n158_271626# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X32 a_100_118738# a_n100_118641# a_n158_118738# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X33 a_100_n129046# a_n100_n129143# a_n158_n129046# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X34 a_100_n334654# a_n100_n334751# a_n158_n334654# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X35 a_100_n173858# a_n100_n173955# a_n158_n173858# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X36 a_100_68654# a_n100_68557# a_n158_68654# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X37 a_100_319074# a_n100_318977# a_n158_319074# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X38 a_100_n134318# a_n100_n134415# a_n158_n134318# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X39 a_100_n131682# a_n100_n131779# a_n158_n131682# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X40 a_100_n94778# a_n100_n94875# a_n158_n94778# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X41 a_100_158278# a_n100_158181# a_n158_158278# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X42 a_100_29114# a_n100_29017# a_n158_29114# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X43 a_100_279534# a_n100_279437# a_n158_279534# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X44 a_100_73926# a_n100_73829# a_n158_73926# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X45 a_100_n55238# a_n100_n55335# a_n158_n55238# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X46 a_100_324346# a_n100_324249# a_n158_324346# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X47 a_100_118# a_n100_21# a_n158_118# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X48 a_100_31750# a_n100_31653# a_n158_31750# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X49 a_100_n13062# a_n100_n13159# a_n158_n13062# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X50 a_100_n295114# a_n100_n295211# a_n158_n295114# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X51 a_100_n226578# a_n100_n226675# a_n158_n226578# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X52 a_100_284806# a_n100_284709# a_n158_284806# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X53 a_100_121374# a_n100_121277# a_n158_121374# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X54 a_100_n60510# a_n100_n60607# a_n158_n60510# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X55 a_100_242630# a_n100_242533# a_n158_242630# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X56 a_100_71290# a_n100_71193# a_n158_71290# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X57 a_100_n231850# a_n100_n231947# a_n158_n231850# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X58 a_100_n144862# a_n100_n144959# a_n158_n144862# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X59 a_100_n65782# a_n100_n65879# a_n158_n65782# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X60 a_100_n105322# a_n100_n105419# a_n158_n105322# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X61 a_100_334890# a_n100_334793# a_n158_334890# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X62 a_100_282170# a_n100_282073# a_n158_282170# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X63 a_100_129282# a_n100_129185# a_n158_129282# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X64 a_100_n68418# a_n100_n68515# a_n158_n68418# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X65 a_100_44930# a_n100_44833# a_n158_44930# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X66 a_100_n271390# a_n100_n271487# a_n158_n271390# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X67 a_100_n187038# a_n100_n187135# a_n158_n187038# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X68 a_100_n26242# a_n100_n26339# a_n158_n26242# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X69 a_100_n239758# a_n100_n239855# a_n158_n239758# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X70 a_100_134554# a_n100_134457# a_n158_134554# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X71 a_100_255810# a_n100_255713# a_n158_255810# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X72 a_100_84470# a_n100_84373# a_n158_84470# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X73 a_100_n192310# a_n100_n192407# a_n158_n192310# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X74 a_100_87106# a_n100_87009# a_n158_87106# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X75 a_100_n31514# a_n100_n31611# a_n158_n31514# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X76 a_100_n279298# a_n100_n279395# a_n158_n279298# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X77 a_100_300622# a_n100_300525# a_n158_300622# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X78 a_100_174094# a_n100_173997# a_n158_174094# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X79 a_100_n2518# a_n100_n2615# a_n158_n2518# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X80 a_100_n150134# a_n100_n150231# a_n158_n150134# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X81 a_100_295350# a_n100_295253# a_n158_295350# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X82 a_100_n78962# a_n100_n79059# a_n158_n78962# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X83 a_100_n202854# a_n100_n202951# a_n158_n202854# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X84 a_100_n118502# a_n100_n118599# a_n158_n118502# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X85 a_100_n71054# a_n100_n71151# a_n158_n71054# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X86 a_100_n284570# a_n100_n284667# a_n158_n284570# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X87 a_100_n197582# a_n100_n197679# a_n158_n197582# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X88 a_100_n39422# a_n100_n39519# a_n158_n39422# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X89 a_100_308530# a_n100_308433# a_n158_308530# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X90 a_100_147734# a_n100_147637# a_n158_147734# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X91 a_100_50202# a_n100_50105# a_n158_50202# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X92 a_100_n245030# a_n100_n245127# a_n158_n245030# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X93 a_100_n242394# a_n100_n242491# a_n158_n242394# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X94 a_100_n158042# a_n100_n158139# a_n158_n158042# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X95 a_100_97650# a_n100_97553# a_n158_97650# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X96 a_100_313802# a_n100_313705# a_n158_313802# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X97 a_100_187274# a_n100_187177# a_n158_187274# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X98 a_100_n163314# a_n100_n163411# a_n158_n163314# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X99 a_100_239994# a_n100_239897# a_n158_239994# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X100 a_100_58110# a_n100_58013# a_n158_58110# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X101 a_100_n337290# a_n100_n337387# a_n158_n337290# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X102 a_100_232086# a_n100_231989# a_n158_232086# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X103 a_100_110830# a_n100_110733# a_n158_110830# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X104 a_100_n15698# a_n100_n15795# a_n158_n15698# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X105 a_100_n84234# a_n100_n84331# a_n158_n84234# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X106 a_100_n297750# a_n100_n297847# a_n158_n297750# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X107 a_100_192546# a_n100_192449# a_n158_192546# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X108 a_100_n255574# a_n100_n255671# a_n158_n255574# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X109 a_100_n258210# a_n100_n258307# a_n158_n258210# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X110 a_100_153006# a_n100_152909# a_n158_153006# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X111 a_100_150370# a_n100_150273# a_n158_150370# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X112 a_100_n20970# a_n100_n21067# a_n158_n20970# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X113 a_100_205726# a_n100_205629# a_n158_205726# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X114 a_100_n300386# a_n100_n300483# a_n158_n300386# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X115 a_100_n216034# a_n100_n216131# a_n158_n216034# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X116 a_100_34386# a_n100_34289# a_n158_34386# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X117 a_100_n260846# a_n100_n260943# a_n158_n260846# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X118 a_100_n107958# a_n100_n108055# a_n158_n107958# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X119 a_100_n100050# a_n100_n100147# a_n158_n100050# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X120 a_100_245266# a_n100_245169# a_n158_245266# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X121 a_100_n28878# a_n100_n28975# a_n158_n28878# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X122 a_100_n221306# a_n100_n221403# a_n158_n221306# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X123 a_100_n97414# a_n100_n97511# a_n158_n97414# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X124 a_100_n308294# a_n100_n308391# a_n158_n308294# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X125 a_100_n147498# a_n100_n147595# a_n158_n147498# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X126 a_100_203090# a_n100_202993# a_n158_203090# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X127 a_100_n268754# a_n100_n268851# a_n158_n268754# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X128 a_100_250538# a_n100_250441# a_n158_250538# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X129 a_100_163550# a_n100_163453# a_n158_163550# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X130 a_100_5390# a_n100_5293# a_n158_5390# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X131 a_100_218906# a_n100_218809# a_n158_218906# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X132 a_100_8026# a_n100_7929# a_n158_8026# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X133 a_100_n313566# a_n100_n313663# a_n158_n313566# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X134 a_100_n229214# a_n100_n229311# a_n158_n229214# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X135 a_100_n152770# a_n100_n152867# a_n158_n152770# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X136 a_100_297986# a_n100_297889# a_n158_297986# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X137 a_100_124010# a_n100_123913# a_n158_124010# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X138 a_100_47566# a_n100_47469# a_n158_47566# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X139 a_100_n73690# a_n100_n73787# a_n158_n73690# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X140 a_100_n113230# a_n100_n113327# a_n158_n113230# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X141 a_100_n110594# a_n100_n110691# a_n158_n110594# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X142 a_100_290078# a_n100_289981# a_n158_290078# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X143 a_100_258446# a_n100_258349# a_n158_258446# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X144 a_100_52838# a_n100_52741# a_n158_52838# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X145 a_100_n34150# a_n100_n34247# a_n158_n34150# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X146 a_100_303258# a_n100_303161# a_n158_303258# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X147 a_100_216270# a_n100_216173# a_n158_216270# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X148 a_100_176730# a_n100_176633# a_n158_176730# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X149 a_100_10662# a_n100_10565# a_n158_10662# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X150 a_100_n274026# a_n100_n274123# a_n158_n274026# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X151 a_100_n205490# a_n100_n205587# a_n158_n205490# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X152 a_100_263718# a_n100_263621# a_n158_263718# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X153 a_100_92378# a_n100_92281# a_n158_92378# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X154 a_100_n326746# a_n100_n326843# a_n158_n326746# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X155 a_100_100286# a_n100_100189# a_n158_100286# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X156 a_100_n165950# a_n100_n166047# a_n158_n165950# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X157 a_100_221542# a_n100_221445# a_n158_221542# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X158 a_100_n126410# a_n100_n126507# a_n158_n126410# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X159 a_100_n123774# a_n100_n123871# a_n158_n123774# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X160 a_100_n86870# a_n100_n86967# a_n158_n86870# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X161 a_100_268990# a_n100_268893# a_n158_268990# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X162 a_100_18570# a_n100_18473# a_n158_18570# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X163 a_100_n44694# a_n100_n44791# a_n158_n44694# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X164 a_100_261082# a_n100_260985# a_n158_261082# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X165 a_100_108194# a_n100_108097# a_n158_108194# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X166 a_100_n47330# a_n100_n47427# a_n158_n47330# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X167 a_100_316438# a_n100_316341# a_n158_316438# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X168 a_100_229450# a_n100_229353# a_n158_229450# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X169 a_100_23842# a_n100_23745# a_n158_23842# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X170 a_100_189910# a_n100_189813# a_n158_189910# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X171 a_100_n287206# a_n100_n287303# a_n158_n287206# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X172 a_100_n218670# a_n100_n218767# a_n158_n218670# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X173 a_100_113466# a_n100_113369# a_n158_113466# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X174 a_100_182002# a_n100_181905# a_n158_182002# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X175 a_100_234722# a_n100_234625# a_n158_234722# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X176 a_100_63382# a_n100_63285# a_n158_63382# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X177 a_100_n332018# a_n100_n332115# a_n158_n332018# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X178 a_100_n136954# a_n100_n137051# a_n158_n136954# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X179 a_100_66018# a_n100_65921# a_n158_66018# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X180 a_100_n10426# a_n100_n10523# a_n158_n10426# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X181 a_100_274262# a_n100_274165# a_n158_274262# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X182 a_100_n57874# a_n100_n57971# a_n158_n57874# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X183 a_100_n250302# a_n100_n250399# a_n158_n250302# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X184 a_100_326982# a_n100_326885# a_n158_326982# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X185 a_100_n176494# a_n100_n176591# a_n158_n176494# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X186 a_100_329618# a_n100_329521# a_n158_329618# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X187 a_100_n179130# a_n100_n179227# a_n158_n179130# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X188 a_100_n18334# a_n100_n18431# a_n158_n18334# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X189 a_100_210998# a_n100_210901# a_n158_210998# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X190 a_100_126646# a_n100_126549# a_n158_126646# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X191 a_100_247902# a_n100_247805# a_n158_247902# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X192 a_100_n181766# a_n100_n181863# a_n158_n181766# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X193 a_100_76562# a_n100_76465# a_n158_76562# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X194 a_100_n23606# a_n100_n23703# a_n158_n23606# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X195 a_100_n303022# a_n100_n303119# a_n158_n303022# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X196 a_100_166186# a_n100_166089# a_n158_166186# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X197 a_100_131918# a_n100_131821# a_n158_131918# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X198 a_100_n142226# a_n100_n142323# a_n158_n142226# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X199 a_100_287442# a_n100_287345# a_n158_287442# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X200 a_100_37022# a_n100_36925# a_n158_37022# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X201 a_100_81834# a_n100_81737# a_n158_81834# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X202 a_100_n63146# a_n100_n63243# a_n158_n63146# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X203 a_100_n189674# a_n100_n189771# a_n158_n189674# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X204 a_100_332254# a_n100_332157# a_n158_332254# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X205 a_100_171458# a_n100_171361# a_n158_171458# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X206 a_100_n234486# a_n100_n234583# a_n158_n234486# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X207 a_100_292714# a_n100_292617# a_n158_292714# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X208 a_100_139826# a_n100_139729# a_n158_139826# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X209 a_100_n194946# a_n100_n195043# a_n158_n194946# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X210 a_100_89742# a_n100_89645# a_n158_89742# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X211 a_100_13298# a_n100_13201# a_n158_13298# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X212 a_100_n316202# a_n100_n316299# a_n158_n316202# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X213 a_100_n155406# a_n100_n155503# a_n158_n155406# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X214 a_100_179366# a_n100_179269# a_n158_179366# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X215 a_100_224178# a_n100_224081# a_n158_224178# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X216 a_100_137190# a_n100_137093# a_n158_137190# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X217 a_100_102922# a_n100_102825# a_n158_102922# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X218 a_100_n76326# a_n100_n76423# a_n158_n76326# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X219 a_100_n200218# a_n100_n200315# a_n158_n200218# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X220 a_100_184638# a_n100_184541# a_n158_184638# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X221 a_100_n247666# a_n100_n247763# a_n158_n247666# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X222 a_100_142462# a_n100_142365# a_n158_142462# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X223 a_100_n5154# a_n100_n5251# a_n158_n5154# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X224 a_100_n208126# a_n100_n208223# a_n158_n208126# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X225 a_100_276898# a_n100_276801# a_n158_276898# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X226 a_100_95014# a_n100_94917# a_n158_95014# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X227 a_100_26478# a_n100_26381# a_n158_26478# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X228 a_100_n252938# a_n100_n253035# a_n158_n252938# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X229 a_100_n210762# a_n100_n210859# a_n158_n210762# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X230 a_100_237358# a_n100_237261# a_n158_237358# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X231 a_100_n89506# a_n100_n89603# a_n158_n89506# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X232 a_100_197818# a_n100_197721# a_n158_197818# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X233 a_100_n292478# a_n100_n292575# a_n158_n292478# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X234 a_100_n139590# a_n100_n139687# a_n158_n139590# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X235 a_100_155642# a_n100_155545# a_n158_155642# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X236 a_100_n305658# a_n100_n305755# a_n158_n305658# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X237 a_100_39658# a_n100_39561# a_n158_39658# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X238 a_100_200454# a_n100_200357# a_n158_200454# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X239 a_100_116102# a_n100_116005# a_n158_116102# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X240 a_100_n52602# a_n100_n52699# a_n158_n52602# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X241 a_100_321710# a_n100_321613# a_n158_321710# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X242 a_100_195182# a_n100_195085# a_n158_195182# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X243 a_100_160914# a_n100_160817# a_n158_160914# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X244 a_100_n171222# a_n100_n171319# a_n158_n171222# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X245 a_100_n102686# a_n100_n102783# a_n158_n102686# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X246 a_100_2754# a_n100_2657# a_n158_2754# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X247 a_100_n310930# a_n100_n311027# a_n158_n310930# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X248 a_100_n223942# a_n100_n224039# a_n158_n223942# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X249 a_100_79198# a_n100_79101# a_n158_79198# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X250 a_100_n92142# a_n100_n92239# a_n158_n92142# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X251 a_100_208362# a_n100_208265# a_n158_208362# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X252 a_100_168822# a_n100_168725# a_n158_168822# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X253 a_100_n266118# a_n100_n266215# a_n158_n266118# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X254 a_100_n263482# a_n100_n263579# a_n158_n263482# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
X255 a_100_n318838# a_n100_n318935# a_n158_n318838# w_n358_n337587# sky130_fd_pr__pfet_g5v0d10v5 ad=3.48 pd=24.58 as=3.48 ps=24.58 w=12 l=1
C0 a_100_n281934# a_n100_n282031# 0.26189f
C1 a_100_303258# a_100_305894# 0.010536f
C2 a_n158_274262# w_n358_n337587# 0.689103f
C3 a_n100_189813# a_n100_192449# 0.205388f
C4 a_n158_150370# w_n358_n337587# 0.689103f
C5 a_n158_n36786# a_n158_n39422# 0.010536f
C6 a_100_121374# a_n158_121374# 0.655843f
C7 a_n100_255713# a_100_255810# 0.26189f
C8 a_n100_n179227# w_n358_n337587# 0.269531f
C9 a_n158_258446# a_n158_261082# 0.010536f
C10 a_n158_n213398# a_n100_n213495# 0.26189f
C11 a_100_89742# a_100_87106# 0.010536f
C12 a_100_n152770# a_100_n155406# 0.010536f
C13 a_n158_216270# a_n158_213634# 0.010536f
C14 a_100_n263482# w_n358_n337587# 0.689103f
C15 a_100_n26242# a_100_n23606# 0.010536f
C16 a_n158_n13062# a_n158_n15698# 0.010536f
C17 a_n100_n289939# a_n100_n292575# 0.205388f
C18 a_n158_284806# a_100_284806# 0.655843f
C19 a_n100_237261# w_n358_n337587# 0.269531f
C20 a_n158_n44694# w_n358_n337587# 0.689103f
C21 a_n158_121374# w_n358_n337587# 0.689103f
C22 a_100_n163314# a_100_n160678# 0.010536f
C23 a_n158_245266# a_100_245266# 0.655843f
C24 a_n100_n266215# a_n100_n268851# 0.205388f
C25 a_100_n123774# a_n100_n123871# 0.26189f
C26 a_100_n250302# a_n158_n250302# 0.655843f
C27 a_n158_5390# a_n158_8026# 0.010536f
C28 a_100_311166# a_100_313802# 0.010536f
C29 a_n100_n155503# a_100_n155406# 0.26189f
C30 a_n158_n229214# a_100_n229214# 0.655843f
C31 a_n100_5293# a_n100_2657# 0.205388f
C32 a_100_200454# w_n358_n337587# 0.689103f
C33 a_n100_34289# a_n158_34386# 0.26189f
C34 a_n158_266354# a_n158_268990# 0.010536f
C35 a_n100_n166047# a_n100_n168683# 0.205388f
C36 a_100_n321474# a_100_n324110# 0.010536f
C37 a_n100_n324207# a_n158_n324110# 0.26189f
C38 a_100_n184402# a_n100_n184499# 0.26189f
C39 a_n100_n42155# a_n100_n39519# 0.205388f
C40 a_n100_n50063# a_n158_n49966# 0.26189f
C41 a_100_295350# a_100_297986# 0.010536f
C42 a_n158_258446# w_n358_n337587# 0.689103f
C43 w_n358_n337587# a_n158_n313566# 0.689103f
C44 a_n158_187274# a_100_187274# 0.655843f
C45 a_n100_187177# a_n100_184541# 0.205388f
C46 a_n158_189910# a_n100_189813# 0.26189f
C47 a_n158_n129046# a_n158_n131682# 0.010536f
C48 a_n158_n31514# a_100_n31514# 0.655843f
C49 a_100_147734# w_n358_n337587# 0.689103f
C50 a_100_118# a_n100_21# 0.26189f
C51 a_n100_303161# w_n358_n337587# 0.269531f
C52 a_n100_318977# a_n158_319074# 0.26189f
C53 a_n100_23745# a_n158_23842# 0.26189f
C54 a_n158_n147498# a_100_n147498# 0.655843f
C55 a_100_n26242# w_n358_n337587# 0.689103f
C56 a_100_158278# w_n358_n337587# 0.689103f
C57 a_n158_n268754# a_100_n268754# 0.655843f
C58 a_n158_n279298# w_n358_n337587# 0.689103f
C59 a_n100_276801# a_100_276898# 0.26189f
C60 a_n158_221542# w_n358_n337587# 0.689103f
C61 a_n158_279534# a_n158_282170# 0.010536f
C62 a_n158_n181766# a_n100_n181863# 0.26189f
C63 a_100_n123774# a_n158_n123774# 0.655843f
C64 a_100_n247666# a_n158_n247666# 0.655843f
C65 a_100_n218670# a_100_n216034# 0.010536f
C66 a_100_239994# a_100_237358# 0.010536f
C67 a_n158_308530# a_n158_305894# 0.010536f
C68 a_n100_192449# a_n158_192546# 0.26189f
C69 a_n100_65921# a_100_66018# 0.26189f
C70 a_n100_279437# w_n358_n337587# 0.269531f
C71 a_n100_n253035# a_n100_n255671# 0.205388f
C72 a_n158_n2518# a_n158_118# 0.010536f
C73 a_100_n284570# a_100_n281934# 0.010536f
C74 a_n100_n289939# a_n158_n289842# 0.26189f
C75 a_n100_n144959# a_n158_n144862# 0.26189f
C76 w_n358_n337587# a_100_n321474# 0.689103f
C77 a_n100_n263579# w_n358_n337587# 0.269531f
C78 a_100_n250302# a_100_n252938# 0.010536f
C79 a_n158_n308294# a_100_n308294# 0.655843f
C80 a_n100_n308391# a_n100_n311027# 0.205388f
C81 a_n100_n10523# w_n358_n337587# 0.269531f
C82 a_n100_326885# w_n358_n337587# 0.269531f
C83 a_100_218906# a_n100_218809# 0.26189f
C84 a_n158_n200218# a_n158_n197582# 0.010536f
C85 a_n100_n152867# a_n100_n150231# 0.205388f
C86 a_n158_55474# a_100_55474# 0.655843f
C87 a_100_13298# a_n100_13201# 0.26189f
C88 a_100_245266# w_n358_n337587# 0.689103f
C89 a_100_n218670# w_n358_n337587# 0.689103f
C90 a_n100_110733# a_n100_113369# 0.205388f
C91 a_n100_245169# a_n100_247805# 0.205388f
C92 a_n100_n258307# w_n358_n337587# 0.269531f
C93 a_n158_n176494# w_n358_n337587# 0.689103f
C94 a_n158_n126410# a_n158_n123774# 0.010536f
C95 a_n100_n292575# a_n100_n295211# 0.205388f
C96 a_n158_n179130# a_100_n179130# 0.655843f
C97 a_100_168822# a_100_166186# 0.010536f
C98 a_n100_166089# a_n158_166186# 0.26189f
C99 a_n158_n165950# a_n158_n168586# 0.010536f
C100 a_n158_23842# w_n358_n337587# 0.689103f
C101 a_100_113466# w_n358_n337587# 0.689103f
C102 a_n100_n253035# a_n158_n252938# 0.26189f
C103 a_n158_n76326# w_n358_n337587# 0.689103f
C104 a_n158_n60510# a_100_n60510# 0.655843f
C105 a_n158_n202854# a_100_n202854# 0.655843f
C106 a_n158_189910# a_n158_192546# 0.010536f
C107 a_n100_60649# a_n100_63285# 0.205388f
C108 a_n100_n123871# w_n358_n337587# 0.269531f
C109 a_n100_n297847# a_100_n297750# 0.26189f
C110 a_n100_n313663# a_100_n313566# 0.26189f
C111 a_n100_n76423# a_n100_n79059# 0.205388f
C112 a_100_n39422# a_100_n42058# 0.010536f
C113 a_n158_179366# w_n358_n337587# 0.689103f
C114 a_n100_258349# a_100_258446# 0.26189f
C115 a_n158_n31514# w_n358_n337587# 0.689103f
C116 a_n100_n226675# a_n100_n224039# 0.205388f
C117 a_100_n44694# a_n100_n44791# 0.26189f
C118 a_100_n263482# a_n100_n263579# 0.26189f
C119 a_n158_311166# w_n358_n337587# 0.689103f
C120 a_n100_89645# a_100_89742# 0.26189f
C121 a_100_142462# a_100_145098# 0.010536f
C122 a_n100_42197# a_n100_44833# 0.205388f
C123 a_100_50202# a_100_47566# 0.010536f
C124 a_n158_n15698# w_n358_n337587# 0.689103f
C125 a_n100_287345# a_100_287442# 0.26189f
C126 a_n100_105461# a_n100_108097# 0.205388f
C127 a_n100_110733# a_100_110830# 0.26189f
C128 a_n158_126646# w_n358_n337587# 0.689103f
C129 a_n158_234722# a_100_234722# 0.655843f
C130 a_100_239994# a_100_242630# 0.010536f
C131 a_100_n250302# w_n358_n337587# 0.689103f
C132 a_n158_n2518# a_n158_n5154# 0.010536f
C133 a_100_29114# a_n100_29017# 0.26189f
C134 a_n100_308433# a_n100_311069# 0.205388f
C135 a_100_287442# w_n358_n337587# 0.689103f
C136 a_n100_10565# a_n100_7929# 0.205388f
C137 a_n100_n247763# a_n100_n245127# 0.205388f
C138 a_n100_131821# a_n158_131918# 0.26189f
C139 a_n158_203090# w_n358_n337587# 0.689103f
C140 a_100_97650# a_100_100286# 0.010536f
C141 w_n358_n337587# a_n158_334890# 0.693647f
C142 a_n158_n123774# w_n358_n337587# 0.689103f
C143 a_n100_152909# a_n100_150273# 0.205388f
C144 a_n158_n258210# a_n158_n260846# 0.010536f
C145 a_n158_295350# a_n100_295253# 0.26189f
C146 a_100_n107958# a_100_n105322# 0.010536f
C147 a_100_n65782# w_n358_n337587# 0.689103f
C148 a_n158_52838# a_100_52838# 0.655843f
C149 a_n158_182002# a_n158_184638# 0.010536f
C150 a_n158_250538# w_n358_n337587# 0.689103f
C151 a_n100_n55335# a_100_n55238# 0.26189f
C152 a_n158_118738# a_100_118738# 0.655843f
C153 a_n158_n2518# a_100_n2518# 0.655843f
C154 a_100_247902# a_n158_247902# 0.655843f
C155 a_n100_250441# a_100_250538# 0.26189f
C156 a_n100_168725# w_n358_n337587# 0.269531f
C157 a_n100_316341# a_n100_318977# 0.205388f
C158 a_100_324346# a_100_321710# 0.010536f
C159 a_100_84470# a_n100_84373# 0.26189f
C160 a_100_n329382# a_100_n332018# 0.010536f
C161 a_n100_n332115# a_n158_n332018# 0.26189f
C162 a_100_n129046# w_n358_n337587# 0.689103f
C163 w_n358_n337587# a_n158_n303022# 0.689103f
C164 a_n158_n36786# w_n358_n337587# 0.689103f
C165 a_n100_39561# a_n158_39658# 0.26189f
C166 a_n158_213634# w_n358_n337587# 0.689103f
C167 a_n100_21# w_n358_n337587# 0.269531f
C168 a_n158_n171222# w_n358_n337587# 0.689103f
C169 a_n158_105558# a_n100_105461# 0.26189f
C170 a_100_34386# w_n358_n337587# 0.689103f
C171 a_n100_184541# w_n358_n337587# 0.269531f
C172 a_100_126646# a_100_124010# 0.010536f
C173 a_n100_123913# a_n158_124010# 0.26189f
C174 a_n158_21206# a_100_21206# 0.655843f
C175 a_n158_n229214# w_n358_n337587# 0.689103f
C176 a_n158_n231850# w_n358_n337587# 0.689103f
C177 w_n358_n337587# a_n158_n310930# 0.689103f
C178 a_n158_329618# a_n158_326982# 0.010536f
C179 a_n158_n107958# a_n158_n105322# 0.010536f
C180 a_n158_87106# a_100_87106# 0.655843f
C181 a_100_92378# a_100_95014# 0.010536f
C182 a_100_216270# a_100_213634# 0.010536f
C183 a_n100_213537# a_n158_213634# 0.26189f
C184 a_n158_n63146# w_n358_n337587# 0.689103f
C185 a_n158_n52602# a_n158_n55238# 0.010536f
C186 a_100_n107958# a_100_n110594# 0.010536f
C187 a_n100_158181# a_n100_155545# 0.205388f
C188 a_n158_245266# a_n158_242630# 0.010536f
C189 a_n158_239994# a_n100_239897# 0.26189f
C190 a_100_n20970# a_100_n23606# 0.010536f
C191 a_100_n110594# a_100_n113230# 0.010536f
C192 a_n100_52741# w_n358_n337587# 0.269531f
C193 a_100_311166# a_n100_311069# 0.26189f
C194 a_n158_n192310# w_n358_n337587# 0.689103f
C195 a_n158_131918# a_n158_134554# 0.010536f
C196 a_n100_n50063# w_n358_n337587# 0.269531f
C197 a_n100_15837# w_n358_n337587# 0.269531f
C198 a_n100_n274123# a_100_n274026# 0.26189f
C199 a_n100_197721# w_n358_n337587# 0.269531f
C200 a_n158_n284570# a_100_n284570# 0.655843f
C201 w_n358_n337587# a_100_n318838# 0.689103f
C202 a_n100_n218767# a_n100_n216131# 0.205388f
C203 a_n100_n181863# w_n358_n337587# 0.269531f
C204 a_100_n18334# a_100_n20970# 0.010536f
C205 a_100_258446# w_n358_n337587# 0.689103f
C206 w_n358_n337587# a_n100_n337387# 0.349164f
C207 a_n158_145098# w_n358_n337587# 0.689103f
C208 a_n158_n78962# w_n358_n337587# 0.689103f
C209 a_n100_n34247# w_n358_n337587# 0.269531f
C210 a_100_n205490# a_100_n202854# 0.010536f
C211 a_n100_n36883# a_100_n36786# 0.26189f
C212 a_n100_73829# w_n358_n337587# 0.269531f
C213 a_n158_15934# a_n158_13298# 0.010536f
C214 a_n100_n47427# a_n100_n50063# 0.205388f
C215 a_n100_139729# a_n100_142365# 0.205388f
C216 a_n158_n84234# a_n158_n81598# 0.010536f
C217 a_n158_174094# a_100_174094# 0.655843f
C218 a_n100_n268851# w_n358_n337587# 0.269531f
C219 a_100_n10426# a_100_n13062# 0.010536f
C220 a_n100_n158139# a_n100_n160775# 0.205388f
C221 a_n100_n147595# a_100_n147498# 0.26189f
C222 a_n158_279534# w_n358_n337587# 0.689103f
C223 a_100_n7790# a_100_n5154# 0.010536f
C224 a_n158_192546# a_100_192546# 0.655843f
C225 a_100_39658# w_n358_n337587# 0.689103f
C226 a_n158_n205490# a_n158_n208126# 0.010536f
C227 a_100_n20970# w_n358_n337587# 0.689103f
C228 a_n158_66018# a_100_66018# 0.655843f
C229 a_n158_n245030# w_n358_n337587# 0.689103f
C230 a_100_n208126# a_n158_n208126# 0.655843f
C231 a_n158_n210762# a_100_n210762# 0.655843f
C232 a_n100_n181863# a_n100_n179227# 0.205388f
C233 a_n100_n23703# a_100_n23606# 0.26189f
C234 a_n100_224081# a_n158_224178# 0.26189f
C235 a_n158_n295114# a_n158_n297750# 0.010536f
C236 a_n158_n310930# a_n158_n313566# 0.010536f
C237 a_n158_326982# w_n358_n337587# 0.689103f
C238 a_n100_97553# a_n158_97650# 0.26189f
C239 a_n100_216173# a_n100_218809# 0.205388f
C240 a_100_n76326# a_n100_n76423# 0.26189f
C241 a_100_n234486# a_n158_n234486# 0.655843f
C242 a_n100_n221403# a_n158_n221306# 0.26189f
C243 a_100_13298# a_n158_13298# 0.655843f
C244 a_n100_10565# a_n100_13201# 0.205388f
C245 a_n158_242630# w_n358_n337587# 0.689103f
C246 a_100_n5154# a_n100_n5251# 0.26189f
C247 a_n100_n202951# a_100_n202854# 0.26189f
C248 a_n100_129185# w_n358_n337587# 0.269531f
C249 a_n158_84470# a_100_84470# 0.655843f
C250 a_n100_300525# w_n358_n337587# 0.269531f
C251 a_n100_n113327# a_100_n113230# 0.26189f
C252 a_n158_271626# a_n158_268990# 0.010536f
C253 a_n100_n89603# a_n158_n89506# 0.26189f
C254 a_n100_n150231# w_n358_n337587# 0.269531f
C255 a_n158_166186# a_100_166186# 0.655843f
C256 a_n100_34289# a_n100_36925# 0.205388f
C257 a_n158_n266118# a_100_n266118# 0.655843f
C258 a_100_n234486# a_n100_n234583# 0.26189f
C259 a_100_100286# a_n100_100189# 0.26189f
C260 a_100_226814# a_n100_226717# 0.26189f
C261 a_n100_229353# a_n158_229450# 0.26189f
C262 a_n100_155545# w_n358_n337587# 0.269531f
C263 a_n158_266354# w_n358_n337587# 0.689103f
C264 a_n100_n316299# a_n100_n318935# 0.205388f
C265 a_n100_58013# a_n158_58110# 0.26189f
C266 a_n158_n57874# a_100_n57874# 0.655843f
C267 a_n100_152909# w_n358_n337587# 0.269531f
C268 a_n100_n123871# a_n158_n123774# 0.26189f
C269 a_n100_n247763# a_n158_n247666# 0.26189f
C270 a_100_n187038# a_100_n189674# 0.010536f
C271 a_n158_n292478# w_n358_n337587# 0.689103f
C272 a_n100_n71151# w_n358_n337587# 0.269531f
C273 a_100_179366# w_n358_n337587# 0.689103f
C274 a_n158_258446# a_100_258446# 0.655843f
C275 a_100_n287206# w_n358_n337587# 0.689103f
C276 a_n158_89742# a_100_89742# 0.655843f
C277 a_100_324346# w_n358_n337587# 0.689103f
C278 a_n100_n23703# w_n358_n337587# 0.269531f
C279 a_100_n28878# a_n100_n28975# 0.26189f
C280 a_100_142462# a_n100_142365# 0.26189f
C281 a_n100_47469# a_100_47566# 0.26189f
C282 a_n158_n150134# w_n358_n337587# 0.689103f
C283 a_n100_n63243# a_100_n63146# 0.26189f
C284 a_n100_110733# a_n100_108097# 0.205388f
C285 a_n100_n210859# a_100_n210762# 0.26189f
C286 a_n100_n266215# a_100_n266118# 0.26189f
C287 a_n158_71290# a_n100_71193# 0.26189f
C288 a_100_47566# w_n358_n337587# 0.689103f
C289 a_100_n5154# w_n358_n337587# 0.689103f
C290 a_n100_202993# a_100_203090# 0.26189f
C291 a_100_266354# a_100_268990# 0.010536f
C292 a_100_18570# a_100_21206# 0.010536f
C293 a_100_n194946# a_n158_n194946# 0.655843f
C294 a_n100_263621# a_n158_263718# 0.26189f
C295 a_100_n318838# a_100_n321474# 0.010536f
C296 a_n100_n321571# a_n158_n321474# 0.26189f
C297 a_n100_n81695# a_100_n81598# 0.26189f
C298 w_n358_n337587# a_n100_332157# 0.269531f
C299 a_n100_334793# a_100_334890# 0.26189f
C300 a_n100_160817# a_n158_160914# 0.26189f
C301 a_100_224178# a_100_221542# 0.010536f
C302 a_n158_n271390# w_n358_n337587# 0.689103f
C303 a_n100_n110691# a_n100_n108055# 0.205388f
C304 a_100_295350# a_n100_295253# 0.26189f
C305 a_n100_247805# w_n358_n337587# 0.269531f
C306 a_n100_n39519# a_100_n39422# 0.26189f
C307 w_n358_n337587# a_n100_n300483# 0.269531f
C308 a_n158_n81598# w_n358_n337587# 0.689103f
C309 a_n158_n155406# a_n158_n158042# 0.010536f
C310 a_n158_n221306# w_n358_n337587# 0.689103f
C311 a_n100_321613# a_n100_318977# 0.205388f
C312 a_n158_n168586# a_100_n168586# 0.655843f
C313 a_100_205726# a_n100_205629# 0.26189f
C314 a_n100_81737# a_n100_84373# 0.205388f
C315 a_n158_81834# a_n158_79198# 0.010536f
C316 a_n100_208265# a_100_208362# 0.26189f
C317 a_n158_n337290# a_100_n337290# 0.655843f
C318 a_n100_n60607# a_n158_n60510# 0.26189f
C319 a_n100_n158139# a_100_n158042# 0.26189f
C320 a_n100_21109# a_n100_23745# 0.205388f
C321 a_100_n57874# w_n358_n337587# 0.689103f
C322 a_n100_n208223# w_n358_n337587# 0.269531f
C323 a_n100_39561# a_n100_36925# 0.205388f
C324 a_100_n255574# a_n100_n255671# 0.26189f
C325 a_100_282170# a_100_279534# 0.010536f
C326 a_n100_279437# a_n158_279534# 0.26189f
C327 a_100_n89506# a_n158_n89506# 0.655843f
C328 a_n100_102825# a_n100_100189# 0.205388f
C329 a_100_105558# a_n100_105461# 0.26189f
C330 a_n100_300525# a_n100_303161# 0.205388f
C331 a_n100_n94875# a_100_n94778# 0.26189f
C332 a_n158_n20970# w_n358_n337587# 0.689103f
C333 a_n100_68557# a_n158_68654# 0.26189f
C334 a_n100_31653# w_n358_n337587# 0.269531f
C335 a_n100_195085# a_n100_192449# 0.205388f
C336 a_n158_n305658# a_100_n305658# 0.655843f
C337 a_n100_n113327# a_n158_n113230# 0.26189f
C338 a_100_n279298# a_100_n281934# 0.010536f
C339 a_n100_123913# a_100_124010# 0.26189f
C340 a_n158_5390# w_n358_n337587# 0.689103f
C341 a_n100_326885# a_n158_326982# 0.26189f
C342 a_100_92378# a_n100_92281# 0.26189f
C343 a_n100_n303119# a_100_n303022# 0.26189f
C344 a_n158_n76326# a_n158_n78962# 0.010536f
C345 a_100_n274026# a_n158_n274026# 0.655843f
C346 w_n358_n337587# a_n100_n334751# 0.269531f
C347 a_100_n44694# a_100_n42058# 0.010536f
C348 a_100_237358# w_n358_n337587# 0.689103f
C349 a_n158_n129046# a_n100_n129143# 0.26189f
C350 a_100_134554# w_n358_n337587# 0.689103f
C351 a_n100_292617# w_n358_n337587# 0.269531f
C352 a_n100_n26339# a_n158_n26242# 0.26189f
C353 a_n158_n255574# a_100_n255574# 0.655843f
C354 a_100_155642# a_n158_155642# 0.655843f
C355 a_n158_29114# a_n100_29017# 0.26189f
C356 a_n100_21109# w_n358_n337587# 0.269531f
C357 a_n100_n86967# a_n100_n89603# 0.205388f
C358 a_n158_210998# w_n358_n337587# 0.689103f
C359 a_n100_n171319# a_n100_n168683# 0.205388f
C360 a_100_58110# a_100_60746# 0.010536f
C361 a_n158_187274# a_n158_184638# 0.010536f
C362 a_100_189910# a_n100_189813# 0.26189f
C363 a_n158_n160678# a_n100_n160775# 0.26189f
C364 a_100_145098# w_n358_n337587# 0.689103f
C365 a_n158_n23606# a_100_n23606# 0.655843f
C366 a_n158_176730# w_n358_n337587# 0.689103f
C367 a_n158_n229214# a_n158_n231850# 0.010536f
C368 a_n100_n287303# w_n358_n337587# 0.269531f
C369 a_100_n200218# a_100_n197582# 0.010536f
C370 a_n158_n68418# a_100_n68418# 0.655843f
C371 a_n100_n55335# a_n158_n55238# 0.26189f
C372 a_n100_318977# a_100_319074# 0.26189f
C373 a_n100_205629# a_n158_205726# 0.26189f
C374 a_100_221542# w_n358_n337587# 0.689103f
C375 a_n100_n239855# a_n100_n237219# 0.205388f
C376 a_n158_n239758# w_n358_n337587# 0.689103f
C377 a_n100_116005# w_n358_n337587# 0.269531f
C378 a_n100_n86967# a_n100_n84331# 0.205388f
C379 a_n100_237261# a_100_237358# 0.26189f
C380 a_100_308530# a_100_305894# 0.010536f
C381 a_n100_305797# a_n158_305894# 0.26189f
C382 a_n100_n147595# a_n100_n144959# 0.205388f
C383 a_n158_n295114# a_100_n295114# 0.655843f
C384 a_n100_n295211# a_n100_n297847# 0.205388f
C385 a_n100_n274123# w_n358_n337587# 0.269531f
C386 a_n158_n71054# w_n358_n337587# 0.689103f
C387 a_100_326982# w_n358_n337587# 0.689103f
C388 a_100_n239758# a_n158_n239758# 0.655843f
C389 a_n100_97553# a_100_97650# 0.26189f
C390 a_n100_224081# a_100_224178# 0.26189f
C391 a_n158_n89506# w_n358_n337587# 0.689103f
C392 a_100_n7790# a_100_n10426# 0.010536f
C393 a_n158_n121138# a_100_n121138# 0.655843f
C394 a_100_242630# w_n358_n337587# 0.689103f
C395 a_n100_n76423# w_n358_n337587# 0.269531f
C396 a_n158_295350# a_100_295350# 0.655843f
C397 a_100_182002# a_100_184638# 0.010536f
C398 a_n158_179366# a_100_179366# 0.655843f
C399 a_100_129282# w_n358_n337587# 0.689103f
C400 a_100_n187038# a_n100_n187135# 0.26189f
C401 a_n158_n197582# w_n358_n337587# 0.689103f
C402 a_n158_n163314# a_100_n163314# 0.655843f
C403 a_n158_n23606# w_n358_n337587# 0.689103f
C404 a_n158_n226578# a_100_n226578# 0.655843f
C405 a_n158_n97414# a_n158_n94778# 0.010536f
C406 a_n100_n192407# w_n358_n337587# 0.269531f
C407 a_100_n102686# a_100_n105322# 0.010536f
C408 a_100_n326746# a_100_n329382# 0.010536f
C409 a_n100_n329479# a_n158_n329382# 0.26189f
C410 a_100_n123774# a_100_n126410# 0.010536f
C411 a_n100_n142323# a_n158_n142226# 0.26189f
C412 a_n100_210901# w_n358_n337587# 0.269531f
C413 a_n100_n60607# a_n100_n63243# 0.205388f
C414 a_n100_n68515# a_100_n68418# 0.26189f
C415 a_n100_n226675# a_100_n226578# 0.26189f
C416 a_n158_n92142# a_n158_n94778# 0.010536f
C417 a_n100_n197679# a_100_n197582# 0.26189f
C418 a_n158_n194946# w_n358_n337587# 0.689103f
C419 a_n100_166089# a_n100_163453# 0.205388f
C420 a_n100_n176591# w_n358_n337587# 0.269531f
C421 a_n158_105558# a_100_105558# 0.655843f
C422 a_100_226814# a_n158_226814# 0.655843f
C423 a_100_300622# a_100_297986# 0.010536f
C424 a_n100_297889# a_n158_297986# 0.26189f
C425 w_n358_n337587# a_n158_n308294# 0.689103f
C426 a_n100_176633# w_n358_n337587# 0.269531f
C427 a_n158_n326746# a_n158_n329382# 0.010536f
C428 a_n100_n234583# a_n100_n237219# 0.205388f
C429 a_n158_81834# w_n358_n337587# 0.689103f
C430 a_n158_89742# a_n158_87106# 0.010536f
C431 a_n100_210901# a_n100_213537# 0.205388f
C432 a_100_147734# a_100_145098# 0.010536f
C433 a_n100_n18431# a_n158_n18334# 0.26189f
C434 a_100_142462# a_n158_142462# 0.655843f
C435 a_100_229450# w_n358_n337587# 0.689103f
C436 a_n158_n258210# w_n358_n337587# 0.689103f
C437 a_n158_n126410# a_100_n126410# 0.655843f
C438 a_100_n78962# a_100_n81598# 0.010536f
C439 a_n100_n131779# a_n158_n131682# 0.26189f
C440 a_n100_n42155# w_n358_n337587# 0.269531f
C441 a_100_n292478# a_n100_n292575# 0.26189f
C442 a_n158_118# a_n158_2754# 0.010536f
C443 a_n100_n176591# a_n100_n179227# 0.205388f
C444 a_100_18570# a_n100_18473# 0.26189f
C445 a_n158_n216034# a_100_n216034# 0.655843f
C446 a_n158_263718# a_100_263718# 0.655843f
C447 a_n158_n26242# a_n158_n28878# 0.010536f
C448 a_n158_155642# a_n158_158278# 0.010536f
C449 a_n158_160914# a_100_160914# 0.655843f
C450 a_n100_n160775# w_n358_n337587# 0.269531f
C451 a_n158_221542# a_100_221542# 0.655843f
C452 a_n158_n242394# a_100_n242394# 0.655843f
C453 a_n100_55377# a_n100_58013# 0.205388f
C454 a_100_n10426# w_n358_n337587# 0.689103f
C455 w_n358_n337587# a_n100_n332115# 0.269531f
C456 a_100_n181766# a_100_n184402# 0.010536f
C457 a_n158_253174# a_n100_253077# 0.26189f
C458 a_100_n202854# w_n358_n337587# 0.689103f
C459 a_n158_208362# a_100_208362# 0.655843f
C460 a_n100_65921# w_n358_n337587# 0.269531f
C461 a_100_n97414# a_100_n94778# 0.010536f
C462 a_n158_n216034# w_n358_n337587# 0.689103f
C463 a_n100_26381# a_100_26478# 0.26189f
C464 a_n100_224081# w_n358_n337587# 0.269531f
C465 a_100_n266118# w_n358_n337587# 0.689103f
C466 a_n158_n129046# a_n158_n126410# 0.010536f
C467 a_n100_n224039# a_n100_n221403# 0.205388f
C468 a_n158_108194# w_n358_n337587# 0.689103f
C469 a_n158_102922# a_100_102922# 0.655843f
C470 a_n158_10662# a_n158_13298# 0.010536f
C471 a_n100_7929# a_n158_8026# 0.26189f
C472 a_n100_102825# a_n100_105461# 0.205388f
C473 a_100_n94778# w_n358_n337587# 0.689103f
C474 a_n158_271626# w_n358_n337587# 0.689103f
C475 a_n100_68557# a_100_68654# 0.26189f
C476 a_n100_308433# a_n158_308530# 0.26189f
C477 a_100_197818# a_n158_197818# 0.655843f
C478 a_n100_123913# a_n100_121277# 0.205388f
C479 a_100_n126410# w_n358_n337587# 0.689103f
C480 a_n158_21206# a_n158_18570# 0.010536f
C481 a_100_n310930# a_n100_n311027# 0.26189f
C482 a_n100_326885# a_100_326982# 0.26189f
C483 a_100_n223942# w_n358_n337587# 0.689103f
C484 a_n100_n86967# w_n358_n337587# 0.269531f
C485 a_n100_234625# w_n358_n337587# 0.269531f
C486 a_100_n92142# a_n100_n92239# 0.26189f
C487 a_n100_n171319# a_100_n171222# 0.26189f
C488 a_n100_n189771# a_n158_n189674# 0.26189f
C489 a_n158_176730# a_n158_179366# 0.010536f
C490 a_100_110830# a_100_108194# 0.010536f
C491 a_n100_131821# w_n358_n337587# 0.269531f
C492 a_100_245266# a_100_242630# 0.010536f
C493 a_n100_n284667# w_n358_n337587# 0.269531f
C494 a_n100_313705# a_n158_313802# 0.26189f
C495 a_n158_52838# w_n358_n337587# 0.689103f
C496 a_n100_n205587# a_n158_n205490# 0.26189f
C497 a_100_n258210# a_100_n260846# 0.010536f
C498 a_n158_n102686# a_n158_n105322# 0.010536f
C499 a_n158_34386# a_n158_31750# 0.010536f
C500 a_100_210998# w_n358_n337587# 0.689103f
C501 a_n158_274262# a_n158_271626# 0.010536f
C502 a_n158_n2518# w_n358_n337587# 0.689103f
C503 a_n100_n129143# a_n100_n126507# 0.205388f
C504 a_100_n263482# a_100_n266118# 0.010536f
C505 a_n100_n86967# a_100_n86870# 0.26189f
C506 a_n158_n250302# a_n158_n252938# 0.010536f
C507 a_n158_n42058# a_100_n42058# 0.655843f
C508 a_n158_n57874# a_n158_n60510# 0.010536f
C509 a_n100_97553# a_n100_100189# 0.205388f
C510 a_100_58110# a_n100_58013# 0.26189f
C511 a_100_63382# a_100_60746# 0.010536f
C512 a_n100_60649# a_n158_60746# 0.26189f
C513 a_n100_n176591# a_n158_n176494# 0.26189f
C514 a_n100_n200315# a_100_n200218# 0.26189f
C515 a_n100_n76423# a_n158_n76326# 0.26189f
C516 a_n158_n165950# a_100_n165950# 0.655843f
C517 a_100_5390# w_n358_n337587# 0.689103f
C518 a_n100_181905# w_n358_n337587# 0.269531f
C519 a_n100_142365# w_n358_n337587# 0.269531f
C520 a_100_n144862# a_n158_n144862# 0.655843f
C521 a_n158_n274026# w_n358_n337587# 0.689103f
C522 a_n158_n129046# w_n358_n337587# 0.689103f
C523 a_n100_n271487# a_100_n271390# 0.26189f
C524 a_100_73926# w_n358_n337587# 0.689103f
C525 a_100_84470# a_100_87106# 0.010536f
C526 a_100_316438# w_n358_n337587# 0.689103f
C527 a_n158_319074# a_100_319074# 0.655843f
C528 a_n158_210998# a_n158_213634# 0.010536f
C529 a_n100_n31611# a_n100_n28975# 0.205388f
C530 a_n158_n81598# a_n158_n78962# 0.010536f
C531 a_n100_n105419# w_n358_n337587# 0.269531f
C532 a_100_42294# a_100_44930# 0.010536f
C533 a_n158_116102# w_n358_n337587# 0.689103f
C534 a_n100_237261# a_n100_234625# 0.205388f
C535 a_n158_26478# a_n158_29114# 0.010536f
C536 a_100_26478# a_100_23842# 0.010536f
C537 a_100_239994# a_n158_239994# 0.655843f
C538 a_n158_276898# w_n358_n337587# 0.689103f
C539 a_n158_37022# w_n358_n337587# 0.689103f
C540 a_n100_305797# a_100_305894# 0.26189f
C541 a_100_71290# a_100_73926# 0.010536f
C542 a_n100_n224039# w_n358_n337587# 0.269531f
C543 a_100_n158042# w_n358_n337587# 0.689103f
C544 a_n100_n258307# a_n158_n258210# 0.26189f
C545 a_n100_n318935# a_n158_n318838# 0.26189f
C546 a_n100_192449# w_n358_n337587# 0.269531f
C547 a_n100_266257# a_100_266354# 0.26189f
C548 a_100_332254# w_n358_n337587# 0.689103f
C549 w_n358_n337587# a_n158_n305658# 0.689103f
C550 a_n100_152909# a_n100_155545# 0.205388f
C551 a_100_n10426# a_n100_n10523# 0.26189f
C552 a_100_n136954# a_n158_n136954# 0.655843f
C553 a_100_n39422# a_n158_n39422# 0.655843f
C554 a_n158_n237122# a_n100_n237219# 0.26189f
C555 a_n100_n163411# a_n158_n163314# 0.26189f
C556 a_100_n252938# a_n158_n252938# 0.655843f
C557 a_100_n184402# a_n158_n184402# 0.655843f
C558 a_100_n110594# a_n158_n110594# 0.655843f
C559 a_100_n260846# a_n100_n260943# 0.26189f
C560 a_n158_n150134# a_n100_n150231# 0.26189f
C561 a_n100_n7887# a_n158_n7790# 0.26189f
C562 a_n100_n326843# a_100_n326746# 0.26189f
C563 a_n158_295350# a_n158_292714# 0.010536f
C564 a_n158_n284570# a_n158_n287206# 0.010536f
C565 a_n158_n60510# w_n358_n337587# 0.689103f
C566 a_n100_166089# w_n358_n337587# 0.269531f
C567 a_100_n237122# a_100_n234486# 0.010536f
C568 a_n158_134554# w_n358_n337587# 0.689103f
C569 a_n158_245266# a_n158_247902# 0.010536f
C570 a_n100_n197679# a_n100_n200315# 0.205388f
C571 a_n158_n334654# a_100_n334654# 0.655843f
C572 a_n100_n334751# a_n100_n337387# 0.205388f
C573 a_n158_n134318# a_n158_n136954# 0.010536f
C574 a_n158_n168586# w_n358_n337587# 0.689103f
C575 a_n158_n281934# a_n100_n282031# 0.26189f
C576 a_100_79198# a_n100_79101# 0.26189f
C577 a_n158_316438# a_n158_319074# 0.010536f
C578 a_n100_n13159# a_n100_n15795# 0.205388f
C579 a_n100_139729# a_n158_139826# 0.26189f
C580 a_100_218906# w_n358_n337587# 0.689103f
C581 a_n158_274262# a_n158_276898# 0.010536f
C582 a_n158_n20970# a_100_n20970# 0.655843f
C583 a_n158_168822# a_100_168822# 0.655843f
C584 a_n158_232086# a_n100_231989# 0.26189f
C585 a_n100_229353# a_n100_226717# 0.205388f
C586 a_n100_n255671# w_n358_n337587# 0.269531f
C587 w_n358_n337587# a_n158_n295114# 0.689103f
C588 a_n158_297986# a_100_297986# 0.655843f
C589 a_n158_63382# a_n158_66018# 0.010536f
C590 a_100_n234486# a_100_n231850# 0.010536f
C591 a_n158_153006# w_n358_n337587# 0.689103f
C592 a_n158_189910# w_n358_n337587# 0.689103f
C593 a_n158_n28878# a_100_n28878# 0.655843f
C594 w_n358_n337587# a_n100_n329479# 0.269531f
C595 a_n100_n55335# a_n100_n57971# 0.205388f
C596 a_100_92378# a_n158_92378# 0.655843f
C597 a_n100_216173# a_n158_216270# 0.26189f
C598 a_n158_145098# a_100_145098# 0.655843f
C599 a_n158_287442# a_n158_284806# 0.010536f
C600 a_100_50202# a_n158_50202# 0.655843f
C601 a_100_n189674# w_n358_n337587# 0.689103f
C602 a_n100_n52699# a_100_n52602# 0.26189f
C603 a_100_n305658# a_n100_n305755# 0.26189f
C604 a_100_n115866# a_100_n113230# 0.010536f
C605 a_n100_n276759# w_n358_n337587# 0.269531f
C606 a_100_n163314# w_n358_n337587# 0.689103f
C607 a_100_284806# w_n358_n337587# 0.689103f
C608 a_100_n300386# a_100_n297750# 0.010536f
C609 a_100_n105322# w_n358_n337587# 0.689103f
C610 a_100_18570# a_n158_18570# 0.655843f
C611 a_n158_131918# a_100_131918# 0.655843f
C612 a_n100_200357# w_n358_n337587# 0.269531f
C613 a_n158_n252938# w_n358_n337587# 0.689103f
C614 a_n158_n255574# w_n358_n337587# 0.689103f
C615 w_n358_n337587# a_n158_n326746# 0.689103f
C616 a_n100_221445# a_n100_218809# 0.205388f
C617 a_n100_289981# a_n158_290078# 0.26189f
C618 a_n158_153006# a_n158_150370# 0.010536f
C619 a_n158_247902# w_n358_n337587# 0.689103f
C620 a_n158_n310930# a_n158_n308294# 0.010536f
C621 a_100_n36786# a_100_n34150# 0.010536f
C622 a_100_184638# a_100_187274# 0.010536f
C623 a_n100_n68515# a_n158_n68418# 0.26189f
C624 a_n100_n108055# a_n158_n107958# 0.26189f
C625 a_n100_n192407# a_n158_n192310# 0.26189f
C626 a_100_253174# a_n100_253077# 0.26189f
C627 a_n158_174094# w_n358_n337587# 0.689103f
C628 a_n158_n192310# a_n158_n194946# 0.010536f
C629 a_n158_66018# w_n358_n337587# 0.689103f
C630 a_n100_208265# a_n100_205629# 0.205388f
C631 a_100_n289842# a_n158_n289842# 0.655843f
C632 a_100_n194946# a_n100_n195043# 0.26189f
C633 a_100_205726# a_n158_205726# 0.655843f
C634 a_100_n139590# a_n158_n139590# 0.655843f
C635 a_n158_26478# a_100_26478# 0.655843f
C636 a_n100_26381# a_n100_23745# 0.205388f
C637 a_n158_137190# a_100_137190# 0.655843f
C638 a_100_n47330# a_100_n49966# 0.010536f
C639 a_n100_n242491# w_n358_n337587# 0.269531f
C640 a_n158_42294# a_n100_42197# 0.26189f
C641 a_100_168822# a_100_171458# 0.010536f
C642 a_n100_n187135# a_n158_n187038# 0.26189f
C643 a_n158_113466# w_n358_n337587# 0.689103f
C644 a_n158_102922# a_n158_100286# 0.010536f
C645 a_100_n115866# a_n158_n115866# 0.655843f
C646 a_n100_n155503# a_n158_n155406# 0.26189f
C647 a_100_n110594# w_n358_n337587# 0.689103f
C648 a_100_271626# w_n358_n337587# 0.689103f
C649 a_n100_308433# a_100_308530# 0.26189f
C650 a_n158_68654# a_100_68654# 0.655843f
C651 a_n158_303258# a_n158_305894# 0.010536f
C652 a_n100_29017# w_n358_n337587# 0.269531f
C653 a_100_n187038# a_100_n184402# 0.010536f
C654 a_100_126646# a_n100_126549# 0.26189f
C655 a_100_261082# a_100_263718# 0.010536f
C656 a_n158_n126410# a_n100_n126507# 0.26189f
C657 a_100_n131682# a_n100_n131779# 0.26189f
C658 a_100_n313566# a_100_n316202# 0.010536f
C659 a_n100_n316299# a_n158_n316202# 0.26189f
C660 a_n158_326982# a_100_326982# 0.655843f
C661 a_n100_89645# a_n100_92281# 0.205388f
C662 a_100_234722# w_n358_n337587# 0.689103f
C663 a_100_50202# a_n100_50105# 0.26189f
C664 a_100_n194946# a_100_n192310# 0.010536f
C665 a_100_n287206# a_n100_n287303# 0.26189f
C666 a_100_n147498# a_100_n150134# 0.010536f
C667 a_n100_108097# a_100_108194# 0.26189f
C668 a_n158_242630# a_100_242630# 0.655843f
C669 a_n100_242533# a_n100_239897# 0.205388f
C670 a_n100_n63243# w_n358_n337587# 0.269531f
C671 a_100_n129046# a_100_n126410# 0.010536f
C672 a_n158_316438# a_n100_316341# 0.26189f
C673 a_n100_n21067# w_n358_n337587# 0.269531f
C674 a_n100_200357# a_100_200454# 0.26189f
C675 a_n100_76465# a_n100_79101# 0.205388f
C676 a_100_203090# a_100_205726# 0.010536f
C677 a_n100_129185# a_100_129282# 0.26189f
C678 a_n100_26381# w_n358_n337587# 0.269531f
C679 a_100_268990# a_n100_268893# 0.26189f
C680 a_n158_102922# w_n358_n337587# 0.689103f
C681 a_n158_97650# a_n158_100286# 0.010536f
C682 a_n158_255810# w_n358_n337587# 0.689103f
C683 a_n100_60649# a_100_60746# 0.26189f
C684 a_100_8026# a_100_10662# 0.010536f
C685 a_100_n276662# a_100_n274026# 0.010536f
C686 a_n158_n71054# a_n100_n71151# 0.26189f
C687 a_n158_142462# w_n358_n337587# 0.689103f
C688 a_n100_118641# a_n100_121277# 0.205388f
C689 a_n100_n142323# a_n100_n144959# 0.205388f
C690 a_n100_n258307# a_n100_n255671# 0.205388f
C691 a_n100_313705# w_n358_n337587# 0.269531f
C692 a_100_324346# a_100_326982# 0.010536f
C693 a_n158_n139590# w_n358_n337587# 0.689103f
C694 a_n100_171361# a_n158_171458# 0.26189f
C695 a_100_116102# w_n358_n337587# 0.689103f
C696 a_n100_23745# a_100_23842# 0.26189f
C697 a_100_n15698# a_n100_n15795# 0.26189f
C698 a_100_n52602# a_100_n49966# 0.010536f
C699 a_n100_n126507# w_n358_n337587# 0.269531f
C700 a_100_n107958# a_n158_n107958# 0.655843f
C701 a_100_308530# a_100_311166# 0.010536f
C702 a_n158_n23606# a_n100_n23703# 0.26189f
C703 a_100_2754# a_100_118# 0.010536f
C704 a_n158_n129046# a_100_n129046# 0.655843f
C705 a_n100_n65879# a_n100_n68515# 0.205388f
C706 a_100_276898# w_n358_n337587# 0.689103f
C707 a_n100_n139687# a_n158_n139590# 0.26189f
C708 a_n100_n218767# a_n158_n218670# 0.26189f
C709 a_n158_n263482# a_n158_n260846# 0.010536f
C710 a_n100_n113327# w_n358_n337587# 0.269531f
C711 a_100_n39422# w_n358_n337587# 0.689103f
C712 a_n100_68557# a_n100_71193# 0.205388f
C713 a_n158_n324110# a_100_n324110# 0.655843f
C714 a_n100_n324207# a_n100_n326843# 0.205388f
C715 a_100_160914# a_100_163550# 0.010536f
C716 a_100_n226578# a_100_n229214# 0.010536f
C717 a_100_192546# w_n358_n337587# 0.689103f
C718 a_n158_261082# a_n158_263718# 0.010536f
C719 w_n358_n337587# a_n100_n316299# 0.269531f
C720 a_n158_97650# w_n358_n337587# 0.689103f
C721 a_n158_n165950# a_n100_n166047# 0.26189f
C722 a_n158_97650# a_n158_95014# 0.010536f
C723 a_n158_92378# a_n100_92281# 0.26189f
C724 a_n100_147637# a_n100_150273# 0.205388f
C725 a_100_n71054# w_n358_n337587# 0.689103f
C726 a_100_290078# a_100_292714# 0.010536f
C727 a_n158_253174# w_n358_n337587# 0.689103f
C728 a_n100_52741# a_n158_52838# 0.26189f
C729 a_n100_181905# a_n100_184541# 0.205388f
C730 a_n100_118641# a_n158_118738# 0.26189f
C731 a_100_166186# w_n358_n337587# 0.689103f
C732 a_n158_n136954# w_n358_n337587# 0.689103f
C733 a_100_n181766# a_100_n179130# 0.010536f
C734 a_100_79198# a_n158_79198# 0.655843f
C735 a_n100_n115963# a_n100_n113327# 0.205388f
C736 a_n100_297889# w_n358_n337587# 0.269531f
C737 a_n158_58110# w_n358_n337587# 0.689103f
C738 a_n100_216173# w_n358_n337587# 0.269531f
C739 a_n158_n305658# a_n158_n303022# 0.010536f
C740 a_n158_42294# a_100_42294# 0.655843f
C741 a_n158_139826# a_100_139826# 0.655843f
C742 a_n100_166089# a_n100_168725# 0.205388f
C743 a_n158_110830# w_n358_n337587# 0.689103f
C744 a_n158_n155406# a_n158_n152770# 0.010536f
C745 a_n100_n131779# a_n100_n129143# 0.205388f
C746 a_100_n165950# a_100_n168586# 0.010536f
C747 a_100_n179130# a_100_n176494# 0.010536f
C748 a_n158_168822# a_n158_166186# 0.010536f
C749 a_100_n237122# a_n100_n237219# 0.26189f
C750 a_n100_n187135# w_n358_n337587# 0.269531f
C751 w_n358_n337587# a_n158_n324110# 0.689103f
C752 a_100_23842# w_n358_n337587# 0.689103f
C753 a_n158_263718# w_n358_n337587# 0.689103f
C754 a_n158_n26242# w_n358_n337587# 0.689103f
C755 a_n158_160914# w_n358_n337587# 0.689103f
C756 a_100_63382# a_100_66018# 0.010536f
C757 a_100_197818# a_100_195182# 0.010536f
C758 a_100_153006# w_n358_n337587# 0.689103f
C759 a_n158_258446# a_n158_255810# 0.010536f
C760 a_n158_n171222# a_n158_n168586# 0.010536f
C761 a_100_n152770# a_100_n150134# 0.010536f
C762 a_100_81834# w_n358_n337587# 0.689103f
C763 a_n100_329521# a_100_329618# 0.26189f
C764 a_n100_216173# a_n100_213537# 0.205388f
C765 a_n100_n195043# w_n358_n337587# 0.269531f
C766 a_n100_87009# a_n158_87106# 0.26189f
C767 a_100_n92142# a_n158_n92142# 0.655843f
C768 a_n158_n23606# a_n158_n20970# 0.010536f
C769 a_n158_n297750# a_100_n297750# 0.655843f
C770 a_n158_160914# a_n158_163550# 0.010536f
C771 a_n100_231989# w_n358_n337587# 0.269531f
C772 a_n100_n163411# w_n358_n337587# 0.269531f
C773 a_n158_47566# a_n158_44930# 0.010536f
C774 a_100_287442# a_100_284806# 0.010536f
C775 a_n158_124010# w_n358_n337587# 0.689103f
C776 a_100_113466# a_n158_113466# 0.655843f
C777 a_n158_n60510# a_n158_n63146# 0.010536f
C778 a_n100_n121235# a_100_n121138# 0.26189f
C779 a_n100_n110691# a_n158_n110594# 0.26189f
C780 a_n100_n131779# a_n100_n134415# 0.205388f
C781 a_n100_n282031# w_n358_n337587# 0.269531f
C782 a_n158_50202# w_n358_n337587# 0.689103f
C783 a_n100_73829# a_100_73926# 0.26189f
C784 a_n158_n13062# a_n158_n10426# 0.010536f
C785 a_100_n76326# a_100_n73690# 0.010536f
C786 a_n158_15934# a_n158_18570# 0.010536f
C787 a_n100_131821# a_n100_129185# 0.205388f
C788 a_100_224178# a_100_226814# 0.010536f
C789 a_n158_n144862# w_n358_n337587# 0.689103f
C790 a_n100_n81695# a_n100_n79059# 0.205388f
C791 a_n100_7929# w_n358_n337587# 0.269531f
C792 a_n100_134457# w_n358_n337587# 0.269531f
C793 a_100_n192310# w_n358_n337587# 0.689103f
C794 a_n158_250538# a_n158_247902# 0.010536f
C795 a_n158_n263482# a_n158_n266118# 0.010536f
C796 a_n100_250441# a_n100_253077# 0.205388f
C797 a_n158_71290# w_n358_n337587# 0.689103f
C798 a_100_n208126# a_100_n210762# 0.010536f
C799 a_n158_305894# w_n358_n337587# 0.689103f
C800 a_n158_321710# a_n158_319074# 0.010536f
C801 a_n158_210998# a_n100_210901# 0.26189f
C802 a_100_8026# a_n158_8026# 0.655843f
C803 a_n100_137093# a_n100_134457# 0.205388f
C804 a_n158_279534# a_n158_276898# 0.010536f
C805 a_100_n155406# w_n358_n337587# 0.689103f
C806 a_n158_n152770# a_100_n152770# 0.655843f
C807 a_n100_308433# a_n100_305797# 0.205388f
C808 a_100_37022# w_n358_n337587# 0.689103f
C809 a_n158_n226578# a_n158_n223942# 0.010536f
C810 a_100_71290# a_n158_71290# 0.655843f
C811 a_n158_195182# a_n158_197818# 0.010536f
C812 a_n158_124010# a_n158_121374# 0.010536f
C813 a_n100_123913# a_n100_126549# 0.205388f
C814 a_n100_18473# a_n158_18570# 0.26189f
C815 a_100_261082# a_n100_260985# 0.26189f
C816 a_100_89742# w_n358_n337587# 0.689103f
C817 a_n100_n94875# a_n158_n94778# 0.26189f
C818 a_100_2754# w_n358_n337587# 0.689103f
C819 a_n158_239994# w_n358_n337587# 0.689103f
C820 a_n100_47469# a_n100_50105# 0.205388f
C821 a_n100_n229311# a_n100_n231947# 0.205388f
C822 a_100_n28878# a_100_n31514# 0.010536f
C823 a_n100_287345# a_n100_289981# 0.205388f
C824 a_n158_176730# a_n100_176633# 0.26189f
C825 a_100_n221306# a_n100_n221403# 0.26189f
C826 a_100_113466# a_100_116102# 0.010536f
C827 a_100_n26242# a_n158_n26242# 0.655843f
C828 a_n158_313802# a_100_313802# 0.655843f
C829 a_n158_n332018# a_100_n332018# 0.655843f
C830 a_n100_n332115# a_n100_n334751# 0.205388f
C831 a_n100_289981# w_n358_n337587# 0.269531f
C832 a_n100_50105# w_n358_n337587# 0.269531f
C833 w_n358_n337587# a_n100_n305755# 0.269531f
C834 a_100_n284570# w_n358_n337587# 0.689103f
C835 a_n100_200357# a_n100_197721# 0.205388f
C836 a_n100_n102783# a_n158_n102686# 0.26189f
C837 a_n100_n123871# a_n100_n126507# 0.205388f
C838 a_n100_n15795# a_n100_n18431# 0.205388f
C839 a_n100_n247763# a_n100_n250399# 0.205388f
C840 a_100_208362# w_n358_n337587# 0.689103f
C841 a_n158_26478# w_n358_n337587# 0.689103f
C842 a_100_268990# a_n158_268990# 0.655843f
C843 a_n100_n168683# a_100_n168586# 0.26189f
C844 a_n158_232086# a_100_232086# 0.655843f
C845 a_100_303258# a_100_300622# 0.010536f
C846 w_n358_n337587# a_n100_n313663# 0.269531f
C847 a_n158_n73690# w_n358_n337587# 0.689103f
C848 a_100_n258210# a_100_n255574# 0.010536f
C849 a_100_255810# w_n358_n337587# 0.689103f
C850 a_n158_60746# a_100_60746# 0.655843f
C851 a_n100_60649# a_n100_58013# 0.205388f
C852 a_n158_n197582# a_n158_n194946# 0.010536f
C853 a_n100_147637# w_n358_n337587# 0.269531f
C854 a_100_n213398# a_n100_n213495# 0.26189f
C855 a_n158_182002# w_n358_n337587# 0.689103f
C856 a_n100_n110691# w_n358_n337587# 0.269531f
C857 a_100_163550# a_n100_163453# 0.26189f
C858 a_100_n226578# w_n358_n337587# 0.689103f
C859 a_n100_321613# a_n100_324249# 0.205388f
C860 a_n158_n271390# a_n158_n274026# 0.010536f
C861 a_n100_84373# a_n100_87009# 0.205388f
C862 a_100_79198# w_n358_n337587# 0.689103f
C863 a_n100_n260943# a_n158_n260846# 0.26189f
C864 a_n100_n118599# a_n158_n118502# 0.26189f
C865 a_100_282170# a_n100_282073# 0.26189f
C866 a_100_226814# w_n358_n337587# 0.689103f
C867 a_100_174094# a_100_171458# 0.010536f
C868 a_100_105558# a_100_108194# 0.010536f
C869 a_n158_237358# a_n158_234722# 0.010536f
C870 a_n158_23842# a_100_23842# 0.655843f
C871 a_n100_n52699# a_n158_n52602# 0.26189f
C872 a_n158_n63146# a_n100_n63243# 0.26189f
C873 a_n100_42197# w_n358_n337587# 0.269531f
C874 a_n100_76465# a_n158_76562# 0.26189f
C875 a_n100_266257# a_n100_263621# 0.205388f
C876 a_n158_197818# w_n358_n337587# 0.689103f
C877 a_n158_n10426# w_n358_n337587# 0.689103f
C878 w_n358_n337587# a_n158_n321474# 0.689103f
C879 a_100_332254# a_n100_332157# 0.26189f
C880 a_n100_n308391# a_100_n308294# 0.26189f
C881 a_100_97650# w_n358_n337587# 0.689103f
C882 a_n158_n292478# a_n158_n295114# 0.010536f
C883 a_n158_n92142# a_n100_n92239# 0.26189f
C884 a_n100_152909# a_n158_153006# 0.26189f
C885 a_100_253174# w_n358_n337587# 0.689103f
C886 a_100_n28878# w_n358_n337587# 0.689103f
C887 a_100_55474# a_100_52838# 0.010536f
C888 a_100_n276662# w_n358_n337587# 0.689103f
C889 a_n158_n184402# a_n100_n184499# 0.26189f
C890 a_100_290078# a_n158_290078# 0.655843f
C891 w_n358_n337587# a_100_n337290# 0.693647f
C892 a_n158_139826# w_n358_n337587# 0.689103f
C893 a_100_5390# a_n158_5390# 0.655843f
C894 a_100_247902# a_100_250538# 0.010536f
C895 a_n100_118641# a_100_118738# 0.26189f
C896 a_n158_253174# a_n158_250538# 0.010536f
C897 a_100_n268754# w_n358_n337587# 0.689103f
C898 a_100_n221306# w_n358_n337587# 0.689103f
C899 a_n100_n73787# w_n358_n337587# 0.269531f
C900 a_100_297986# w_n358_n337587# 0.689103f
C901 a_n158_210998# a_100_210998# 0.655843f
C902 a_n100_13201# w_n358_n337587# 0.269531f
C903 a_n158_n210762# w_n358_n337587# 0.689103f
C904 a_n158_2754# w_n358_n337587# 0.689103f
C905 a_n100_2657# w_n358_n337587# 0.269531f
C906 a_n100_n284667# a_n100_n287303# 0.205388f
C907 a_n100_n171319# a_n100_n173955# 0.205388f
C908 a_n158_229450# a_n158_226814# 0.010536f
C909 a_n100_195085# a_100_195182# 0.26189f
C910 a_n158_126646# a_n158_124010# 0.010536f
C911 a_100_121374# a_100_124010# 0.010536f
C912 a_100_n310930# a_100_n313566# 0.010536f
C913 a_n100_n313663# a_n158_n313566# 0.26189f
C914 a_100_261082# a_n158_261082# 0.655843f
C915 a_100_189910# w_n358_n337587# 0.689103f
C916 a_100_n234486# w_n358_n337587# 0.689103f
C917 a_100_n295114# a_100_n297750# 0.010536f
C918 a_n100_n297847# a_n158_n297750# 0.26189f
C919 a_n100_n158139# a_n158_n158042# 0.26189f
C920 a_n100_n13159# a_100_n13062# 0.26189f
C921 a_n158_216270# a_100_216270# 0.655843f
C922 a_n158_145098# a_n158_142462# 0.010536f
C923 a_100_147734# a_n100_147637# 0.26189f
C924 a_n100_44833# a_n158_44930# 0.26189f
C925 a_n100_n213495# w_n358_n337587# 0.269531f
C926 a_100_n47330# w_n358_n337587# 0.689103f
C927 a_n100_284709# a_n158_284806# 0.26189f
C928 a_100_n20970# a_n100_n21067# 0.26189f
C929 a_100_124010# w_n358_n337587# 0.689103f
C930 a_n100_n131779# w_n358_n337587# 0.269531f
C931 a_n100_55377# w_n358_n337587# 0.269531f
C932 a_n158_n234486# a_n100_n234583# 0.26189f
C933 a_n158_n121138# a_n158_n118502# 0.010536f
C934 a_n158_n147498# w_n358_n337587# 0.689103f
C935 a_100_n78962# a_n100_n79059# 0.26189f
C936 a_100_134554# a_n158_134554# 0.655843f
C937 a_100_n73690# w_n358_n337587# 0.689103f
C938 a_n100_266257# a_n100_268893# 0.205388f
C939 a_n158_n316202# a_n158_n318838# 0.010536f
C940 a_100_n44694# w_n358_n337587# 0.689103f
C941 a_n100_n47427# a_100_n47330# 0.26189f
C942 a_n100_n274123# a_n158_n274026# 0.26189f
C943 a_n158_295350# a_n158_297986# 0.010536f
C944 a_100_261082# w_n358_n337587# 0.689103f
C945 a_n100_n210859# w_n358_n337587# 0.269531f
C946 a_n100_187177# a_n158_187274# 0.26189f
C947 a_100_184638# a_n158_184638# 0.655843f
C948 a_n158_147734# w_n358_n337587# 0.689103f
C949 a_100_n289842# a_n100_n289939# 0.26189f
C950 a_n100_n39519# a_n100_n36883# 0.205388f
C951 a_n100_116005# a_n158_116102# 0.26189f
C952 a_n100_247805# a_n158_247902# 0.26189f
C953 a_n158_171458# w_n358_n337587# 0.689103f
C954 a_n100_76465# w_n358_n337587# 0.269531f
C955 a_100_305894# w_n358_n337587# 0.689103f
C956 a_100_210998# a_n100_210901# 0.26189f
C957 a_n100_n279395# w_n358_n337587# 0.269531f
C958 a_n158_26478# a_n158_23842# 0.010536f
C959 a_100_282170# a_n158_282170# 0.655843f
C960 a_100_n55238# w_n358_n337587# 0.689103f
C961 a_n100_n292575# w_n358_n337587# 0.269531f
C962 w_n358_n337587# a_n100_n303119# 0.269531f
C963 a_n100_100189# a_n158_100286# 0.26189f
C964 a_100_176730# a_100_174094# 0.010536f
C965 a_n100_n81695# a_n100_n84331# 0.205388f
C966 a_100_n26242# a_100_n28878# 0.010536f
C967 a_n158_n181766# a_n158_n179130# 0.010536f
C968 a_100_42294# w_n358_n337587# 0.689103f
C969 a_n158_308530# a_100_308530# 0.655843f
C970 a_n158_n73690# a_n158_n76326# 0.010536f
C971 a_n158_n5154# a_n158_n7790# 0.010536f
C972 a_n100_n231947# a_n100_n234583# 0.205388f
C973 a_n158_n321474# a_100_n321474# 0.655843f
C974 a_n100_n321571# a_n100_n324207# 0.205388f
C975 a_n100_n21067# a_n100_n23703# 0.205388f
C976 a_n100_n10523# a_n158_n10426# 0.26189f
C977 a_n158_n200218# a_100_n200218# 0.655843f
C978 a_n158_n42058# a_n158_n39422# 0.010536f
C979 a_n158_n94778# w_n358_n337587# 0.689103f
C980 a_n100_n118599# a_n100_n121235# 0.205388f
C981 a_n158_87106# w_n358_n337587# 0.689103f
C982 a_100_218906# a_100_221542# 0.010536f
C983 a_100_n171222# a_100_n168586# 0.010536f
C984 a_n158_147734# a_n158_150370# 0.010536f
C985 a_n158_287442# a_n158_290078# 0.010536f
C986 a_n158_182002# a_n158_179366# 0.010536f
C987 a_100_n247666# w_n358_n337587# 0.689103f
C988 a_n158_n44694# a_100_n44694# 0.655843f
C989 a_100_131918# w_n358_n337587# 0.689103f
C990 a_100_n184402# w_n358_n337587# 0.689103f
C991 a_100_58110# w_n358_n337587# 0.689103f
C992 a_100_n52602# w_n358_n337587# 0.689103f
C993 a_100_n221306# a_100_n218670# 0.010536f
C994 a_100_34386# a_100_37022# 0.010536f
C995 a_n158_31750# a_100_31750# 0.655843f
C996 a_n100_31653# a_n100_29017# 0.205388f
C997 a_n100_100189# w_n358_n337587# 0.269531f
C998 a_100_163550# w_n358_n337587# 0.689103f
C999 a_100_n165950# w_n358_n337587# 0.689103f
C1000 a_100_18570# a_100_15934# 0.010536f
C1001 w_n358_n337587# a_n158_n318838# 0.689103f
C1002 a_n158_n305658# a_n158_n308294# 0.010536f
C1003 a_n100_300525# a_n100_297889# 0.205388f
C1004 a_n158_n192310# a_100_n192310# 0.655843f
C1005 a_n158_63382# a_n100_63285# 0.26189f
C1006 a_100_155642# w_n358_n337587# 0.689103f
C1007 a_n158_n263482# w_n358_n337587# 0.689103f
C1008 a_n158_n289842# w_n358_n337587# 0.689103f
C1009 a_100_182002# w_n358_n337587# 0.689103f
C1010 a_100_163550# a_n158_163550# 0.655843f
C1011 w_n358_n337587# a_100_n334654# 0.689103f
C1012 a_n100_89645# a_n158_89742# 0.26189f
C1013 a_100_n71054# a_n100_n71151# 0.26189f
C1014 a_100_313802# w_n358_n337587# 0.689103f
C1015 a_n100_n229311# a_n100_n226675# 0.205388f
C1016 a_n158_147734# a_100_147734# 0.655843f
C1017 a_100_232086# w_n358_n337587# 0.689103f
C1018 a_n100_n276759# a_n100_n274123# 0.205388f
C1019 a_n100_171361# a_100_171458# 0.26189f
C1020 a_n158_174094# a_n158_176730# 0.010536f
C1021 a_n158_n20970# a_n100_n21067# 0.26189f
C1022 a_n100_113369# w_n358_n337587# 0.269531f
C1023 a_100_237358# a_100_234722# 0.010536f
C1024 a_100_13298# a_100_10662# 0.010536f
C1025 a_n100_10565# a_n158_10662# 0.26189f
C1026 a_n158_n173858# a_n100_n173955# 0.26189f
C1027 a_n158_266354# a_n158_263718# 0.010536f
C1028 a_n100_202993# w_n358_n337587# 0.269531f
C1029 a_n100_158181# a_n158_158278# 0.26189f
C1030 a_n158_n279298# a_n100_n279395# 0.26189f
C1031 a_n100_94917# a_100_95014# 0.26189f
C1032 a_n158_218906# a_n100_218809# 0.26189f
C1033 a_n158_n208126# w_n358_n337587# 0.689103f
C1034 a_n100_152909# a_100_153006# 0.26189f
C1035 a_100_295350# a_100_292714# 0.010536f
C1036 a_n100_250441# w_n358_n337587# 0.269531f
C1037 a_n100_52741# a_n100_50105# 0.205388f
C1038 a_100_n245030# w_n358_n337587# 0.689103f
C1039 a_100_n15698# a_100_n13062# 0.010536f
C1040 a_100_n263482# a_n158_n263482# 0.655843f
C1041 a_n100_n121235# a_n158_n121138# 0.26189f
C1042 a_100_n118502# a_100_n115866# 0.010536f
C1043 a_n100_63285# w_n358_n337587# 0.269531f
C1044 a_n100_321613# a_n158_321710# 0.26189f
C1045 a_n158_13298# w_n358_n337587# 0.689103f
C1046 a_n158_n13062# a_n100_n13159# 0.26189f
C1047 a_n158_42294# a_n158_39658# 0.010536f
C1048 a_100_216270# w_n358_n337587# 0.689103f
C1049 a_100_37022# a_100_39658# 0.010536f
C1050 a_n158_n234486# a_n158_n237122# 0.010536f
C1051 a_n158_n160678# a_n158_n158042# 0.010536f
C1052 a_100_110830# w_n358_n337587# 0.689103f
C1053 a_n100_n55335# a_n100_n52699# 0.205388f
C1054 a_100_n76326# a_100_n78962# 0.010536f
C1055 a_n100_34289# w_n358_n337587# 0.269531f
C1056 a_100_268990# w_n358_n337587# 0.689103f
C1057 a_100_n115866# w_n358_n337587# 0.689103f
C1058 a_n158_195182# a_100_195182# 0.655843f
C1059 a_100_n271390# a_100_n274026# 0.010536f
C1060 a_100_121374# a_n100_121277# 0.26189f
C1061 a_n100_n224039# a_100_n223942# 0.26189f
C1062 a_100_n2518# a_n100_n2615# 0.26189f
C1063 a_n100_n205587# a_100_n205490# 0.26189f
C1064 a_n100_n216131# a_100_n216034# 0.26189f
C1065 a_n158_187274# w_n358_n337587# 0.689103f
C1066 a_100_258446# a_100_255810# 0.010536f
C1067 a_100_n34150# a_n158_n34150# 0.655843f
C1068 a_n100_318977# w_n358_n337587# 0.269531f
C1069 a_n158_329618# a_100_329618# 0.655843f
C1070 a_n100_84373# w_n358_n337587# 0.269531f
C1071 a_n158_324346# a_n100_324249# 0.26189f
C1072 a_n158_89742# a_n158_92378# 0.010536f
C1073 a_n100_n81695# w_n358_n337587# 0.269531f
C1074 a_n100_n31611# a_100_n31514# 0.26189f
C1075 a_n158_n202854# a_n158_n205490# 0.010536f
C1076 a_n100_2657# a_n100_21# 0.205388f
C1077 a_n158_n47330# a_n158_n49966# 0.010536f
C1078 a_n158_n255574# a_n158_n258210# 0.010536f
C1079 a_n100_44833# a_100_44930# 0.26189f
C1080 a_n158_n142226# a_100_n142226# 0.655843f
C1081 a_n100_121277# w_n358_n337587# 0.269531f
C1082 a_n158_n329382# a_100_n329382# 0.655843f
C1083 a_n100_n329479# a_n100_n332115# 0.205388f
C1084 a_n100_245169# a_n100_242533# 0.205388f
C1085 a_n158_239994# a_n158_242630# 0.010536f
C1086 a_n100_n237219# w_n358_n337587# 0.269531f
C1087 a_n100_n115963# a_100_n115866# 0.26189f
C1088 a_100_155642# a_100_158278# 0.010536f
C1089 a_n158_n107958# a_n158_n110594# 0.010536f
C1090 a_100_290078# w_n358_n337587# 0.689103f
C1091 a_n158_55474# w_n358_n337587# 0.689103f
C1092 a_n100_n216131# w_n358_n337587# 0.269531f
C1093 a_100_n279298# w_n358_n337587# 0.689103f
C1094 a_n158_197818# a_n100_197721# 0.26189f
C1095 a_n158_131918# a_n158_129282# 0.010536f
C1096 a_n158_200454# w_n358_n337587# 0.689103f
C1097 a_n158_n276662# w_n358_n337587# 0.689103f
C1098 a_n100_n147595# w_n358_n337587# 0.269531f
C1099 a_100_8026# w_n358_n337587# 0.689103f
C1100 a_n158_n49966# a_n158_n52602# 0.010536f
C1101 a_n100_n168683# w_n358_n337587# 0.269531f
C1102 a_n100_150273# a_100_150370# 0.26189f
C1103 a_n100_n202951# a_n100_n205587# 0.205388f
C1104 w_n358_n337587# a_n100_n311027# 0.269531f
C1105 a_n100_n137051# a_100_n136954# 0.26189f
C1106 a_n158_63382# a_100_63382# 0.655843f
C1107 a_n100_n263579# a_n158_n263482# 0.26189f
C1108 a_n158_n179130# w_n358_n337587# 0.689103f
C1109 a_n100_187177# a_100_187274# 0.26189f
C1110 w_n358_n337587# a_100_n297750# 0.689103f
C1111 a_n100_116005# a_100_116102# 0.26189f
C1112 a_n100_n137051# a_n100_n134415# 0.205388f
C1113 a_100_n123774# a_100_n121138# 0.010536f
C1114 a_100_n258210# w_n358_n337587# 0.689103f
C1115 a_n100_15837# a_n100_13201# 0.205388f
C1116 a_n158_n68418# a_n158_n65782# 0.010536f
C1117 a_n100_n337387# a_100_n337290# 0.26189f
C1118 a_100_n36786# w_n358_n337587# 0.689103f
C1119 a_n158_208362# a_n158_205726# 0.010536f
C1120 a_n158_158278# w_n358_n337587# 0.689103f
C1121 a_n100_221445# w_n358_n337587# 0.269531f
C1122 a_n100_173997# a_100_174094# 0.26189f
C1123 a_n158_n42058# w_n358_n337587# 0.689103f
C1124 a_n158_118738# w_n358_n337587# 0.689103f
C1125 a_100_n287206# a_100_n284570# 0.010536f
C1126 a_100_68654# a_100_66018# 0.010536f
C1127 a_n100_65921# a_n158_66018# 0.26189f
C1128 a_100_282170# w_n358_n337587# 0.689103f
C1129 a_n100_39561# w_n358_n337587# 0.269531f
C1130 a_n100_121277# a_n158_121374# 0.26189f
C1131 a_100_n250302# a_100_n247666# 0.010536f
C1132 a_100_n144862# a_100_n147498# 0.010536f
C1133 a_100_n268754# a_n100_n268851# 0.26189f
C1134 a_100_195182# w_n358_n337587# 0.689103f
C1135 a_n158_21206# w_n358_n337587# 0.689103f
C1136 a_100_329618# w_n358_n337587# 0.689103f
C1137 a_n158_n71054# a_100_n71054# 0.655843f
C1138 a_n158_n57874# a_n158_n55238# 0.010536f
C1139 a_n158_n179130# a_n100_n179227# 0.26189f
C1140 a_100_n300386# a_100_n303022# 0.010536f
C1141 a_n100_n303119# a_n158_n303022# 0.26189f
C1142 a_n100_55377# a_n100_52741# 0.205388f
C1143 w_n358_n337587# a_100_n332018# 0.689103f
C1144 a_n100_n31611# w_n358_n337587# 0.269531f
C1145 a_100_113466# a_n100_113369# 0.26189f
C1146 a_100_n242394# w_n358_n337587# 0.689103f
C1147 a_100_63382# w_n358_n337587# 0.689103f
C1148 a_n100_295253# w_n358_n337587# 0.269531f
C1149 a_n158_n158042# w_n358_n337587# 0.689103f
C1150 a_n158_200454# a_100_200454# 0.655843f
C1151 a_n100_n60607# a_n100_n57971# 0.205388f
C1152 a_100_134554# a_n100_134457# 0.26189f
C1153 a_n100_n200315# a_n158_n200218# 0.26189f
C1154 a_n100_205629# w_n358_n337587# 0.269531f
C1155 a_n158_271626# a_100_271626# 0.655843f
C1156 a_n100_271529# a_n100_268893# 0.205388f
C1157 a_n100_n13159# w_n358_n337587# 0.269531f
C1158 a_n100_n260943# w_n358_n337587# 0.269531f
C1159 a_n100_105461# w_n358_n337587# 0.269531f
C1160 a_n158_15934# a_100_15934# 0.655843f
C1161 a_n158_232086# a_n158_229450# 0.010536f
C1162 a_n158_n44694# a_n158_n42058# 0.010536f
C1163 a_n158_300622# a_100_300622# 0.655843f
C1164 a_100_n239758# a_100_n242394# 0.010536f
C1165 a_100_303258# a_n158_303258# 0.655843f
C1166 a_100_n118502# a_100_n121138# 0.010536f
C1167 a_n158_118738# a_n158_121374# 0.010536f
C1168 a_100_261082# a_100_258446# 0.010536f
C1169 a_n100_253077# a_n100_255713# 0.205388f
C1170 a_n100_179269# w_n358_n337587# 0.269531f
C1171 a_n100_n105419# a_100_n105322# 0.26189f
C1172 a_n100_311069# w_n358_n337587# 0.269531f
C1173 a_n158_84470# w_n358_n337587# 0.689103f
C1174 a_n158_n279298# a_100_n279298# 0.655843f
C1175 a_n158_147734# a_n158_145098# 0.010536f
C1176 a_n158_n276662# a_n158_n279298# 0.010536f
C1177 a_n158_n107958# w_n358_n337587# 0.689103f
C1178 a_n158_n23606# a_n158_n26242# 0.010536f
C1179 a_n100_287345# a_n158_287442# 0.26189f
C1180 a_n100_229353# w_n358_n337587# 0.269531f
C1181 a_n100_n71151# a_n100_n73787# 0.205388f
C1182 a_100_113466# a_100_110830# 0.010536f
C1183 a_100_n121138# w_n358_n337587# 0.689103f
C1184 a_n100_234625# a_100_234722# 0.26189f
C1185 a_100_29114# a_100_31750# 0.010536f
C1186 a_n158_n55238# w_n358_n337587# 0.689103f
C1187 a_n158_287442# w_n358_n337587# 0.689103f
C1188 a_n158_76562# a_100_76562# 0.655843f
C1189 a_n100_76465# a_n100_73829# 0.205388f
C1190 a_100_n205490# a_n158_n205490# 0.655843f
C1191 a_n100_n247763# w_n358_n337587# 0.269531f
C1192 a_n100_202993# a_n158_203090# 0.26189f
C1193 a_n158_n287206# w_n358_n337587# 0.689103f
C1194 a_n100_10565# a_100_10662# 0.26189f
C1195 a_100_13298# a_100_15934# 0.010536f
C1196 a_n100_n192407# a_n100_n195043# 0.205388f
C1197 a_100_n208126# a_100_n205490# 0.010536f
C1198 a_n100_n295211# a_100_n295114# 0.26189f
C1199 a_n100_n166047# w_n358_n337587# 0.269531f
C1200 a_n100_n65879# a_n158_n65782# 0.26189f
C1201 a_n100_n189771# w_n358_n337587# 0.269531f
C1202 a_n158_158278# a_100_158278# 0.655843f
C1203 a_100_266354# a_100_263718# 0.010536f
C1204 a_n100_n195043# a_n158_n194946# 0.26189f
C1205 a_n158_95014# a_100_95014# 0.655843f
C1206 a_n100_94917# a_n100_92281# 0.205388f
C1207 a_100_95014# w_n358_n337587# 0.689103f
C1208 w_n358_n337587# a_n100_334793# 0.349164f
C1209 a_n100_221445# a_n158_221542# 0.26189f
C1210 a_n100_n245127# w_n358_n337587# 0.269531f
C1211 a_n158_292714# a_100_292714# 0.655843f
C1212 a_n100_292617# a_n100_289981# 0.205388f
C1213 a_n158_n268754# a_n158_n266118# 0.010536f
C1214 a_100_n194946# a_100_n197582# 0.010536f
C1215 a_n158_113466# a_n158_116102# 0.010536f
C1216 a_n100_250441# a_n158_250538# 0.26189f
C1217 a_100_n68418# w_n358_n337587# 0.689103f
C1218 a_n158_168822# w_n358_n337587# 0.689103f
C1219 a_n100_308433# w_n358_n337587# 0.269531f
C1220 a_n158_81834# a_100_81834# 0.655843f
C1221 a_n100_81737# a_n100_79101# 0.205388f
C1222 a_n100_68557# w_n358_n337587# 0.269531f
C1223 a_n100_n142323# a_100_n142226# 0.26189f
C1224 a_n158_n179130# a_n158_n176494# 0.010536f
C1225 a_100_42294# a_100_39658# 0.010536f
C1226 a_100_n221306# a_n158_n221306# 0.655843f
C1227 a_100_n258210# a_n100_n258307# 0.26189f
C1228 a_n158_n255574# a_n100_n255671# 0.26189f
C1229 a_n100_n126507# a_100_n126410# 0.26189f
C1230 a_100_105558# a_100_102922# 0.010536f
C1231 a_n100_108097# w_n358_n337587# 0.269531f
C1232 a_n100_226717# a_n158_226814# 0.26189f
C1233 a_n100_n192407# a_100_n192310# 0.26189f
C1234 a_n158_34386# w_n358_n337587# 0.689103f
C1235 a_100_n78962# w_n358_n337587# 0.689103f
C1236 a_n158_n318838# a_100_n318838# 0.655843f
C1237 a_n100_n318935# a_n100_n321571# 0.205388f
C1238 w_n358_n337587# a_n100_n308391# 0.269531f
C1239 a_100_150370# w_n358_n337587# 0.689103f
C1240 a_100_n171222# a_100_n173858# 0.010536f
C1241 a_n158_n47330# w_n358_n337587# 0.689103f
C1242 a_100_187274# w_n358_n337587# 0.689103f
C1243 a_n158_n150134# a_n158_n147498# 0.010536f
C1244 a_n158_319074# w_n358_n337587# 0.689103f
C1245 a_n100_87009# a_100_87106# 0.26189f
C1246 a_100_92378# w_n358_n337587# 0.689103f
C1247 a_100_n89506# a_100_n92142# 0.010536f
C1248 a_n158_n250302# a_n158_n247666# 0.010536f
C1249 a_n100_142365# a_n158_142462# 0.26189f
C1250 a_100_n107958# a_n100_n108055# 0.26189f
C1251 a_100_n171222# w_n358_n337587# 0.689103f
C1252 a_n158_44930# a_100_44930# 0.655843f
C1253 a_100_287442# a_100_290078# 0.010536f
C1254 a_n100_284709# a_n100_282073# 0.205388f
C1255 a_n158_n334654# a_n158_n337290# 0.010536f
C1256 a_n158_110830# a_n158_108194# 0.010536f
C1257 a_n100_n163411# a_n100_n160775# 0.205388f
C1258 a_n158_n223942# w_n358_n337587# 0.689103f
C1259 a_n158_295350# w_n358_n337587# 0.689103f
C1260 a_100_55474# w_n358_n337587# 0.689103f
C1261 a_100_n179130# w_n358_n337587# 0.689103f
C1262 a_n158_203090# a_n158_200454# 0.010536f
C1263 a_100_n18334# a_n158_n18334# 0.655843f
C1264 a_n100_n47427# a_n158_n47330# 0.26189f
C1265 a_n100_n263579# a_n100_n260943# 0.205388f
C1266 a_n158_23842# a_n158_21206# 0.010536f
C1267 a_n100_n13159# a_n100_n10523# 0.205388f
C1268 a_n158_n255574# a_n158_n252938# 0.010536f
C1269 a_n100_n102783# a_n100_n100147# 0.205388f
C1270 a_n100_n26339# a_n100_n28975# 0.205388f
C1271 a_n158_n52602# w_n358_n337587# 0.689103f
C1272 a_n158_n292478# a_n100_n292575# 0.26189f
C1273 a_n100_n155503# a_n100_n158139# 0.205388f
C1274 a_n158_n105322# w_n358_n337587# 0.689103f
C1275 a_n158_5390# a_n158_2754# 0.010536f
C1276 a_n158_29114# a_n158_31750# 0.010536f
C1277 a_100_18570# w_n358_n337587# 0.689103f
C1278 a_n100_34289# a_100_34386# 0.26189f
C1279 w_n358_n337587# a_n100_n297847# 0.269531f
C1280 a_n158_105558# w_n358_n337587# 0.689103f
C1281 a_100_n18334# a_100_n15698# 0.010536f
C1282 a_n158_n71054# a_n158_n73690# 0.010536f
C1283 a_n158_150370# a_100_150370# 0.655843f
C1284 a_n100_n202951# a_n100_n200315# 0.205388f
C1285 a_100_n271390# w_n358_n337587# 0.689103f
C1286 a_n100_145001# w_n358_n337587# 0.269531f
C1287 a_100_118738# a_100_121374# 0.010536f
C1288 a_n100_n258307# a_n100_n260943# 0.205388f
C1289 a_n158_116102# a_100_116102# 0.655843f
C1290 a_n158_10662# a_100_10662# 0.655843f
C1291 w_n358_n337587# a_100_n329382# 0.689103f
C1292 a_100_171458# w_n358_n337587# 0.689103f
C1293 a_n158_n142226# w_n358_n337587# 0.689103f
C1294 a_n100_n137051# w_n358_n337587# 0.269531f
C1295 a_100_76562# w_n358_n337587# 0.689103f
C1296 a_100_311166# w_n358_n337587# 0.689103f
C1297 a_n158_321710# a_n158_324346# 0.010536f
C1298 a_n158_n47330# a_n158_n44694# 0.010536f
C1299 a_100_n213398# a_n158_n213398# 0.655843f
C1300 a_n158_n31514# a_n100_n31611# 0.26189f
C1301 a_n100_173997# a_n100_171361# 0.205388f
C1302 a_n158_276898# a_100_276898# 0.655843f
C1303 a_n158_n18334# w_n358_n337587# 0.689103f
C1304 a_n100_n92239# a_n100_n94875# 0.205388f
C1305 a_n100_n139687# a_n100_n137051# 0.205388f
C1306 a_n100_n97511# a_n158_n97414# 0.26189f
C1307 a_100_118738# w_n358_n337587# 0.689103f
C1308 a_n100_231989# a_n100_234625# 0.205388f
C1309 a_100_n179130# a_n100_n179227# 0.26189f
C1310 a_100_n300386# a_n158_n300386# 0.655843f
C1311 a_n100_n303119# a_n100_n300483# 0.205388f
C1312 a_n100_n210859# a_n100_n208223# 0.205388f
C1313 a_n158_39658# w_n358_n337587# 0.689103f
C1314 a_100_n15698# w_n358_n337587# 0.689103f
C1315 a_n100_192449# a_100_192546# 0.26189f
C1316 a_n158_n115866# a_n158_n118502# 0.010536f
C1317 a_100_155642# a_n100_155545# 0.26189f
C1318 a_100_n310930# a_100_n308294# 0.010536f
C1319 a_n158_n310930# a_n100_n311027# 0.26189f
C1320 a_100_21206# w_n358_n337587# 0.689103f
C1321 a_100_n245030# a_n158_n245030# 0.655843f
C1322 a_100_n57874# a_100_n55238# 0.010536f
C1323 a_100_n144862# a_n100_n144959# 0.26189f
C1324 a_n100_n92239# a_n100_n89603# 0.205388f
C1325 a_n100_n282031# a_n100_n284667# 0.205388f
C1326 a_n158_n36786# a_100_n36786# 0.655843f
C1327 a_n100_n152867# a_100_n152770# 0.26189f
C1328 a_100_n7790# a_n158_n7790# 0.655843f
C1329 a_100_n200218# w_n358_n337587# 0.689103f
C1330 a_100_147734# a_100_150370# 0.010536f
C1331 a_n100_242533# w_n358_n337587# 0.269531f
C1332 a_n158_50202# a_n158_52838# 0.010536f
C1333 a_n158_n281934# a_100_n281934# 0.655843f
C1334 a_n100_n218767# a_n100_n221403# 0.205388f
C1335 a_100_n231850# a_n100_n231947# 0.26189f
C1336 a_n158_n292478# a_n158_n289842# 0.010536f
C1337 a_100_182002# a_100_179366# 0.010536f
C1338 a_n100_179269# a_n158_179366# 0.26189f
C1339 a_n100_n184499# w_n358_n337587# 0.269531f
C1340 a_100_303258# w_n358_n337587# 0.689103f
C1341 a_n100_311069# a_n158_311166# 0.26189f
C1342 a_n100_60649# w_n358_n337587# 0.269531f
C1343 a_n100_131821# a_n100_134457# 0.205388f
C1344 a_100_n102686# a_n158_n102686# 0.655843f
C1345 a_n100_n76423# a_n100_n73787# 0.205388f
C1346 a_n100_n155503# a_n100_n152867# 0.205388f
C1347 a_n100_n229311# a_100_n229214# 0.26189f
C1348 a_100_n92142# w_n358_n337587# 0.689103f
C1349 a_n100_166089# a_100_166186# 0.26189f
C1350 a_100_274262# a_n100_274165# 0.26189f
C1351 a_100_100286# a_100_102922# 0.010536f
C1352 a_n100_110733# w_n358_n337587# 0.269531f
C1353 a_n100_n289939# w_n358_n337587# 0.269531f
C1354 a_100_226814# a_100_229450# 0.010536f
C1355 a_n100_n205587# w_n358_n337587# 0.269531f
C1356 a_n100_266257# w_n358_n337587# 0.269531f
C1357 a_n158_300622# a_n158_297986# 0.010536f
C1358 a_n158_n316202# a_100_n316202# 0.655843f
C1359 a_100_n197582# w_n358_n337587# 0.689103f
C1360 a_n100_258349# a_n100_255713# 0.205388f
C1361 a_n100_316341# w_n358_n337587# 0.269531f
C1362 a_n100_89645# a_n100_87009# 0.205388f
C1363 a_100_84470# w_n358_n337587# 0.689103f
C1364 a_n158_n247666# w_n358_n337587# 0.689103f
C1365 a_n158_229450# w_n358_n337587# 0.689103f
C1366 a_n158_287442# a_100_287442# 0.655843f
C1367 a_n100_47469# a_n158_47566# 0.26189f
C1368 a_n100_n197679# w_n358_n337587# 0.269531f
C1369 a_100_239994# a_n100_239897# 0.26189f
C1370 a_n100_26381# a_n100_29017# 0.205388f
C1371 a_n158_n213398# w_n358_n337587# 0.689103f
C1372 a_n158_47566# w_n358_n337587# 0.689103f
C1373 a_n158_76562# a_n158_73926# 0.010536f
C1374 a_100_134554# a_100_131918# 0.010536f
C1375 a_n100_n36883# w_n358_n337587# 0.269531f
C1376 w_n358_n337587# a_100_334890# 0.693647f
C1377 a_n100_334793# a_n158_334890# 0.26189f
C1378 a_n100_92281# w_n358_n337587# 0.269531f
C1379 a_n158_n7790# w_n358_n337587# 0.689103f
C1380 a_n158_n57874# a_n100_n57971# 0.26189f
C1381 a_100_n260846# a_n158_n260846# 0.655843f
C1382 a_n158_153006# a_100_153006# 0.655843f
C1383 a_n158_n28878# a_n100_n28975# 0.26189f
C1384 a_100_n10426# a_n158_n10426# 0.655843f
C1385 a_100_n284570# a_n100_n284667# 0.26189f
C1386 a_n158_292714# a_n158_290078# 0.010536f
C1387 a_100_250538# w_n358_n337587# 0.689103f
C1388 a_n158_137190# w_n358_n337587# 0.689103f
C1389 a_100_n324110# a_100_n326746# 0.010536f
C1390 a_n100_n218767# w_n358_n337587# 0.269531f
C1391 a_n100_250441# a_n100_247805# 0.205388f
C1392 a_100_176730# w_n358_n337587# 0.689103f
C1393 a_100_n223942# a_100_n226578# 0.010536f
C1394 a_100_5390# a_100_2754# 0.010536f
C1395 a_n100_321613# a_100_321710# 0.26189f
C1396 a_100_210998# a_100_208362# 0.010536f
C1397 a_n100_208265# a_n158_208362# 0.26189f
C1398 a_n158_68654# w_n358_n337587# 0.689103f
C1399 a_100_n158042# a_100_n155406# 0.010536f
C1400 a_n100_n334751# a_100_n334654# 0.26189f
C1401 a_n158_134554# a_n100_134457# 0.26189f
C1402 a_n100_n147595# a_n100_n150231# 0.205388f
C1403 a_100_n65782# a_100_n68418# 0.010536f
C1404 a_100_139826# a_100_137190# 0.010536f
C1405 a_n100_137093# a_n158_137190# 0.26189f
C1406 a_n100_n34247# a_n100_n31611# 0.205388f
C1407 a_100_n289842# a_100_n292478# 0.010536f
C1408 a_100_213634# w_n358_n337587# 0.689103f
C1409 a_n100_n102783# a_100_n102686# 0.26189f
C1410 a_100_37022# a_n158_37022# 0.655843f
C1411 a_n100_39561# a_100_39658# 0.26189f
C1412 a_n100_102825# a_100_102922# 0.26189f
C1413 a_n158_168822# a_n100_168725# 0.26189f
C1414 a_n100_n226675# a_n158_n226578# 0.26189f
C1415 a_n158_n208126# a_n100_n208223# 0.26189f
C1416 a_n100_n118599# a_100_n118502# 0.26189f
C1417 a_n158_10662# a_n158_8026# 0.010536f
C1418 a_100_n237122# a_n158_n237122# 0.655843f
C1419 a_100_n147498# w_n358_n337587# 0.689103f
C1420 a_n100_n253035# a_n100_n250399# 0.205388f
C1421 a_100_n84234# a_100_n81598# 0.010536f
C1422 a_100_303258# a_n100_303161# 0.26189f
C1423 a_n158_n324110# a_n158_n326746# 0.010536f
C1424 a_100_274262# w_n358_n337587# 0.689103f
C1425 w_n358_n337587# a_n100_n295211# 0.269531f
C1426 a_100_n18334# a_n100_n18431# 0.26189f
C1427 a_n100_n5251# a_n100_n2615# 0.205388f
C1428 w_n358_n337587# a_100_n316202# 0.689103f
C1429 a_100_n268754# a_100_n266118# 0.010536f
C1430 a_n100_n163411# a_100_n163314# 0.26189f
C1431 a_n100_5293# w_n358_n337587# 0.269531f
C1432 a_100_n7790# a_n100_n7887# 0.26189f
C1433 a_n100_213537# a_100_213634# 0.26189f
C1434 a_n158_216270# a_n158_218906# 0.010536f
C1435 a_n100_n118599# w_n358_n337587# 0.269531f
C1436 a_n158_237358# w_n358_n337587# 0.689103f
C1437 w_n358_n337587# a_100_n326746# 0.689103f
C1438 a_n100_n142323# w_n358_n337587# 0.269531f
C1439 a_n100_181905# a_n158_182002# 0.26189f
C1440 a_n100_n81695# a_n158_n81598# 0.26189f
C1441 a_n100_126549# w_n358_n337587# 0.269531f
C1442 a_n158_110830# a_n158_113466# 0.010536f
C1443 a_n100_n57971# w_n358_n337587# 0.269531f
C1444 a_100_n60510# a_100_n63146# 0.010536f
C1445 a_n100_n7887# a_n100_n5251# 0.205388f
C1446 a_100_n305658# a_100_n303022# 0.010536f
C1447 a_n158_n305658# a_n100_n305755# 0.26189f
C1448 a_n158_n155406# w_n358_n337587# 0.689103f
C1449 a_n100_n152867# a_n158_n152770# 0.26189f
C1450 a_100_295350# w_n358_n337587# 0.689103f
C1451 a_100_311166# a_n158_311166# 0.655843f
C1452 a_n158_316438# a_n158_313802# 0.010536f
C1453 a_100_n221306# a_100_n223942# 0.010536f
C1454 a_100_131918# a_100_129282# 0.010536f
C1455 a_n100_n139687# a_n100_n142323# 0.205388f
C1456 a_n158_34386# a_100_34386# 0.655843f
C1457 a_n100_34289# a_n100_31653# 0.205388f
C1458 a_n158_274262# a_100_274262# 0.655843f
C1459 a_n158_15934# w_n358_n337587# 0.689103f
C1460 a_n100_n18431# w_n358_n337587# 0.269531f
C1461 a_100_205726# w_n358_n337587# 0.689103f
C1462 a_n158_n113230# a_100_n113230# 0.655843f
C1463 a_100_n189674# a_100_n192310# 0.010536f
C1464 w_n358_n337587# a_n100_n326843# 0.269531f
C1465 a_100_105558# w_n358_n337587# 0.689103f
C1466 a_n100_n118599# a_n100_n115963# 0.205388f
C1467 a_n158_n68418# w_n358_n337587# 0.689103f
C1468 a_n158_n15698# a_n158_n18334# 0.010536f
C1469 a_100_n171222# a_n158_n171222# 0.655843f
C1470 a_n158_63382# a_n158_60746# 0.010536f
C1471 a_n158_n268754# w_n358_n337587# 0.689103f
C1472 a_n100_255713# w_n358_n337587# 0.269531f
C1473 a_n158_253174# a_n158_255810# 0.010536f
C1474 a_n100_116005# a_n100_113369# 0.205388f
C1475 a_n100_n44791# w_n358_n337587# 0.269531f
C1476 a_n158_n15698# a_100_n15698# 0.655843f
C1477 a_n158_n281934# a_n158_n284570# 0.010536f
C1478 a_100_321710# a_100_319074# 0.010536f
C1479 a_n158_n297750# a_n158_n300386# 0.010536f
C1480 a_n158_73926# w_n358_n337587# 0.689103f
C1481 a_n158_42294# a_n158_44930# 0.010536f
C1482 a_n100_n2615# w_n358_n337587# 0.269531f
C1483 a_n100_n92239# w_n358_n337587# 0.269531f
C1484 a_n158_n205490# w_n358_n337587# 0.689103f
C1485 a_n100_237261# a_n158_237358# 0.26189f
C1486 a_100_29114# a_n158_29114# 0.655843f
C1487 a_100_13298# w_n358_n337587# 0.689103f
C1488 a_100_279534# w_n358_n337587# 0.689103f
C1489 a_n100_n55335# w_n358_n337587# 0.269531f
C1490 a_n158_n139590# a_n158_n136954# 0.010536f
C1491 a_n100_36925# w_n358_n337587# 0.269531f
C1492 a_n100_n47427# a_n100_n44791# 0.205388f
C1493 a_100_n208126# w_n358_n337587# 0.689103f
C1494 a_n158_n115866# a_n158_n113230# 0.010536f
C1495 a_n158_n245030# a_n100_n245127# 0.26189f
C1496 a_n100_n229311# w_n358_n337587# 0.269531f
C1497 a_n100_18473# w_n358_n337587# 0.269531f
C1498 a_n158_329618# a_n158_332254# 0.010536f
C1499 a_100_87106# w_n358_n337587# 0.689103f
C1500 a_n158_n189674# a_n158_n187038# 0.010536f
C1501 a_100_n78962# a_n158_n78962# 0.655843f
C1502 a_n100_n7887# w_n358_n337587# 0.269531f
C1503 a_n100_n68515# w_n358_n337587# 0.269531f
C1504 a_n100_179269# a_100_179366# 0.26189f
C1505 a_n158_129282# w_n358_n337587# 0.689103f
C1506 a_n158_60746# w_n358_n337587# 0.689103f
C1507 a_n158_n84234# a_n158_n86870# 0.010536f
C1508 a_n158_n121138# w_n358_n337587# 0.689103f
C1509 a_100_n152770# w_n358_n337587# 0.689103f
C1510 a_n100_n218767# a_100_n218670# 0.26189f
C1511 a_n158_205726# w_n358_n337587# 0.689103f
C1512 a_n158_n44694# a_n100_n44791# 0.26189f
C1513 a_n100_271529# a_n100_274165# 0.205388f
C1514 a_100_n81598# w_n358_n337587# 0.689103f
C1515 a_100_n94778# a_n158_n94778# 0.655843f
C1516 a_100_100286# a_n158_100286# 0.655843f
C1517 a_100_232086# a_100_229450# 0.010536f
C1518 a_n158_300622# a_n158_303258# 0.010536f
C1519 a_100_266354# w_n358_n337587# 0.689103f
C1520 a_n100_n200315# w_n358_n337587# 0.269531f
C1521 a_100_n287206# a_n158_n287206# 0.655843f
C1522 a_n100_n155503# w_n358_n337587# 0.269531f
C1523 a_n100_321613# w_n358_n337587# 0.269531f
C1524 a_n100_81737# w_n358_n337587# 0.269531f
C1525 a_100_n131682# a_n158_n131682# 0.655843f
C1526 a_n100_145001# a_n158_145098# 0.26189f
C1527 a_100_n281934# w_n358_n337587# 0.689103f
C1528 a_n158_282170# a_n158_284806# 0.010536f
C1529 a_n100_287345# a_n100_284709# 0.205388f
C1530 a_n100_n65879# w_n358_n337587# 0.269531f
C1531 a_n100_47469# a_n100_44833# 0.205388f
C1532 a_n158_n332018# a_n158_n334654# 0.010536f
C1533 a_100_126646# w_n358_n337587# 0.689103f
C1534 a_n100_284709# w_n358_n337587# 0.269531f
C1535 a_n100_44833# w_n358_n337587# 0.269531f
C1536 a_n158_n100050# a_n158_n102686# 0.010536f
C1537 a_n100_n276759# a_100_n276662# 0.26189f
C1538 a_n100_131821# a_100_131918# 0.26189f
C1539 a_n100_21109# a_n158_21206# 0.26189f
C1540 a_100_203090# w_n358_n337587# 0.689103f
C1541 a_n100_263621# a_100_263718# 0.26189f
C1542 a_n100_n171319# w_n358_n337587# 0.269531f
C1543 a_n100_n324207# a_100_n324110# 0.26189f
C1544 a_n158_n102686# w_n358_n337587# 0.689103f
C1545 a_n100_160817# a_100_160914# 0.26189f
C1546 a_100_100286# w_n358_n337587# 0.689103f
C1547 a_n158_334890# a_100_334890# 0.655843f
C1548 w_n358_n337587# a_n158_332254# 0.689103f
C1549 a_n100_334793# a_n100_332157# 0.205388f
C1550 w_n358_n337587# a_100_n313566# 0.689103f
C1551 a_n100_221445# a_100_221542# 0.26189f
C1552 a_n100_n97511# a_n100_n100147# 0.205388f
C1553 a_n100_n110691# a_100_n110594# 0.26189f
C1554 a_n100_292617# a_n100_295253# 0.205388f
C1555 a_n100_n271487# w_n358_n337587# 0.269531f
C1556 a_n158_189910# a_100_189910# 0.655843f
C1557 a_100_n213398# a_100_n210762# 0.010536f
C1558 a_100_137190# w_n358_n337587# 0.689103f
C1559 a_n100_173997# w_n358_n337587# 0.269531f
C1560 a_n158_250538# a_100_250538# 0.655843f
C1561 a_n158_308530# w_n358_n337587# 0.689103f
C1562 a_n100_n181863# a_n100_n184499# 0.205388f
C1563 a_100_68654# w_n358_n337587# 0.689103f
C1564 a_n100_137093# a_100_137190# 0.26189f
C1565 a_100_29114# a_100_26478# 0.010536f
C1566 a_n100_26381# a_n158_26478# 0.26189f
C1567 a_n158_n36786# a_n100_n36883# 0.26189f
C1568 a_100_n150134# w_n358_n337587# 0.689103f
C1569 a_n100_274165# a_n100_276801# 0.205388f
C1570 a_n158_218906# w_n358_n337587# 0.689103f
C1571 a_n100_279437# a_100_279534# 0.26189f
C1572 a_n158_39658# a_100_39658# 0.655843f
C1573 a_n100_n60607# a_100_n60510# 0.26189f
C1574 a_n158_232086# a_n158_234722# 0.010536f
C1575 a_n158_31750# w_n358_n337587# 0.689103f
C1576 a_n100_271529# w_n358_n337587# 0.269531f
C1577 a_100_71290# a_100_68654# 0.010536f
C1578 a_n100_n144959# w_n358_n337587# 0.269531f
C1579 a_n100_63285# a_n100_65921# 0.205388f
C1580 a_n100_n239855# w_n358_n337587# 0.269531f
C1581 w_n358_n337587# a_n100_n324207# 0.269531f
C1582 a_n158_255810# a_100_255810# 0.655843f
C1583 a_n158_184638# w_n358_n337587# 0.689103f
C1584 a_n158_126646# a_n100_126549# 0.26189f
C1585 a_100_n292478# a_100_n295114# 0.010536f
C1586 a_100_319074# w_n358_n337587# 0.689103f
C1587 a_100_329618# a_100_326982# 0.010536f
C1588 a_n100_89645# w_n358_n337587# 0.269531f
C1589 a_n100_n7887# a_n100_n10523# 0.205388f
C1590 a_n158_n86870# w_n358_n337587# 0.689103f
C1591 a_n158_213634# a_100_213634# 0.655843f
C1592 a_n158_n189674# w_n358_n337587# 0.689103f
C1593 a_n158_n200218# a_n158_n202854# 0.010536f
C1594 a_n100_181905# a_100_182002# 0.26189f
C1595 a_n100_242533# a_n158_242630# 0.26189f
C1596 a_100_n239758# a_n100_n239855# 0.26189f
C1597 a_n158_n34150# w_n358_n337587# 0.689103f
C1598 a_100_316438# a_100_313802# 0.010536f
C1599 a_n158_292714# w_n358_n337587# 0.689103f
C1600 a_100_203090# a_100_200454# 0.010536f
C1601 a_n158_n242394# w_n358_n337587# 0.689103f
C1602 a_100_n258210# a_n158_n258210# 0.655843f
C1603 a_n100_n102783# w_n358_n337587# 0.269531f
C1604 a_n158_n223942# a_n158_n221306# 0.010536f
C1605 a_n158_n86870# a_100_n86870# 0.655843f
C1606 a_n158_224178# a_n158_226814# 0.010536f
C1607 a_n100_102825# w_n358_n337587# 0.269531f
C1608 a_100_n131682# a_100_n134318# 0.010536f
C1609 a_n158_n160678# a_100_n160678# 0.655843f
C1610 a_n158_n163314# a_n158_n165950# 0.010536f
C1611 a_n158_n234486# w_n358_n337587# 0.689103f
C1612 a_n100_n276759# a_n100_n279395# 0.205388f
C1613 a_n158_n287206# a_n100_n287303# 0.26189f
C1614 a_n100_n110691# a_n100_n113327# 0.205388f
C1615 a_n100_n297847# a_n100_n300483# 0.205388f
C1616 a_n100_187177# a_n100_189813# 0.205388f
C1617 a_n158_n152770# w_n358_n337587# 0.689103f
C1618 a_n158_n313566# a_100_n313566# 0.655843f
C1619 a_n100_n313663# a_n100_n316299# 0.205388f
C1620 a_n100_n34247# a_n100_n36883# 0.205388f
C1621 a_n100_n216131# a_n158_n216034# 0.26189f
C1622 a_100_n271390# a_n158_n271390# 0.655843f
C1623 a_n100_n42155# a_n158_n42058# 0.26189f
C1624 a_n158_n245030# a_n158_n247666# 0.010536f
C1625 a_n158_316438# w_n358_n337587# 0.689103f
C1626 a_n158_n218670# w_n358_n337587# 0.689103f
C1627 a_100_n181766# a_n158_n181766# 0.655843f
C1628 a_n158_139826# a_n158_142462# 0.010536f
C1629 a_n158_155642# w_n358_n337587# 0.689103f
C1630 a_100_n210762# w_n358_n337587# 0.689103f
C1631 a_n158_174094# a_n158_171458# 0.010536f
C1632 a_n100_n234583# w_n358_n337587# 0.269531f
C1633 a_n100_10565# w_n358_n337587# 0.269531f
C1634 a_n100_276801# w_n358_n337587# 0.269531f
C1635 a_n158_126646# a_n158_129282# 0.010536f
C1636 a_n100_266257# a_n158_266354# 0.26189f
C1637 a_100_n316202# a_100_n318838# 0.010536f
C1638 a_n158_18570# w_n358_n337587# 0.689103f
C1639 a_n100_324249# w_n358_n337587# 0.269531f
C1640 a_n158_218906# a_n158_221542# 0.010536f
C1641 a_n158_97650# a_100_97650# 0.655843f
C1642 a_n100_97553# a_n100_94917# 0.205388f
C1643 a_n100_224081# a_n100_221445# 0.205388f
C1644 a_n158_n134318# a_n158_n131682# 0.010536f
C1645 a_n158_92378# a_n158_95014# 0.010536f
C1646 a_n158_92378# w_n358_n337587# 0.689103f
C1647 a_n100_21# a_n100_n2615# 0.205388f
C1648 a_n158_50202# a_n100_50105# 0.26189f
C1649 a_n100_n231947# w_n358_n337587# 0.269531f
C1650 a_n100_239897# w_n358_n337587# 0.269531f
C1651 a_n158_55474# a_n158_52838# 0.010536f
C1652 a_n100_179269# a_n100_176633# 0.205388f
C1653 a_100_168822# w_n358_n337587# 0.689103f
C1654 a_n158_253174# a_100_253174# 0.655843f
C1655 a_n158_n284570# w_n358_n337587# 0.689103f
C1656 a_n100_n189771# a_n100_n192407# 0.205388f
C1657 a_n158_n20970# a_n158_n18334# 0.010536f
C1658 a_n158_84470# a_n158_81834# 0.010536f
C1659 a_n100_n173955# a_100_n173858# 0.26189f
C1660 a_n100_n332115# a_100_n332018# 0.26189f
C1661 a_100_79198# a_100_81834# 0.010536f
C1662 a_100_60746# w_n358_n337587# 0.689103f
C1663 a_n158_300622# w_n358_n337587# 0.689103f
C1664 a_n100_15837# a_n158_15934# 0.26189f
C1665 a_n158_203090# a_n158_205726# 0.010536f
C1666 w_n358_n337587# a_100_n303022# 0.689103f
C1667 a_100_n163314# a_100_n165950# 0.010536f
C1668 a_n158_n173858# a_100_n173858# 0.655843f
C1669 a_n158_n121138# a_n158_n123774# 0.010536f
C1670 a_n100_268893# a_n158_268990# 0.26189f
C1671 a_n100_229353# a_100_229450# 0.26189f
C1672 a_n100_n173955# w_n358_n337587# 0.269531f
C1673 a_n158_n321474# a_n158_n324110# 0.010536f
C1674 a_n100_297889# a_100_297986# 0.26189f
C1675 a_100_189910# a_100_192546# 0.010536f
C1676 a_n158_n173858# w_n358_n337587# 0.689103f
C1677 w_n358_n337587# a_100_n310930# 0.689103f
C1678 a_100_8026# a_100_5390# 0.010536f
C1679 a_n158_126646# a_100_126646# 0.655843f
C1680 a_n158_n276662# a_n158_n274026# 0.010536f
C1681 a_n158_n229214# a_n100_n229311# 0.26189f
C1682 a_100_184638# w_n358_n337587# 0.689103f
C1683 a_n100_n28975# w_n358_n337587# 0.269531f
C1684 a_100_218906# a_100_216270# 0.010536f
C1685 a_100_n42058# w_n358_n337587# 0.689103f
C1686 a_n100_160817# a_n100_163453# 0.205388f
C1687 a_n100_145001# a_100_145098# 0.26189f
C1688 a_100_n260846# w_n358_n337587# 0.689103f
C1689 a_n158_47566# a_100_47566# 0.655843f
C1690 a_n100_226717# w_n358_n337587# 0.269531f
C1691 a_100_176730# a_100_179366# 0.010536f
C1692 a_n100_123913# w_n358_n337587# 0.269531f
C1693 a_n100_237261# a_n100_239897# 0.205388f
C1694 a_n100_n65879# a_100_n65782# 0.26189f
C1695 a_n100_n202951# a_n158_n202854# 0.26189f
C1696 a_n158_n268754# a_n100_n268851# 0.26189f
C1697 a_n100_n205587# a_n100_n208223# 0.205388f
C1698 a_n158_308530# a_n158_311166# 0.010536f
C1699 a_n100_73829# a_n158_73926# 0.26189f
C1700 a_n158_284806# w_n358_n337587# 0.689103f
C1701 a_n158_44930# w_n358_n337587# 0.689103f
C1702 a_100_n160678# w_n358_n337587# 0.689103f
C1703 a_n158_203090# a_100_203090# 0.655843f
C1704 a_n100_202993# a_n100_200357# 0.205388f
C1705 a_n100_126549# a_n100_129185# 0.205388f
C1706 a_n100_15837# a_n100_18473# 0.205388f
C1707 a_n100_21109# a_100_21206# 0.26189f
C1708 a_n100_263621# a_n100_260985# 0.205388f
C1709 a_n100_n15795# w_n358_n337587# 0.269531f
C1710 a_100_n71054# a_100_n73690# 0.010536f
C1711 w_n358_n337587# a_n100_n321571# 0.269531f
C1712 a_n158_334890# a_n158_332254# 0.010536f
C1713 a_100_n305658# a_100_n308294# 0.010536f
C1714 a_n100_n308391# a_n158_n308294# 0.26189f
C1715 a_n158_10662# w_n358_n337587# 0.689103f
C1716 a_n158_189910# a_n158_187274# 0.010536f
C1717 a_100_n97414# a_n158_n97414# 0.655843f
C1718 a_n158_118738# a_n158_116102# 0.010536f
C1719 a_100_n252938# a_n100_n253035# 0.26189f
C1720 a_100_n136954# a_100_n134318# 0.010536f
C1721 a_n158_113466# a_n100_113369# 0.26189f
C1722 a_n100_n97511# a_n100_n94875# 0.205388f
C1723 w_n358_n337587# a_n158_n337290# 0.693647f
C1724 a_n158_n100050# a_n158_n97414# 0.010536f
C1725 a_n158_n181766# a_n158_n184402# 0.010536f
C1726 a_100_n134318# a_n100_n134415# 0.26189f
C1727 a_n158_321710# a_100_321710# 0.655843f
C1728 a_100_308530# w_n358_n337587# 0.689103f
C1729 a_n100_n171319# a_n158_n171222# 0.26189f
C1730 a_n158_n97414# w_n358_n337587# 0.689103f
C1731 a_n158_n168586# a_n100_n168683# 0.26189f
C1732 a_100_n134318# a_n158_n134318# 0.655843f
C1733 a_n158_279534# a_100_279534# 0.655843f
C1734 a_n100_279437# a_n100_276801# 0.205388f
C1735 a_n158_n92142# w_n358_n337587# 0.689103f
C1736 a_100_118# a_n158_118# 0.655843f
C1737 a_100_n118502# a_n158_n118502# 0.655843f
C1738 a_100_n34150# a_100_n31514# 0.010536f
C1739 a_n100_n39519# a_n158_n39422# 0.26189f
C1740 a_n158_n31514# a_n158_n34150# 0.010536f
C1741 a_100_n218670# a_n158_n218670# 0.655843f
C1742 a_100_232086# a_100_234722# 0.010536f
C1743 a_100_108194# w_n358_n337587# 0.689103f
C1744 a_100_n263482# a_100_n260846# 0.010536f
C1745 a_n100_68557# a_n100_65921# 0.205388f
C1746 a_100_31750# w_n358_n337587# 0.689103f
C1747 a_n100_n108055# w_n358_n337587# 0.269531f
C1748 a_n158_195182# a_n158_192546# 0.010536f
C1749 a_n158_124010# a_100_124010# 0.655843f
C1750 a_n100_189813# w_n358_n337587# 0.269531f
C1751 a_n100_n289939# a_n100_n287303# 0.205388f
C1752 a_100_329618# a_100_332254# 0.010536f
C1753 a_n158_89742# w_n358_n337587# 0.689103f
C1754 a_n158_324346# w_n358_n337587# 0.689103f
C1755 a_n100_326885# a_n100_324249# 0.205388f
C1756 a_n158_n118502# w_n358_n337587# 0.689103f
C1757 a_n158_234722# w_n358_n337587# 0.689103f
C1758 a_100_50202# a_100_52838# 0.010536f
C1759 a_n100_181905# a_n100_179269# 0.205388f
C1760 a_n158_n158042# a_100_n158042# 0.655843f
C1761 a_n100_108097# a_n158_108194# 0.26189f
C1762 a_n100_n276759# a_n158_n276662# 0.26189f
C1763 a_n100_160817# a_n100_158181# 0.205388f
C1764 a_n100_242533# a_100_242630# 0.26189f
C1765 a_n100_313705# a_100_313802# 0.26189f
C1766 a_n158_n184402# a_n158_n187038# 0.010536f
C1767 a_n158_n237122# w_n358_n337587# 0.689103f
C1768 a_n100_200357# a_n158_200454# 0.26189f
C1769 a_n100_129185# a_n158_129282# 0.26189f
C1770 a_100_n181766# w_n358_n337587# 0.689103f
C1771 a_100_n176494# a_100_n173858# 0.010536f
C1772 a_n158_n147498# a_n158_n144862# 0.010536f
C1773 a_n100_208265# w_n358_n337587# 0.269531f
C1774 a_100_29114# w_n358_n337587# 0.689103f
C1775 a_100_268990# a_100_271626# 0.010536f
C1776 a_n100_2657# a_100_2754# 0.26189f
C1777 a_100_2754# a_n158_2754# 0.655843f
C1778 a_n100_n253035# w_n358_n337587# 0.269531f
C1779 a_100_58110# a_n158_58110# 0.655843f
C1780 a_100_n57874# a_n100_n57971# 0.26189f
C1781 a_n100_n279395# a_n100_n282031# 0.205388f
C1782 a_n100_184541# a_n158_184638# 0.26189f
C1783 a_n158_n36786# a_n158_n34150# 0.010536f
C1784 a_n158_n268754# a_n158_n271390# 0.010536f
C1785 a_100_n176494# w_n358_n337587# 0.689103f
C1786 a_100_253174# a_100_255810# 0.010536f
C1787 a_n100_5293# a_n158_5390# 0.26189f
C1788 a_100_n292478# w_n358_n337587# 0.689103f
C1789 a_100_163550# a_100_166186# 0.010536f
C1790 a_n100_71193# w_n358_n337587# 0.269531f
C1791 a_n100_n68515# a_n100_n71151# 0.205388f
C1792 a_n158_n173858# a_n158_n176494# 0.010536f
C1793 a_100_282170# a_100_284806# 0.010536f
C1794 a_n158_n73690# a_n100_n73787# 0.26189f
C1795 a_n100_218809# w_n358_n337587# 0.269531f
C1796 a_100_176730# a_n158_176730# 0.655843f
C1797 a_n158_n329382# a_n158_n332018# 0.010536f
C1798 a_n158_105558# a_n158_108194# 0.010536f
C1799 w_n358_n337587# a_100_n300386# 0.689103f
C1800 a_n158_n197582# a_100_n197582# 0.655843f
C1801 a_n158_237358# a_100_237358# 0.655843f
C1802 a_100_n34150# w_n358_n337587# 0.689103f
C1803 a_n158_305894# a_100_305894# 0.655843f
C1804 a_100_n223942# a_n158_n223942# 0.655843f
C1805 a_n100_n271487# a_n100_n268851# 0.205388f
C1806 a_100_71290# a_n100_71193# 0.26189f
C1807 a_n100_n197679# a_n158_n197582# 0.26189f
C1808 a_n100_n321571# a_100_n321474# 0.26189f
C1809 a_n158_266354# a_100_266354# 0.655843f
C1810 a_n158_n131682# w_n358_n337587# 0.689103f
C1811 a_n158_192546# w_n358_n337587# 0.689103f
C1812 a_n100_97553# w_n358_n337587# 0.269531f
C1813 a_100_118# a_100_n2518# 0.010536f
C1814 a_n158_n189674# a_n158_n192310# 0.010536f
C1815 a_n158_n234486# a_n158_n231850# 0.010536f
C1816 a_100_155642# a_100_153006# 0.010536f
C1817 w_n358_n337587# a_n158_n300386# 0.689103f
C1818 a_n158_n165950# w_n358_n337587# 0.689103f
C1819 a_100_247902# w_n358_n337587# 0.689103f
C1820 a_n158_166186# w_n358_n337587# 0.689103f
C1821 a_100_n107958# w_n358_n337587# 0.689103f
C1822 a_100_300622# w_n358_n337587# 0.689103f
C1823 a_n100_58013# w_n358_n337587# 0.269531f
C1824 a_100_n208126# a_n100_n208223# 0.26189f
C1825 a_n158_n113230# a_n158_n110594# 0.010536f
C1826 a_100_n200218# a_100_n202854# 0.010536f
C1827 a_100_n60510# w_n358_n337587# 0.689103f
C1828 a_100_n231850# a_100_n229214# 0.010536f
C1829 a_n100_139729# a_100_139826# 0.26189f
C1830 a_100_n113230# w_n358_n337587# 0.689103f
C1831 a_n158_166186# a_n158_163550# 0.010536f
C1832 a_n158_34386# a_n158_37022# 0.010536f
C1833 a_100_168822# a_n100_168725# 0.26189f
C1834 a_n100_n34247# a_n158_n34150# 0.26189f
C1835 a_n158_n73690# a_100_n73690# 0.655843f
C1836 a_n158_229450# a_100_229450# 0.655843f
C1837 a_100_232086# a_n100_231989# 0.26189f
C1838 a_n158_n81598# a_100_n81598# 0.655843f
C1839 a_n100_263621# w_n358_n337587# 0.269531f
C1840 a_n158_n250302# a_n100_n250399# 0.26189f
C1841 w_n358_n337587# a_n100_n318935# 0.269531f
C1842 a_n100_160817# w_n358_n337587# 0.269531f
C1843 a_n100_n242491# a_100_n242394# 0.26189f
C1844 a_n158_118# w_n358_n337587# 0.689103f
C1845 a_n158_321710# w_n358_n337587# 0.689103f
C1846 a_n100_329521# a_n158_329618# 0.26189f
C1847 a_n158_n303022# a_100_n303022# 0.655843f
C1848 a_n100_n303119# a_n100_n305755# 0.205388f
C1849 a_n100_216173# a_100_216270# 0.26189f
C1850 w_n358_n337587# a_n158_n334654# 0.689103f
C1851 a_100_n187038# a_n158_n187038# 0.655843f
C1852 a_n158_n226578# w_n358_n337587# 0.689103f
C1853 a_n100_n150231# a_100_n150134# 0.26189f
C1854 a_n158_n49966# a_100_n49966# 0.655843f
C1855 a_n100_n231947# a_n158_n231850# 0.26189f
C1856 a_n158_147734# a_n100_147637# 0.26189f
C1857 a_n158_n5154# a_n100_n5251# 0.26189f
C1858 a_n158_n15698# a_n100_n15795# 0.26189f
C1859 a_n100_n105419# a_n158_n105322# 0.26189f
C1860 a_n100_145001# a_n100_142365# 0.205388f
C1861 a_n100_n224039# a_n158_n223942# 0.26189f
C1862 a_n100_2657# a_n158_2754# 0.26189f
C1863 a_n158_282170# a_n100_282073# 0.26189f
C1864 a_n158_226814# w_n358_n337587# 0.689103f
C1865 a_100_n144862# a_100_n142226# 0.010536f
C1866 a_n100_n226675# w_n358_n337587# 0.269531f
C1867 a_100_176730# a_n100_176633# 0.26189f
C1868 a_n100_n189771# a_100_n189674# 0.26189f
C1869 a_100_n92142# a_100_n94778# 0.010536f
C1870 a_n158_n242394# a_n158_n245030# 0.010536f
C1871 a_n158_110830# a_100_110830# 0.655843f
C1872 a_n158_n171222# a_n158_n173858# 0.010536f
C1873 a_100_44930# w_n358_n337587# 0.689103f
C1874 a_100_76562# a_100_73926# 0.010536f
C1875 a_n158_n184402# w_n358_n337587# 0.689103f
C1876 a_n158_n115866# w_n358_n337587# 0.689103f
C1877 a_n100_21109# a_n100_18473# 0.205388f
C1878 a_n100_n121235# w_n358_n337587# 0.269531f
C1879 a_n100_n97511# a_100_n97414# 0.26189f
C1880 a_n158_n71054# a_n158_n68418# 0.010536f
C1881 a_n100_332157# a_n158_332254# 0.26189f
C1882 a_n158_n150134# a_100_n150134# 0.655843f
C1883 a_n158_55474# a_n158_58110# 0.010536f
C1884 a_n158_n310930# a_100_n310930# 0.655843f
C1885 a_100_184638# a_n100_184541# 0.26189f
C1886 a_100_10662# w_n358_n337587# 0.689103f
C1887 a_n100_n97511# w_n358_n337587# 0.269531f
C1888 a_n158_n213398# a_n158_n216034# 0.010536f
C1889 a_n100_n266215# a_n158_n266118# 0.26189f
C1890 a_100_n39422# a_100_n36786# 0.010536f
C1891 a_n100_n271487# a_n158_n271390# 0.26189f
C1892 a_n100_n73787# a_100_n73690# 0.26189f
C1893 a_100_174094# w_n358_n337587# 0.689103f
C1894 a_n100_n39519# w_n358_n337587# 0.269531f
C1895 a_100_66018# w_n358_n337587# 0.689103f
C1896 a_n100_305797# w_n358_n337587# 0.269531f
C1897 a_n100_79101# a_n158_79198# 0.26189f
C1898 a_n100_n115963# a_n158_n115866# 0.26189f
C1899 a_100_139826# a_100_142462# 0.010536f
C1900 a_100_n134318# w_n358_n337587# 0.689103f
C1901 a_100_n176494# a_n158_n176494# 0.655843f
C1902 a_n158_39658# a_n158_37022# 0.010536f
C1903 a_100_42294# a_n100_42197# 0.26189f
C1904 a_n100_n26339# w_n358_n337587# 0.269531f
C1905 a_n100_n210859# a_n158_n210762# 0.26189f
C1906 a_n100_n242491# a_n100_n245127# 0.205388f
C1907 a_n100_118641# w_n358_n337587# 0.269531f
C1908 a_n100_268893# w_n358_n337587# 0.269531f
C1909 a_n158_n5154# w_n358_n337587# 0.689103f
C1910 a_100_195182# a_100_192546# 0.010536f
C1911 a_100_197818# w_n358_n337587# 0.689103f
C1912 a_100_n63146# w_n358_n337587# 0.689103f
C1913 a_n100_n52699# w_n358_n337587# 0.269531f
C1914 a_n100_329521# w_n358_n337587# 0.269531f
C1915 a_n158_n113230# w_n358_n337587# 0.689103f
C1916 a_100_n289842# w_n358_n337587# 0.689103f
C1917 a_n158_182002# a_100_182002# 0.655843f
C1918 a_100_n47330# a_100_n44694# 0.010536f
C1919 a_n158_160914# a_n158_158278# 0.010536f
C1920 a_n158_155642# a_n100_155545# 0.26189f
C1921 a_n158_131918# w_n358_n337587# 0.689103f
C1922 a_100_n2518# w_n358_n337587# 0.689103f
C1923 a_100_245266# a_100_247902# 0.010536f
C1924 a_n100_n210859# a_n100_n213495# 0.205388f
C1925 a_n100_313705# a_n100_311069# 0.205388f
C1926 a_100_292714# w_n358_n337587# 0.689103f
C1927 a_100_52838# w_n358_n337587# 0.689103f
C1928 a_100_n105322# a_n158_n105322# 0.655843f
C1929 a_n100_n329479# a_100_n329382# 0.26189f
C1930 a_100_316438# a_n100_316341# 0.26189f
C1931 a_n158_n150134# a_n158_n152770# 0.010536f
C1932 a_n158_n202854# w_n358_n337587# 0.689103f
C1933 a_n158_129282# a_100_129282# 0.655843f
C1934 a_100_134554# a_100_137190# 0.010536f
C1935 a_100_34386# a_100_31750# 0.010536f
C1936 a_n100_31653# a_n158_31750# 0.26189f
C1937 a_n158_208362# w_n358_n337587# 0.689103f
C1938 a_n100_n42155# a_n100_n44791# 0.205388f
C1939 w_n358_n337587# a_100_n308294# 0.689103f
C1940 a_n100_n250399# w_n358_n337587# 0.269531f
C1941 a_n158_n318838# a_n158_n321474# 0.010536f
C1942 a_100_8026# a_n100_7929# 0.26189f
C1943 a_n100_295253# a_n100_297889# 0.205388f
C1944 a_n100_300525# a_n158_300622# 0.26189f
C1945 w_n358_n337587# a_n158_n297750# 0.689103f
C1946 a_100_n237122# w_n358_n337587# 0.689103f
C1947 a_100_324346# a_n100_324249# 0.26189f
C1948 a_n158_n13062# a_100_n13062# 0.655843f
C1949 a_100_210998# a_100_213634# 0.010536f
C1950 a_100_n334654# a_100_n337290# 0.010536f
C1951 a_n100_n337387# a_n158_n337290# 0.26189f
C1952 a_100_n187038# w_n358_n337587# 0.689103f
C1953 a_100_n237122# a_100_n239758# 0.010536f
C1954 a_n100_305797# a_n100_303161# 0.205388f
C1955 a_n158_n218670# a_n158_n221306# 0.010536f
C1956 a_n158_n100050# a_n100_n100147# 0.26189f
C1957 a_100_197818# a_100_200454# 0.010536f
C1958 a_n158_n200218# w_n358_n337587# 0.689103f
C1959 a_n100_n100147# a_100_n100050# 0.26189f
C1960 a_100_126646# a_100_129282# 0.010536f
C1961 a_n100_n100147# w_n358_n337587# 0.269531f
C1962 a_100_n231850# w_n358_n337587# 0.689103f
C1963 a_100_n252938# a_100_n255574# 0.010536f
C1964 a_n100_n271487# a_n100_n274123# 0.205388f
C1965 a_100_332254# a_100_334890# 0.010536f
C1966 a_n158_n134318# a_n100_n134415# 0.26189f
C1967 a_100_n26242# a_n100_n26339# 0.26189f
C1968 a_n158_224178# a_100_224178# 0.655843f
C1969 a_100_290078# a_n100_289981# 0.26189f
C1970 a_n100_292617# a_n158_292714# 0.26189f
C1971 w_n358_n337587# a_n158_n332018# 0.689103f
C1972 a_n100_139729# w_n358_n337587# 0.269531f
C1973 a_100_5390# a_n100_5293# 0.26189f
C1974 a_n158_n65782# w_n358_n337587# 0.689103f
C1975 a_n100_n239855# a_n158_n239758# 0.26189f
C1976 a_n100_81737# a_n158_81834# 0.26189f
C1977 a_100_n71054# a_100_n68418# 0.010536f
C1978 a_n158_297986# w_n358_n337587# 0.689103f
C1979 a_n158_8026# w_n358_n337587# 0.689103f
C1980 a_n158_134554# a_n158_137190# 0.010536f
C1981 a_n158_n210762# a_n158_n208126# 0.010536f
C1982 a_n100_139729# a_n100_137093# 0.205388f
C1983 a_n158_n260846# w_n358_n337587# 0.689103f
C1984 a_n158_n303022# a_n158_n300386# 0.010536f
C1985 a_n100_n189771# a_n100_n187135# 0.205388f
C1986 a_n158_105558# a_n158_102922# 0.010536f
C1987 a_100_n181766# a_n100_n181863# 0.26189f
C1988 a_n100_229353# a_n100_231989# 0.205388f
C1989 a_n100_n79059# w_n358_n337587# 0.269531f
C1990 a_100_263718# w_n358_n337587# 0.689103f
C1991 a_n158_29114# w_n358_n337587# 0.689103f
C1992 a_n158_n160678# a_n158_n163314# 0.010536f
C1993 a_n100_n121235# a_n100_n123871# 0.205388f
C1994 a_n158_n28878# w_n358_n337587# 0.689103f
C1995 a_100_160914# w_n358_n337587# 0.689103f
C1996 a_n100_195085# a_n158_195182# 0.26189f
C1997 a_n100_n313663# a_n100_n311027# 0.205388f
C1998 a_100_n52602# a_100_n55238# 0.010536f
C1999 a_n100_13201# a_n158_13298# 0.26189f
C2000 a_n158_n242394# a_n158_n239758# 0.010536f
C2001 a_100_n49966# w_n358_n337587# 0.689103f
C2002 a_n158_324346# a_n158_326982# 0.010536f
C2003 a_n100_329521# a_n100_326885# 0.205388f
C2004 a_n100_n163411# a_n100_n166047# 0.205388f
C2005 a_n100_79101# w_n358_n337587# 0.269531f
C2006 a_n158_n2518# a_n100_n2615# 0.26189f
C2007 a_100_n131682# w_n358_n337587# 0.689103f
C2008 a_100_239994# w_n358_n337587# 0.689103f
C2009 a_n158_n86870# a_n158_n89506# 0.010536f
C2010 a_n100_173997# a_n100_176633# 0.205388f
C2011 a_n100_245169# a_n158_245266# 0.26189f
C2012 a_n158_73926# a_100_73926# 0.655843f
C2013 a_n100_73829# a_n100_71193# 0.205388f
C2014 a_n100_282073# w_n358_n337587# 0.269531f
C2015 a_n158_n139590# a_n158_n142226# 0.010536f
C2016 a_n158_118# a_n100_21# 0.26189f
C2017 a_n158_197818# a_n158_200454# 0.010536f
C2018 a_100_n255574# w_n358_n337587# 0.689103f
C2019 a_n100_n295211# a_n158_n295114# 0.26189f
C2020 a_100_n168586# w_n358_n337587# 0.689103f
C2021 a_100_n276662# a_100_n279298# 0.010536f
C2022 a_n100_n34247# a_100_n34150# 0.26189f
C2023 a_100_n205490# w_n358_n337587# 0.689103f
C2024 a_n100_253077# w_n358_n337587# 0.269531f
C2025 a_n158_n276662# a_100_n276662# 0.655843f
C2026 a_100_153006# a_100_150370# 0.010536f
C2027 a_n100_n60607# w_n358_n337587# 0.269531f
C2028 a_100_15934# w_n358_n337587# 0.689103f
C2029 a_100_n139590# a_100_n142226# 0.010536f
C2030 a_100_142462# w_n358_n337587# 0.689103f
C2031 a_100_n144862# w_n358_n337587# 0.689103f
C2032 a_100_118738# a_100_116102# 0.010536f
C2033 a_n100_171361# w_n358_n337587# 0.269531f
C2034 a_100_324346# a_n158_324346# 0.655843f
C2035 a_100_n13062# w_n358_n337587# 0.689103f
C2036 a_n158_n229214# a_n158_n226578# 0.010536f
C2037 a_n158_224178# w_n358_n337587# 0.689103f
C2038 a_n100_39561# a_n100_42197# 0.205388f
C2039 a_n100_36925# a_n158_37022# 0.26189f
C2040 a_n100_n158139# w_n358_n337587# 0.269531f
C2041 a_n100_n137051# a_n158_n136954# 0.26189f
C2042 a_100_n139590# a_100_n136954# 0.010536f
C2043 a_n158_42294# w_n358_n337587# 0.689103f
C2044 a_n158_268990# w_n358_n337587# 0.689103f
C2045 a_n158_68654# a_n158_66018# 0.010536f
C2046 a_n100_195085# w_n358_n337587# 0.269531f
C2047 a_n100_258349# a_n100_260985# 0.205388f
C2048 a_n100_n202951# w_n358_n337587# 0.269531f
C2049 a_n100_n318935# a_100_n318838# 0.26189f
C2050 w_n358_n337587# a_100_n305658# 0.689103f
C2051 a_100_n89506# a_n100_n89603# 0.26189f
C2052 a_n100_n216131# a_n100_n213495# 0.205388f
C2053 a_n100_87009# w_n358_n337587# 0.269531f
C2054 a_n158_n266118# w_n358_n337587# 0.689103f
C2055 a_n158_n326746# a_100_n326746# 0.655843f
C2056 a_n100_n326843# a_n100_n329479# 0.205388f
C2057 a_n100_245169# w_n358_n337587# 0.269531f
C2058 a_n100_55377# a_n158_55474# 0.26189f
C2059 a_100_n65782# a_100_n63146# 0.010536f
C2060 a_n158_n292478# a_100_n292478# 0.655843f
C2061 a_100_160914# a_100_158278# 0.010536f
C2062 a_n158_76562# a_n158_79198# 0.010536f
C2063 a_n158_290078# w_n358_n337587# 0.689103f
C2064 a_n100_313705# a_n100_316341# 0.205388f
C2065 a_100_n247666# a_100_n245030# 0.010536f
C2066 a_n100_n147595# a_n158_n147498# 0.26189f
C2067 a_100_n250302# a_n100_n250399# 0.26189f
C2068 a_n100_n84331# a_100_n84234# 0.26189f
C2069 a_100_n102686# a_100_n100050# 0.010536f
C2070 a_n158_n84234# a_n100_n84331# 0.26189f
C2071 a_100_26478# w_n358_n337587# 0.689103f
C2072 a_100_n102686# w_n358_n337587# 0.689103f
C2073 a_100_274262# a_100_271626# 0.010536f
C2074 a_n100_271529# a_n158_271626# 0.26189f
C2075 a_n100_31653# a_100_31750# 0.26189f
C2076 a_n158_n163314# w_n358_n337587# 0.689103f
C2077 a_100_102922# w_n358_n337587# 0.689103f
C2078 a_100_n274026# w_n358_n337587# 0.689103f
C2079 a_n100_n326843# a_n158_n326746# 0.26189f
C2080 a_100_21206# a_100_23842# 0.010536f
C2081 w_n358_n337587# a_100_n295114# 0.689103f
C2082 a_n158_n281934# w_n358_n337587# 0.689103f
C2083 a_n100_300525# a_100_300622# 0.26189f
C2084 a_n100_n266215# w_n358_n337587# 0.269531f
C2085 a_n100_n129143# w_n358_n337587# 0.269531f
C2086 a_100_n142226# w_n358_n337587# 0.689103f
C2087 a_100_n279298# a_n100_n279395# 0.26189f
C2088 a_n158_n144862# a_n158_n142226# 0.010536f
C2089 a_n158_n63146# a_100_n63146# 0.655843f
C2090 a_n158_313802# w_n358_n337587# 0.689103f
C2091 a_100_92378# a_100_89742# 0.010536f
C2092 a_n100_n187135# a_n100_n184499# 0.205388f
C2093 w_n358_n337587# a_n158_n329382# 0.689103f
C2094 a_n100_279437# a_n100_282073# 0.205388f
C2095 a_n100_n86967# a_n158_n86870# 0.26189f
C2096 a_n158_n84234# a_100_n84234# 0.655843f
C2097 a_n158_232086# w_n358_n337587# 0.689103f
C2098 a_n100_n152867# w_n358_n337587# 0.269531f
C2099 a_n100_n308391# a_n100_n305755# 0.205388f
C2100 a_n100_n176591# a_n100_n173955# 0.205388f
C2101 a_n100_110733# a_n158_110830# 0.26189f
C2102 a_100_50202# w_n358_n337587# 0.689103f
C2103 a_n158_282170# w_n358_n337587# 0.689103f
C2104 a_100_n136954# w_n358_n337587# 0.689103f
C2105 a_100_197818# a_n100_197721# 0.26189f
C2106 a_100_n300386# a_n100_n300483# 0.26189f
C2107 a_n100_n52699# a_n100_n50063# 0.205388f
C2108 a_n158_261082# a_n100_260985# 0.26189f
C2109 a_100_n76326# w_n358_n337587# 0.689103f
C2110 a_n100_n134415# w_n358_n337587# 0.269531f
C2111 a_n158_n216034# a_n158_n218670# 0.010536f
C2112 a_100_97650# a_100_95014# 0.010536f
C2113 a_n100_94917# a_n158_95014# 0.26189f
C2114 a_n100_94917# w_n358_n337587# 0.269531f
C2115 a_100_332254# a_n158_332254# 0.655843f
C2116 a_n100_n94875# w_n358_n337587# 0.269531f
C2117 a_n158_224178# a_n158_221542# 0.010536f
C2118 a_n158_n31514# a_n158_n28878# 0.010536f
C2119 a_n158_n134318# w_n358_n337587# 0.689103f
C2120 a_n100_52741# a_100_52838# 0.26189f
C2121 a_n158_n49966# w_n358_n337587# 0.689103f
C2122 a_100_139826# w_n358_n337587# 0.689103f
C2123 a_n100_163453# w_n358_n337587# 0.269531f
C2124 a_n158_n39422# w_n358_n337587# 0.689103f
C2125 a_n100_n300483# a_n158_n300386# 0.26189f
C2126 a_100_247902# a_n100_247805# 0.26189f
C2127 a_n100_n21067# a_n100_n18431# 0.205388f
C2128 a_100_316438# a_100_319074# 0.010536f
C2129 a_n158_303258# w_n358_n337587# 0.689103f
C2130 a_100_84470# a_100_81834# 0.010536f
C2131 a_n100_n89603# w_n358_n337587# 0.269531f
C2132 a_100_n229214# w_n358_n337587# 0.689103f
C2133 a_n158_216270# w_n358_n337587# 0.689103f
C2134 a_100_n65782# a_n158_n65782# 0.655843f
C2135 a_100_274262# a_100_276898# 0.010536f
C2136 a_n100_163453# a_n158_163550# 0.26189f
C2137 a_n158_n181766# w_n358_n337587# 0.689103f
C2138 a_n158_n92142# a_n158_n89506# 0.010536f
C2139 a_n100_n197679# a_n100_n195043# 0.205388f
C2140 a_n100_n42155# a_100_n42058# 0.26189f
C2141 a_n100_260985# w_n358_n337587# 0.269531f
C2142 a_100_n231850# a_n158_n231850# 0.655843f
C2143 a_n100_150273# w_n358_n337587# 0.269531f
C2144 a_n100_n316299# a_100_n316202# 0.26189f
C2145 a_n158_n237122# a_n158_n239758# 0.010536f
C2146 a_100_n194946# w_n358_n337587# 0.689103f
C2147 a_n100_255713# a_n158_255810# 0.26189f
C2148 a_100_n60510# a_100_n57874# 0.010536f
C2149 a_n100_187177# w_n358_n337587# 0.269531f
C2150 a_n158_79198# w_n358_n337587# 0.689103f
C2151 a_100_321710# w_n358_n337587# 0.689103f
C2152 a_100_218906# a_n158_218906# 0.655843f
C2153 a_n100_n102783# a_n100_n105419# 0.205388f
C2154 a_n100_145001# a_n100_147637# 0.205388f
C2155 a_n100_284709# a_100_284806# 0.26189f
C2156 a_100_47566# a_100_44930# 0.010536f
C2157 a_n100_n84331# w_n358_n337587# 0.269531f
C2158 a_n158_47566# a_n158_50202# 0.010536f
C2159 a_n100_245169# a_100_245266# 0.26189f
C2160 a_100_118# w_n358_n337587# 0.689103f
C2161 a_n158_n281934# a_n158_n279298# 0.010536f
C2162 a_n158_316438# a_100_316438# 0.655843f
C2163 a_100_76562# a_100_79198# 0.010536f
C2164 a_n158_n63146# a_n158_n65782# 0.010536f
C2165 a_n158_n187038# w_n358_n337587# 0.689103f
C2166 a_100_n160678# a_n100_n160775# 0.26189f
C2167 a_n158_n13062# w_n358_n337587# 0.689103f
C2168 a_n100_n26339# a_n100_n23703# 0.205388f
C2169 a_100_n131682# a_100_n129046# 0.010536f
C2170 a_n158_n284570# a_n100_n284667# 0.26189f
C2171 a_n100_224081# a_n100_226717# 0.205388f
C2172 a_n158_n250302# w_n358_n337587# 0.689103f
C2173 a_n100_n263579# a_n100_n266215# 0.205388f
C2174 a_100_n213398# a_100_n216034# 0.010536f
C2175 a_n100_258349# w_n358_n337587# 0.269531f
C2176 a_n100_150273# a_n158_150370# 0.26189f
C2177 a_100_189910# a_100_187274# 0.010536f
C2178 a_100_n84234# w_n358_n337587# 0.689103f
C2179 a_n158_n55238# a_100_n55238# 0.655843f
C2180 a_n158_n160678# w_n358_n337587# 0.689103f
C2181 a_n158_n110594# w_n358_n337587# 0.689103f
C2182 a_n158_n84234# w_n358_n337587# 0.689103f
C2183 a_n158_84470# a_n158_87106# 0.010536f
C2184 a_n158_76562# w_n358_n337587# 0.689103f
C2185 a_n100_208265# a_n100_210901# 0.205388f
C2186 a_100_n332018# a_100_n334654# 0.010536f
C2187 a_n100_n334751# a_n158_n334654# 0.26189f
C2188 a_100_n271390# a_100_n268754# 0.010536f
C2189 a_100_n89506# w_n358_n337587# 0.689103f
C2190 a_n100_158181# w_n358_n337587# 0.269531f
C2191 a_n158_n47330# a_100_n47330# 0.655843f
C2192 a_100_224178# w_n358_n337587# 0.689103f
C2193 a_100_n289842# a_100_n287206# 0.010536f
C2194 a_100_279534# a_100_276898# 0.010536f
C2195 a_n100_276801# a_n158_276898# 0.26189f
C2196 a_100_n123774# w_n358_n337587# 0.689103f
C2197 a_n100_173997# a_n158_174094# 0.26189f
C2198 a_n158_n5154# a_100_n5154# 0.655843f
C2199 a_n100_168725# a_n100_171361# 0.205388f
C2200 a_n158_168822# a_n158_171458# 0.010536f
C2201 a_100_n213398# w_n358_n337587# 0.689103f
C2202 a_100_n84234# a_100_n86870# 0.010536f
C2203 a_n100_274165# w_n358_n337587# 0.269531f
C2204 a_n100_n176591# a_100_n176494# 0.26189f
C2205 a_n158_68654# a_n158_71290# 0.010536f
C2206 a_n158_303258# a_n100_303161# 0.26189f
C2207 a_n100_n50063# a_100_n49966# 0.26189f
C2208 a_n100_n65879# a_n100_n63243# 0.205388f
C2209 a_n100_n221403# w_n358_n337587# 0.269531f
C2210 a_n158_195182# w_n358_n337587# 0.689103f
C2211 a_n158_n189674# a_100_n189674# 0.655843f
C2212 a_100_n31514# w_n358_n337587# 0.689103f
C2213 a_100_n247666# a_n100_n247763# 0.26189f
C2214 w_n358_n337587# a_n158_n316202# 0.689103f
C2215 a_100_n7790# w_n358_n337587# 0.689103f
C2216 a_100_n139590# w_n358_n337587# 0.689103f
C2217 a_n100_329521# a_n100_332157# 0.205388f
C2218 a_n100_n79059# a_n158_n78962# 0.26189f
C2219 a_n158_329618# w_n358_n337587# 0.689103f
C2220 a_100_n89506# a_100_n86870# 0.010536f
C2221 a_n158_245266# w_n358_n337587# 0.689103f
C2222 a_100_n5154# a_100_n2518# 0.010536f
C2223 a_n100_55377# a_100_55474# 0.26189f
C2224 a_n100_7929# a_n100_5293# 0.205388f
C2225 a_100_n252938# w_n358_n337587# 0.689103f
C2226 a_n100_n139687# a_100_n139590# 0.26189f
C2227 a_n158_108194# a_100_108194# 0.655843f
C2228 a_n158_n126410# w_n358_n337587# 0.689103f
C2229 a_n100_n5251# w_n358_n337587# 0.269531f
C2230 a_n158_153006# a_n158_155642# 0.010536f
C2231 a_n158_313802# a_n158_311166# 0.010536f
C2232 a_n158_63382# w_n358_n337587# 0.689103f
C2233 a_n100_n242491# a_n100_n239855# 0.205388f
C2234 a_n158_n57874# w_n358_n337587# 0.689103f
C2235 a_n100_202993# a_n100_205629# 0.205388f
C2236 a_100_n245030# a_100_n242394# 0.010536f
C2237 a_100_n23606# w_n358_n337587# 0.689103f
C2238 a_n100_23745# w_n358_n337587# 0.269531f
C2239 a_n100_n166047# a_100_n165950# 0.26189f
C2240 a_n100_271529# a_100_271626# 0.26189f
C2241 a_n158_274262# a_n100_274165# 0.26189f
C2242 a_n158_100286# w_n358_n337587# 0.689103f
C2243 a_100_n76326# a_n158_n76326# 0.655843f
C2244 a_n158_n289842# a_n158_n287206# 0.010536f
C2245 w_n358_n337587# a_100_n324110# 0.689103f
C2246 a_n100_15837# a_100_15934# 0.26189f
C2247 a_100_63382# a_n100_63285# 0.26189f
C2248 a_n158_60746# a_n158_58110# 0.010536f
C2249 a_n158_261082# w_n358_n337587# 0.689103f
C2250 a_n100_258349# a_n158_258446# 0.26189f
C2251 a_n100_n242491# a_n158_n242394# 0.26189f
C2252 a_100_n18334# w_n358_n337587# 0.689103f
C2253 a_n158_n155406# a_100_n155406# 0.655843f
C2254 a_100_n216034# w_n358_n337587# 0.689103f
C2255 a_n158_171458# a_100_171458# 0.655843f
C2256 a_100_n118502# w_n358_n337587# 0.689103f
C2257 a_100_121374# w_n358_n337587# 0.689103f
C2258 a_100_n160678# a_100_n158042# 0.010536f
C2259 a_n100_n129143# a_100_n129046# 0.26189f
C2260 a_100_n173858# w_n358_n337587# 0.689103f
C2261 a_n158_237358# a_n158_239994# 0.010536f
C2262 a_100_n97414# a_100_n100050# 0.010536f
C2263 a_n100_234625# a_n158_234722# 0.26189f
C2264 a_n100_47469# w_n358_n337587# 0.269531f
C2265 a_n158_71290# a_n158_73926# 0.010536f
C2266 a_n100_76465# a_100_76562# 0.26189f
C2267 a_n158_n100050# a_100_n100050# 0.655843f
C2268 a_n100_287345# w_n358_n337587# 0.269531f
C2269 a_n100_195085# a_n100_197721# 0.205388f
C2270 a_n158_n100050# w_n358_n337587# 0.689103f
C2271 a_100_n97414# w_n358_n337587# 0.689103f
C2272 a_n100_158181# a_100_158278# 0.26189f
C2273 a_100_n100050# w_n358_n337587# 0.689103f
C2274 a_n158_95014# w_n358_n337587# 0.689103f
C2275 a_n158_n7790# a_n158_n10426# 0.010536f
C2276 a_n158_n313566# a_n158_n316202# 0.010536f
C2277 a_100_55474# a_100_58110# 0.010536f
C2278 a_n100_292617# a_100_292714# 0.26189f
C2279 a_n100_137093# w_n358_n337587# 0.269531f
C2280 a_n100_118641# a_n100_116005# 0.205388f
C2281 a_100_n245030# a_n100_n245127# 0.26189f
C2282 a_n158_n213398# a_n158_n210762# 0.010536f
C2283 a_100_n52602# a_n158_n52602# 0.655843f
C2284 a_n100_n139687# w_n358_n337587# 0.269531f
C2285 a_100_253174# a_100_250538# 0.010536f
C2286 a_n158_163550# w_n358_n337587# 0.689103f
C2287 a_n100_n105419# a_n100_n108055# 0.205388f
C2288 a_n100_81737# a_100_81834# 0.26189f
C2289 a_n158_84470# a_n100_84373# 0.26189f
C2290 a_100_71290# w_n358_n337587# 0.689103f
C2291 a_100_n239758# w_n358_n337587# 0.689103f
C2292 a_n158_210998# a_n158_208362# 0.010536f
C2293 a_100_205726# a_100_208362# 0.010536f
C2294 a_n158_139826# a_n158_137190# 0.010536f
C2295 a_n100_213537# w_n358_n337587# 0.269531f
C2296 a_100_37022# a_n100_36925# 0.26189f
C2297 a_100_n86870# w_n358_n337587# 0.689103f
C2298 a_n100_n47427# w_n358_n337587# 0.269531f
C2299 a_n100_n115963# w_n358_n337587# 0.269531f
C2300 a_n100_102825# a_n158_102922# 0.26189f
C2301 a_100_n337290# VSUBS 0.58217f
C2302 a_n158_n337290# VSUBS 0.58217f
C2303 a_n100_n337387# VSUBS 0.291162f
C2304 a_100_n334654# VSUBS 0.576721f
C2305 a_n158_n334654# VSUBS 0.576721f
C2306 a_n100_n334751# VSUBS 0.247431f
C2307 a_100_n332018# VSUBS 0.576721f
C2308 a_n158_n332018# VSUBS 0.576721f
C2309 a_n100_n332115# VSUBS 0.247431f
C2310 a_100_n329382# VSUBS 0.576721f
C2311 a_n158_n329382# VSUBS 0.576721f
C2312 a_n100_n329479# VSUBS 0.247431f
C2313 a_100_n326746# VSUBS 0.576721f
C2314 a_n158_n326746# VSUBS 0.576721f
C2315 a_n100_n326843# VSUBS 0.247431f
C2316 a_100_n324110# VSUBS 0.576721f
C2317 a_n158_n324110# VSUBS 0.576721f
C2318 a_n100_n324207# VSUBS 0.247431f
C2319 a_100_n321474# VSUBS 0.576721f
C2320 a_n158_n321474# VSUBS 0.576721f
C2321 a_n100_n321571# VSUBS 0.247431f
C2322 a_100_n318838# VSUBS 0.576721f
C2323 a_n158_n318838# VSUBS 0.576721f
C2324 a_n100_n318935# VSUBS 0.247431f
C2325 a_100_n316202# VSUBS 0.576721f
C2326 a_n158_n316202# VSUBS 0.576721f
C2327 a_n100_n316299# VSUBS 0.247431f
C2328 a_100_n313566# VSUBS 0.576721f
C2329 a_n158_n313566# VSUBS 0.576721f
C2330 a_n100_n313663# VSUBS 0.247431f
C2331 a_100_n310930# VSUBS 0.576721f
C2332 a_n158_n310930# VSUBS 0.576721f
C2333 a_n100_n311027# VSUBS 0.247431f
C2334 a_100_n308294# VSUBS 0.576721f
C2335 a_n158_n308294# VSUBS 0.576721f
C2336 a_n100_n308391# VSUBS 0.247431f
C2337 a_100_n305658# VSUBS 0.576721f
C2338 a_n158_n305658# VSUBS 0.576721f
C2339 a_n100_n305755# VSUBS 0.247431f
C2340 a_100_n303022# VSUBS 0.576721f
C2341 a_n158_n303022# VSUBS 0.576721f
C2342 a_n100_n303119# VSUBS 0.247431f
C2343 a_100_n300386# VSUBS 0.576721f
C2344 a_n158_n300386# VSUBS 0.576721f
C2345 a_n100_n300483# VSUBS 0.247431f
C2346 a_100_n297750# VSUBS 0.576721f
C2347 a_n158_n297750# VSUBS 0.576721f
C2348 a_n100_n297847# VSUBS 0.247431f
C2349 a_100_n295114# VSUBS 0.576721f
C2350 a_n158_n295114# VSUBS 0.576721f
C2351 a_n100_n295211# VSUBS 0.247431f
C2352 a_100_n292478# VSUBS 0.576721f
C2353 a_n158_n292478# VSUBS 0.576721f
C2354 a_n100_n292575# VSUBS 0.247431f
C2355 a_100_n289842# VSUBS 0.576721f
C2356 a_n158_n289842# VSUBS 0.576721f
C2357 a_n100_n289939# VSUBS 0.247431f
C2358 a_100_n287206# VSUBS 0.576721f
C2359 a_n158_n287206# VSUBS 0.576721f
C2360 a_n100_n287303# VSUBS 0.247431f
C2361 a_100_n284570# VSUBS 0.576721f
C2362 a_n158_n284570# VSUBS 0.576721f
C2363 a_n100_n284667# VSUBS 0.247431f
C2364 a_100_n281934# VSUBS 0.576721f
C2365 a_n158_n281934# VSUBS 0.576721f
C2366 a_n100_n282031# VSUBS 0.247431f
C2367 a_100_n279298# VSUBS 0.576721f
C2368 a_n158_n279298# VSUBS 0.576721f
C2369 a_n100_n279395# VSUBS 0.247431f
C2370 a_100_n276662# VSUBS 0.576721f
C2371 a_n158_n276662# VSUBS 0.576721f
C2372 a_n100_n276759# VSUBS 0.247431f
C2373 a_100_n274026# VSUBS 0.576721f
C2374 a_n158_n274026# VSUBS 0.576721f
C2375 a_n100_n274123# VSUBS 0.247431f
C2376 a_100_n271390# VSUBS 0.576721f
C2377 a_n158_n271390# VSUBS 0.576721f
C2378 a_n100_n271487# VSUBS 0.247431f
C2379 a_100_n268754# VSUBS 0.576721f
C2380 a_n158_n268754# VSUBS 0.576721f
C2381 a_n100_n268851# VSUBS 0.247431f
C2382 a_100_n266118# VSUBS 0.576721f
C2383 a_n158_n266118# VSUBS 0.576721f
C2384 a_n100_n266215# VSUBS 0.247431f
C2385 a_100_n263482# VSUBS 0.576721f
C2386 a_n158_n263482# VSUBS 0.576721f
C2387 a_n100_n263579# VSUBS 0.247431f
C2388 a_100_n260846# VSUBS 0.576721f
C2389 a_n158_n260846# VSUBS 0.576721f
C2390 a_n100_n260943# VSUBS 0.247431f
C2391 a_100_n258210# VSUBS 0.576721f
C2392 a_n158_n258210# VSUBS 0.576721f
C2393 a_n100_n258307# VSUBS 0.247431f
C2394 a_100_n255574# VSUBS 0.576721f
C2395 a_n158_n255574# VSUBS 0.576721f
C2396 a_n100_n255671# VSUBS 0.247431f
C2397 a_100_n252938# VSUBS 0.576721f
C2398 a_n158_n252938# VSUBS 0.576721f
C2399 a_n100_n253035# VSUBS 0.247431f
C2400 a_100_n250302# VSUBS 0.576721f
C2401 a_n158_n250302# VSUBS 0.576721f
C2402 a_n100_n250399# VSUBS 0.247431f
C2403 a_100_n247666# VSUBS 0.576721f
C2404 a_n158_n247666# VSUBS 0.576721f
C2405 a_n100_n247763# VSUBS 0.247431f
C2406 a_100_n245030# VSUBS 0.576721f
C2407 a_n158_n245030# VSUBS 0.576721f
C2408 a_n100_n245127# VSUBS 0.247431f
C2409 a_100_n242394# VSUBS 0.576721f
C2410 a_n158_n242394# VSUBS 0.576721f
C2411 a_n100_n242491# VSUBS 0.247431f
C2412 a_100_n239758# VSUBS 0.576721f
C2413 a_n158_n239758# VSUBS 0.576721f
C2414 a_n100_n239855# VSUBS 0.247431f
C2415 a_100_n237122# VSUBS 0.576721f
C2416 a_n158_n237122# VSUBS 0.576721f
C2417 a_n100_n237219# VSUBS 0.247431f
C2418 a_100_n234486# VSUBS 0.576721f
C2419 a_n158_n234486# VSUBS 0.576721f
C2420 a_n100_n234583# VSUBS 0.247431f
C2421 a_100_n231850# VSUBS 0.576721f
C2422 a_n158_n231850# VSUBS 0.576721f
C2423 a_n100_n231947# VSUBS 0.247431f
C2424 a_100_n229214# VSUBS 0.576721f
C2425 a_n158_n229214# VSUBS 0.576721f
C2426 a_n100_n229311# VSUBS 0.247431f
C2427 a_100_n226578# VSUBS 0.576721f
C2428 a_n158_n226578# VSUBS 0.576721f
C2429 a_n100_n226675# VSUBS 0.247431f
C2430 a_100_n223942# VSUBS 0.576721f
C2431 a_n158_n223942# VSUBS 0.576721f
C2432 a_n100_n224039# VSUBS 0.247431f
C2433 a_100_n221306# VSUBS 0.576721f
C2434 a_n158_n221306# VSUBS 0.576721f
C2435 a_n100_n221403# VSUBS 0.247431f
C2436 a_100_n218670# VSUBS 0.576721f
C2437 a_n158_n218670# VSUBS 0.576721f
C2438 a_n100_n218767# VSUBS 0.247431f
C2439 a_100_n216034# VSUBS 0.576721f
C2440 a_n158_n216034# VSUBS 0.576721f
C2441 a_n100_n216131# VSUBS 0.247431f
C2442 a_100_n213398# VSUBS 0.576721f
C2443 a_n158_n213398# VSUBS 0.576721f
C2444 a_n100_n213495# VSUBS 0.247431f
C2445 a_100_n210762# VSUBS 0.576721f
C2446 a_n158_n210762# VSUBS 0.576721f
C2447 a_n100_n210859# VSUBS 0.247431f
C2448 a_100_n208126# VSUBS 0.576721f
C2449 a_n158_n208126# VSUBS 0.576721f
C2450 a_n100_n208223# VSUBS 0.247431f
C2451 a_100_n205490# VSUBS 0.576721f
C2452 a_n158_n205490# VSUBS 0.576721f
C2453 a_n100_n205587# VSUBS 0.247431f
C2454 a_100_n202854# VSUBS 0.576721f
C2455 a_n158_n202854# VSUBS 0.576721f
C2456 a_n100_n202951# VSUBS 0.247431f
C2457 a_100_n200218# VSUBS 0.576721f
C2458 a_n158_n200218# VSUBS 0.576721f
C2459 a_n100_n200315# VSUBS 0.247431f
C2460 a_100_n197582# VSUBS 0.576721f
C2461 a_n158_n197582# VSUBS 0.576721f
C2462 a_n100_n197679# VSUBS 0.247431f
C2463 a_100_n194946# VSUBS 0.576721f
C2464 a_n158_n194946# VSUBS 0.576721f
C2465 a_n100_n195043# VSUBS 0.247431f
C2466 a_100_n192310# VSUBS 0.576721f
C2467 a_n158_n192310# VSUBS 0.576721f
C2468 a_n100_n192407# VSUBS 0.247431f
C2469 a_100_n189674# VSUBS 0.576721f
C2470 a_n158_n189674# VSUBS 0.576721f
C2471 a_n100_n189771# VSUBS 0.247431f
C2472 a_100_n187038# VSUBS 0.576721f
C2473 a_n158_n187038# VSUBS 0.576721f
C2474 a_n100_n187135# VSUBS 0.247431f
C2475 a_100_n184402# VSUBS 0.576721f
C2476 a_n158_n184402# VSUBS 0.576721f
C2477 a_n100_n184499# VSUBS 0.247431f
C2478 a_100_n181766# VSUBS 0.576721f
C2479 a_n158_n181766# VSUBS 0.576721f
C2480 a_n100_n181863# VSUBS 0.247431f
C2481 a_100_n179130# VSUBS 0.576721f
C2482 a_n158_n179130# VSUBS 0.576721f
C2483 a_n100_n179227# VSUBS 0.247431f
C2484 a_100_n176494# VSUBS 0.576721f
C2485 a_n158_n176494# VSUBS 0.576721f
C2486 a_n100_n176591# VSUBS 0.247431f
C2487 a_100_n173858# VSUBS 0.576721f
C2488 a_n158_n173858# VSUBS 0.576721f
C2489 a_n100_n173955# VSUBS 0.247431f
C2490 a_100_n171222# VSUBS 0.576721f
C2491 a_n158_n171222# VSUBS 0.576721f
C2492 a_n100_n171319# VSUBS 0.247431f
C2493 a_100_n168586# VSUBS 0.576721f
C2494 a_n158_n168586# VSUBS 0.576721f
C2495 a_n100_n168683# VSUBS 0.247431f
C2496 a_100_n165950# VSUBS 0.576721f
C2497 a_n158_n165950# VSUBS 0.576721f
C2498 a_n100_n166047# VSUBS 0.247431f
C2499 a_100_n163314# VSUBS 0.576721f
C2500 a_n158_n163314# VSUBS 0.576721f
C2501 a_n100_n163411# VSUBS 0.247431f
C2502 a_100_n160678# VSUBS 0.576721f
C2503 a_n158_n160678# VSUBS 0.576721f
C2504 a_n100_n160775# VSUBS 0.247431f
C2505 a_100_n158042# VSUBS 0.576721f
C2506 a_n158_n158042# VSUBS 0.576721f
C2507 a_n100_n158139# VSUBS 0.247431f
C2508 a_100_n155406# VSUBS 0.576721f
C2509 a_n158_n155406# VSUBS 0.576721f
C2510 a_n100_n155503# VSUBS 0.247431f
C2511 a_100_n152770# VSUBS 0.576721f
C2512 a_n158_n152770# VSUBS 0.576721f
C2513 a_n100_n152867# VSUBS 0.247431f
C2514 a_100_n150134# VSUBS 0.576721f
C2515 a_n158_n150134# VSUBS 0.576721f
C2516 a_n100_n150231# VSUBS 0.247431f
C2517 a_100_n147498# VSUBS 0.576721f
C2518 a_n158_n147498# VSUBS 0.576721f
C2519 a_n100_n147595# VSUBS 0.247431f
C2520 a_100_n144862# VSUBS 0.576721f
C2521 a_n158_n144862# VSUBS 0.576721f
C2522 a_n100_n144959# VSUBS 0.247431f
C2523 a_100_n142226# VSUBS 0.576721f
C2524 a_n158_n142226# VSUBS 0.576721f
C2525 a_n100_n142323# VSUBS 0.247431f
C2526 a_100_n139590# VSUBS 0.576721f
C2527 a_n158_n139590# VSUBS 0.576721f
C2528 a_n100_n139687# VSUBS 0.247431f
C2529 a_100_n136954# VSUBS 0.576721f
C2530 a_n158_n136954# VSUBS 0.576721f
C2531 a_n100_n137051# VSUBS 0.247431f
C2532 a_100_n134318# VSUBS 0.576721f
C2533 a_n158_n134318# VSUBS 0.576721f
C2534 a_n100_n134415# VSUBS 0.247431f
C2535 a_100_n131682# VSUBS 0.576721f
C2536 a_n158_n131682# VSUBS 0.576721f
C2537 a_n100_n131779# VSUBS 0.247431f
C2538 a_100_n129046# VSUBS 0.576721f
C2539 a_n158_n129046# VSUBS 0.576721f
C2540 a_n100_n129143# VSUBS 0.247431f
C2541 a_100_n126410# VSUBS 0.576721f
C2542 a_n158_n126410# VSUBS 0.576721f
C2543 a_n100_n126507# VSUBS 0.247431f
C2544 a_100_n123774# VSUBS 0.576721f
C2545 a_n158_n123774# VSUBS 0.576721f
C2546 a_n100_n123871# VSUBS 0.247431f
C2547 a_100_n121138# VSUBS 0.576721f
C2548 a_n158_n121138# VSUBS 0.576721f
C2549 a_n100_n121235# VSUBS 0.247431f
C2550 a_100_n118502# VSUBS 0.576721f
C2551 a_n158_n118502# VSUBS 0.576721f
C2552 a_n100_n118599# VSUBS 0.247431f
C2553 a_100_n115866# VSUBS 0.576721f
C2554 a_n158_n115866# VSUBS 0.576721f
C2555 a_n100_n115963# VSUBS 0.247431f
C2556 a_100_n113230# VSUBS 0.576721f
C2557 a_n158_n113230# VSUBS 0.576721f
C2558 a_n100_n113327# VSUBS 0.247431f
C2559 a_100_n110594# VSUBS 0.576721f
C2560 a_n158_n110594# VSUBS 0.576721f
C2561 a_n100_n110691# VSUBS 0.247431f
C2562 a_100_n107958# VSUBS 0.576721f
C2563 a_n158_n107958# VSUBS 0.576721f
C2564 a_n100_n108055# VSUBS 0.247431f
C2565 a_100_n105322# VSUBS 0.576721f
C2566 a_n158_n105322# VSUBS 0.576721f
C2567 a_n100_n105419# VSUBS 0.247431f
C2568 a_100_n102686# VSUBS 0.576721f
C2569 a_n158_n102686# VSUBS 0.576721f
C2570 a_n100_n102783# VSUBS 0.247431f
C2571 a_100_n100050# VSUBS 0.576721f
C2572 a_n158_n100050# VSUBS 0.576721f
C2573 a_n100_n100147# VSUBS 0.247431f
C2574 a_100_n97414# VSUBS 0.576721f
C2575 a_n158_n97414# VSUBS 0.576721f
C2576 a_n100_n97511# VSUBS 0.247431f
C2577 a_100_n94778# VSUBS 0.576721f
C2578 a_n158_n94778# VSUBS 0.576721f
C2579 a_n100_n94875# VSUBS 0.247431f
C2580 a_100_n92142# VSUBS 0.576721f
C2581 a_n158_n92142# VSUBS 0.576721f
C2582 a_n100_n92239# VSUBS 0.247431f
C2583 a_100_n89506# VSUBS 0.576721f
C2584 a_n158_n89506# VSUBS 0.576721f
C2585 a_n100_n89603# VSUBS 0.247431f
C2586 a_100_n86870# VSUBS 0.576721f
C2587 a_n158_n86870# VSUBS 0.576721f
C2588 a_n100_n86967# VSUBS 0.247431f
C2589 a_100_n84234# VSUBS 0.576721f
C2590 a_n158_n84234# VSUBS 0.576721f
C2591 a_n100_n84331# VSUBS 0.247431f
C2592 a_100_n81598# VSUBS 0.576721f
C2593 a_n158_n81598# VSUBS 0.576721f
C2594 a_n100_n81695# VSUBS 0.247431f
C2595 a_100_n78962# VSUBS 0.576721f
C2596 a_n158_n78962# VSUBS 0.576721f
C2597 a_n100_n79059# VSUBS 0.247431f
C2598 a_100_n76326# VSUBS 0.576721f
C2599 a_n158_n76326# VSUBS 0.576721f
C2600 a_n100_n76423# VSUBS 0.247431f
C2601 a_100_n73690# VSUBS 0.576721f
C2602 a_n158_n73690# VSUBS 0.576721f
C2603 a_n100_n73787# VSUBS 0.247431f
C2604 a_100_n71054# VSUBS 0.576721f
C2605 a_n158_n71054# VSUBS 0.576721f
C2606 a_n100_n71151# VSUBS 0.247431f
C2607 a_100_n68418# VSUBS 0.576721f
C2608 a_n158_n68418# VSUBS 0.576721f
C2609 a_n100_n68515# VSUBS 0.247431f
C2610 a_100_n65782# VSUBS 0.576721f
C2611 a_n158_n65782# VSUBS 0.576721f
C2612 a_n100_n65879# VSUBS 0.247431f
C2613 a_100_n63146# VSUBS 0.576721f
C2614 a_n158_n63146# VSUBS 0.576721f
C2615 a_n100_n63243# VSUBS 0.247431f
C2616 a_100_n60510# VSUBS 0.576721f
C2617 a_n158_n60510# VSUBS 0.576721f
C2618 a_n100_n60607# VSUBS 0.247431f
C2619 a_100_n57874# VSUBS 0.576721f
C2620 a_n158_n57874# VSUBS 0.576721f
C2621 a_n100_n57971# VSUBS 0.247431f
C2622 a_100_n55238# VSUBS 0.576721f
C2623 a_n158_n55238# VSUBS 0.576721f
C2624 a_n100_n55335# VSUBS 0.247431f
C2625 a_100_n52602# VSUBS 0.576721f
C2626 a_n158_n52602# VSUBS 0.576721f
C2627 a_n100_n52699# VSUBS 0.247431f
C2628 a_100_n49966# VSUBS 0.576721f
C2629 a_n158_n49966# VSUBS 0.576721f
C2630 a_n100_n50063# VSUBS 0.247431f
C2631 a_100_n47330# VSUBS 0.576721f
C2632 a_n158_n47330# VSUBS 0.576721f
C2633 a_n100_n47427# VSUBS 0.247431f
C2634 a_100_n44694# VSUBS 0.576721f
C2635 a_n158_n44694# VSUBS 0.576721f
C2636 a_n100_n44791# VSUBS 0.247431f
C2637 a_100_n42058# VSUBS 0.576721f
C2638 a_n158_n42058# VSUBS 0.576721f
C2639 a_n100_n42155# VSUBS 0.247431f
C2640 a_100_n39422# VSUBS 0.576721f
C2641 a_n158_n39422# VSUBS 0.576721f
C2642 a_n100_n39519# VSUBS 0.247431f
C2643 a_100_n36786# VSUBS 0.576721f
C2644 a_n158_n36786# VSUBS 0.576721f
C2645 a_n100_n36883# VSUBS 0.247431f
C2646 a_100_n34150# VSUBS 0.576721f
C2647 a_n158_n34150# VSUBS 0.576721f
C2648 a_n100_n34247# VSUBS 0.247431f
C2649 a_100_n31514# VSUBS 0.576721f
C2650 a_n158_n31514# VSUBS 0.576721f
C2651 a_n100_n31611# VSUBS 0.247431f
C2652 a_100_n28878# VSUBS 0.576721f
C2653 a_n158_n28878# VSUBS 0.576721f
C2654 a_n100_n28975# VSUBS 0.247431f
C2655 a_100_n26242# VSUBS 0.576721f
C2656 a_n158_n26242# VSUBS 0.576721f
C2657 a_n100_n26339# VSUBS 0.247431f
C2658 a_100_n23606# VSUBS 0.576721f
C2659 a_n158_n23606# VSUBS 0.576721f
C2660 a_n100_n23703# VSUBS 0.247431f
C2661 a_100_n20970# VSUBS 0.576721f
C2662 a_n158_n20970# VSUBS 0.576721f
C2663 a_n100_n21067# VSUBS 0.247431f
C2664 a_100_n18334# VSUBS 0.576721f
C2665 a_n158_n18334# VSUBS 0.576721f
C2666 a_n100_n18431# VSUBS 0.247431f
C2667 a_100_n15698# VSUBS 0.576721f
C2668 a_n158_n15698# VSUBS 0.576721f
C2669 a_n100_n15795# VSUBS 0.247431f
C2670 a_100_n13062# VSUBS 0.576721f
C2671 a_n158_n13062# VSUBS 0.576721f
C2672 a_n100_n13159# VSUBS 0.247431f
C2673 a_100_n10426# VSUBS 0.576721f
C2674 a_n158_n10426# VSUBS 0.576721f
C2675 a_n100_n10523# VSUBS 0.247431f
C2676 a_100_n7790# VSUBS 0.576721f
C2677 a_n158_n7790# VSUBS 0.576721f
C2678 a_n100_n7887# VSUBS 0.247431f
C2679 a_100_n5154# VSUBS 0.576721f
C2680 a_n158_n5154# VSUBS 0.576721f
C2681 a_n100_n5251# VSUBS 0.247431f
C2682 a_100_n2518# VSUBS 0.576721f
C2683 a_n158_n2518# VSUBS 0.576721f
C2684 a_n100_n2615# VSUBS 0.247431f
C2685 a_100_118# VSUBS 0.576721f
C2686 a_n158_118# VSUBS 0.576721f
C2687 a_n100_21# VSUBS 0.247431f
C2688 a_100_2754# VSUBS 0.576721f
C2689 a_n158_2754# VSUBS 0.576721f
C2690 a_n100_2657# VSUBS 0.247431f
C2691 a_100_5390# VSUBS 0.576721f
C2692 a_n158_5390# VSUBS 0.576721f
C2693 a_n100_5293# VSUBS 0.247431f
C2694 a_100_8026# VSUBS 0.576721f
C2695 a_n158_8026# VSUBS 0.576721f
C2696 a_n100_7929# VSUBS 0.247431f
C2697 a_100_10662# VSUBS 0.576721f
C2698 a_n158_10662# VSUBS 0.576721f
C2699 a_n100_10565# VSUBS 0.247431f
C2700 a_100_13298# VSUBS 0.576721f
C2701 a_n158_13298# VSUBS 0.576721f
C2702 a_n100_13201# VSUBS 0.247431f
C2703 a_100_15934# VSUBS 0.576721f
C2704 a_n158_15934# VSUBS 0.576721f
C2705 a_n100_15837# VSUBS 0.247431f
C2706 a_100_18570# VSUBS 0.576721f
C2707 a_n158_18570# VSUBS 0.576721f
C2708 a_n100_18473# VSUBS 0.247431f
C2709 a_100_21206# VSUBS 0.576721f
C2710 a_n158_21206# VSUBS 0.576721f
C2711 a_n100_21109# VSUBS 0.247431f
C2712 a_100_23842# VSUBS 0.576721f
C2713 a_n158_23842# VSUBS 0.576721f
C2714 a_n100_23745# VSUBS 0.247431f
C2715 a_100_26478# VSUBS 0.576721f
C2716 a_n158_26478# VSUBS 0.576721f
C2717 a_n100_26381# VSUBS 0.247431f
C2718 a_100_29114# VSUBS 0.576721f
C2719 a_n158_29114# VSUBS 0.576721f
C2720 a_n100_29017# VSUBS 0.247431f
C2721 a_100_31750# VSUBS 0.576721f
C2722 a_n158_31750# VSUBS 0.576721f
C2723 a_n100_31653# VSUBS 0.247431f
C2724 a_100_34386# VSUBS 0.576721f
C2725 a_n158_34386# VSUBS 0.576721f
C2726 a_n100_34289# VSUBS 0.247431f
C2727 a_100_37022# VSUBS 0.576721f
C2728 a_n158_37022# VSUBS 0.576721f
C2729 a_n100_36925# VSUBS 0.247431f
C2730 a_100_39658# VSUBS 0.576721f
C2731 a_n158_39658# VSUBS 0.576721f
C2732 a_n100_39561# VSUBS 0.247431f
C2733 a_100_42294# VSUBS 0.576721f
C2734 a_n158_42294# VSUBS 0.576721f
C2735 a_n100_42197# VSUBS 0.247431f
C2736 a_100_44930# VSUBS 0.576721f
C2737 a_n158_44930# VSUBS 0.576721f
C2738 a_n100_44833# VSUBS 0.247431f
C2739 a_100_47566# VSUBS 0.576721f
C2740 a_n158_47566# VSUBS 0.576721f
C2741 a_n100_47469# VSUBS 0.247431f
C2742 a_100_50202# VSUBS 0.576721f
C2743 a_n158_50202# VSUBS 0.576721f
C2744 a_n100_50105# VSUBS 0.247431f
C2745 a_100_52838# VSUBS 0.576721f
C2746 a_n158_52838# VSUBS 0.576721f
C2747 a_n100_52741# VSUBS 0.247431f
C2748 a_100_55474# VSUBS 0.576721f
C2749 a_n158_55474# VSUBS 0.576721f
C2750 a_n100_55377# VSUBS 0.247431f
C2751 a_100_58110# VSUBS 0.576721f
C2752 a_n158_58110# VSUBS 0.576721f
C2753 a_n100_58013# VSUBS 0.247431f
C2754 a_100_60746# VSUBS 0.576721f
C2755 a_n158_60746# VSUBS 0.576721f
C2756 a_n100_60649# VSUBS 0.247431f
C2757 a_100_63382# VSUBS 0.576721f
C2758 a_n158_63382# VSUBS 0.576721f
C2759 a_n100_63285# VSUBS 0.247431f
C2760 a_100_66018# VSUBS 0.576721f
C2761 a_n158_66018# VSUBS 0.576721f
C2762 a_n100_65921# VSUBS 0.247431f
C2763 a_100_68654# VSUBS 0.576721f
C2764 a_n158_68654# VSUBS 0.576721f
C2765 a_n100_68557# VSUBS 0.247431f
C2766 a_100_71290# VSUBS 0.576721f
C2767 a_n158_71290# VSUBS 0.576721f
C2768 a_n100_71193# VSUBS 0.247431f
C2769 a_100_73926# VSUBS 0.576721f
C2770 a_n158_73926# VSUBS 0.576721f
C2771 a_n100_73829# VSUBS 0.247431f
C2772 a_100_76562# VSUBS 0.576721f
C2773 a_n158_76562# VSUBS 0.576721f
C2774 a_n100_76465# VSUBS 0.247431f
C2775 a_100_79198# VSUBS 0.576721f
C2776 a_n158_79198# VSUBS 0.576721f
C2777 a_n100_79101# VSUBS 0.247431f
C2778 a_100_81834# VSUBS 0.576721f
C2779 a_n158_81834# VSUBS 0.576721f
C2780 a_n100_81737# VSUBS 0.247431f
C2781 a_100_84470# VSUBS 0.576721f
C2782 a_n158_84470# VSUBS 0.576721f
C2783 a_n100_84373# VSUBS 0.247431f
C2784 a_100_87106# VSUBS 0.576721f
C2785 a_n158_87106# VSUBS 0.576721f
C2786 a_n100_87009# VSUBS 0.247431f
C2787 a_100_89742# VSUBS 0.576721f
C2788 a_n158_89742# VSUBS 0.576721f
C2789 a_n100_89645# VSUBS 0.247431f
C2790 a_100_92378# VSUBS 0.576721f
C2791 a_n158_92378# VSUBS 0.576721f
C2792 a_n100_92281# VSUBS 0.247431f
C2793 a_100_95014# VSUBS 0.576721f
C2794 a_n158_95014# VSUBS 0.576721f
C2795 a_n100_94917# VSUBS 0.247431f
C2796 a_100_97650# VSUBS 0.576721f
C2797 a_n158_97650# VSUBS 0.576721f
C2798 a_n100_97553# VSUBS 0.247431f
C2799 a_100_100286# VSUBS 0.576721f
C2800 a_n158_100286# VSUBS 0.576721f
C2801 a_n100_100189# VSUBS 0.247431f
C2802 a_100_102922# VSUBS 0.576721f
C2803 a_n158_102922# VSUBS 0.576721f
C2804 a_n100_102825# VSUBS 0.247431f
C2805 a_100_105558# VSUBS 0.576721f
C2806 a_n158_105558# VSUBS 0.576721f
C2807 a_n100_105461# VSUBS 0.247431f
C2808 a_100_108194# VSUBS 0.576721f
C2809 a_n158_108194# VSUBS 0.576721f
C2810 a_n100_108097# VSUBS 0.247431f
C2811 a_100_110830# VSUBS 0.576721f
C2812 a_n158_110830# VSUBS 0.576721f
C2813 a_n100_110733# VSUBS 0.247431f
C2814 a_100_113466# VSUBS 0.576721f
C2815 a_n158_113466# VSUBS 0.576721f
C2816 a_n100_113369# VSUBS 0.247431f
C2817 a_100_116102# VSUBS 0.576721f
C2818 a_n158_116102# VSUBS 0.576721f
C2819 a_n100_116005# VSUBS 0.247431f
C2820 a_100_118738# VSUBS 0.576721f
C2821 a_n158_118738# VSUBS 0.576721f
C2822 a_n100_118641# VSUBS 0.247431f
C2823 a_100_121374# VSUBS 0.576721f
C2824 a_n158_121374# VSUBS 0.576721f
C2825 a_n100_121277# VSUBS 0.247431f
C2826 a_100_124010# VSUBS 0.576721f
C2827 a_n158_124010# VSUBS 0.576721f
C2828 a_n100_123913# VSUBS 0.247431f
C2829 a_100_126646# VSUBS 0.576721f
C2830 a_n158_126646# VSUBS 0.576721f
C2831 a_n100_126549# VSUBS 0.247431f
C2832 a_100_129282# VSUBS 0.576721f
C2833 a_n158_129282# VSUBS 0.576721f
C2834 a_n100_129185# VSUBS 0.247431f
C2835 a_100_131918# VSUBS 0.576721f
C2836 a_n158_131918# VSUBS 0.576721f
C2837 a_n100_131821# VSUBS 0.247431f
C2838 a_100_134554# VSUBS 0.576721f
C2839 a_n158_134554# VSUBS 0.576721f
C2840 a_n100_134457# VSUBS 0.247431f
C2841 a_100_137190# VSUBS 0.576721f
C2842 a_n158_137190# VSUBS 0.576721f
C2843 a_n100_137093# VSUBS 0.247431f
C2844 a_100_139826# VSUBS 0.576721f
C2845 a_n158_139826# VSUBS 0.576721f
C2846 a_n100_139729# VSUBS 0.247431f
C2847 a_100_142462# VSUBS 0.576721f
C2848 a_n158_142462# VSUBS 0.576721f
C2849 a_n100_142365# VSUBS 0.247431f
C2850 a_100_145098# VSUBS 0.576721f
C2851 a_n158_145098# VSUBS 0.576721f
C2852 a_n100_145001# VSUBS 0.247431f
C2853 a_100_147734# VSUBS 0.576721f
C2854 a_n158_147734# VSUBS 0.576721f
C2855 a_n100_147637# VSUBS 0.247431f
C2856 a_100_150370# VSUBS 0.576721f
C2857 a_n158_150370# VSUBS 0.576721f
C2858 a_n100_150273# VSUBS 0.247431f
C2859 a_100_153006# VSUBS 0.576721f
C2860 a_n158_153006# VSUBS 0.576721f
C2861 a_n100_152909# VSUBS 0.247431f
C2862 a_100_155642# VSUBS 0.576721f
C2863 a_n158_155642# VSUBS 0.576721f
C2864 a_n100_155545# VSUBS 0.247431f
C2865 a_100_158278# VSUBS 0.576721f
C2866 a_n158_158278# VSUBS 0.576721f
C2867 a_n100_158181# VSUBS 0.247431f
C2868 a_100_160914# VSUBS 0.576721f
C2869 a_n158_160914# VSUBS 0.576721f
C2870 a_n100_160817# VSUBS 0.247431f
C2871 a_100_163550# VSUBS 0.576721f
C2872 a_n158_163550# VSUBS 0.576721f
C2873 a_n100_163453# VSUBS 0.247431f
C2874 a_100_166186# VSUBS 0.576721f
C2875 a_n158_166186# VSUBS 0.576721f
C2876 a_n100_166089# VSUBS 0.247431f
C2877 a_100_168822# VSUBS 0.576721f
C2878 a_n158_168822# VSUBS 0.576721f
C2879 a_n100_168725# VSUBS 0.247431f
C2880 a_100_171458# VSUBS 0.576721f
C2881 a_n158_171458# VSUBS 0.576721f
C2882 a_n100_171361# VSUBS 0.247431f
C2883 a_100_174094# VSUBS 0.576721f
C2884 a_n158_174094# VSUBS 0.576721f
C2885 a_n100_173997# VSUBS 0.247431f
C2886 a_100_176730# VSUBS 0.576721f
C2887 a_n158_176730# VSUBS 0.576721f
C2888 a_n100_176633# VSUBS 0.247431f
C2889 a_100_179366# VSUBS 0.576721f
C2890 a_n158_179366# VSUBS 0.576721f
C2891 a_n100_179269# VSUBS 0.247431f
C2892 a_100_182002# VSUBS 0.576721f
C2893 a_n158_182002# VSUBS 0.576721f
C2894 a_n100_181905# VSUBS 0.247431f
C2895 a_100_184638# VSUBS 0.576721f
C2896 a_n158_184638# VSUBS 0.576721f
C2897 a_n100_184541# VSUBS 0.247431f
C2898 a_100_187274# VSUBS 0.576721f
C2899 a_n158_187274# VSUBS 0.576721f
C2900 a_n100_187177# VSUBS 0.247431f
C2901 a_100_189910# VSUBS 0.576721f
C2902 a_n158_189910# VSUBS 0.576721f
C2903 a_n100_189813# VSUBS 0.247431f
C2904 a_100_192546# VSUBS 0.576721f
C2905 a_n158_192546# VSUBS 0.576721f
C2906 a_n100_192449# VSUBS 0.247431f
C2907 a_100_195182# VSUBS 0.576721f
C2908 a_n158_195182# VSUBS 0.576721f
C2909 a_n100_195085# VSUBS 0.247431f
C2910 a_100_197818# VSUBS 0.576721f
C2911 a_n158_197818# VSUBS 0.576721f
C2912 a_n100_197721# VSUBS 0.247431f
C2913 a_100_200454# VSUBS 0.576721f
C2914 a_n158_200454# VSUBS 0.576721f
C2915 a_n100_200357# VSUBS 0.247431f
C2916 a_100_203090# VSUBS 0.576721f
C2917 a_n158_203090# VSUBS 0.576721f
C2918 a_n100_202993# VSUBS 0.247431f
C2919 a_100_205726# VSUBS 0.576721f
C2920 a_n158_205726# VSUBS 0.576721f
C2921 a_n100_205629# VSUBS 0.247431f
C2922 a_100_208362# VSUBS 0.576721f
C2923 a_n158_208362# VSUBS 0.576721f
C2924 a_n100_208265# VSUBS 0.247431f
C2925 a_100_210998# VSUBS 0.576721f
C2926 a_n158_210998# VSUBS 0.576721f
C2927 a_n100_210901# VSUBS 0.247431f
C2928 a_100_213634# VSUBS 0.576721f
C2929 a_n158_213634# VSUBS 0.576721f
C2930 a_n100_213537# VSUBS 0.247431f
C2931 a_100_216270# VSUBS 0.576721f
C2932 a_n158_216270# VSUBS 0.576721f
C2933 a_n100_216173# VSUBS 0.247431f
C2934 a_100_218906# VSUBS 0.576721f
C2935 a_n158_218906# VSUBS 0.576721f
C2936 a_n100_218809# VSUBS 0.247431f
C2937 a_100_221542# VSUBS 0.576721f
C2938 a_n158_221542# VSUBS 0.576721f
C2939 a_n100_221445# VSUBS 0.247431f
C2940 a_100_224178# VSUBS 0.576721f
C2941 a_n158_224178# VSUBS 0.576721f
C2942 a_n100_224081# VSUBS 0.247431f
C2943 a_100_226814# VSUBS 0.576721f
C2944 a_n158_226814# VSUBS 0.576721f
C2945 a_n100_226717# VSUBS 0.247431f
C2946 a_100_229450# VSUBS 0.576721f
C2947 a_n158_229450# VSUBS 0.576721f
C2948 a_n100_229353# VSUBS 0.247431f
C2949 a_100_232086# VSUBS 0.576721f
C2950 a_n158_232086# VSUBS 0.576721f
C2951 a_n100_231989# VSUBS 0.247431f
C2952 a_100_234722# VSUBS 0.576721f
C2953 a_n158_234722# VSUBS 0.576721f
C2954 a_n100_234625# VSUBS 0.247431f
C2955 a_100_237358# VSUBS 0.576721f
C2956 a_n158_237358# VSUBS 0.576721f
C2957 a_n100_237261# VSUBS 0.247431f
C2958 a_100_239994# VSUBS 0.576721f
C2959 a_n158_239994# VSUBS 0.576721f
C2960 a_n100_239897# VSUBS 0.247431f
C2961 a_100_242630# VSUBS 0.576721f
C2962 a_n158_242630# VSUBS 0.576721f
C2963 a_n100_242533# VSUBS 0.247431f
C2964 a_100_245266# VSUBS 0.576721f
C2965 a_n158_245266# VSUBS 0.576721f
C2966 a_n100_245169# VSUBS 0.247431f
C2967 a_100_247902# VSUBS 0.576721f
C2968 a_n158_247902# VSUBS 0.576721f
C2969 a_n100_247805# VSUBS 0.247431f
C2970 a_100_250538# VSUBS 0.576721f
C2971 a_n158_250538# VSUBS 0.576721f
C2972 a_n100_250441# VSUBS 0.247431f
C2973 a_100_253174# VSUBS 0.576721f
C2974 a_n158_253174# VSUBS 0.576721f
C2975 a_n100_253077# VSUBS 0.247431f
C2976 a_100_255810# VSUBS 0.576721f
C2977 a_n158_255810# VSUBS 0.576721f
C2978 a_n100_255713# VSUBS 0.247431f
C2979 a_100_258446# VSUBS 0.576721f
C2980 a_n158_258446# VSUBS 0.576721f
C2981 a_n100_258349# VSUBS 0.247431f
C2982 a_100_261082# VSUBS 0.576721f
C2983 a_n158_261082# VSUBS 0.576721f
C2984 a_n100_260985# VSUBS 0.247431f
C2985 a_100_263718# VSUBS 0.576721f
C2986 a_n158_263718# VSUBS 0.576721f
C2987 a_n100_263621# VSUBS 0.247431f
C2988 a_100_266354# VSUBS 0.576721f
C2989 a_n158_266354# VSUBS 0.576721f
C2990 a_n100_266257# VSUBS 0.247431f
C2991 a_100_268990# VSUBS 0.576721f
C2992 a_n158_268990# VSUBS 0.576721f
C2993 a_n100_268893# VSUBS 0.247431f
C2994 a_100_271626# VSUBS 0.576721f
C2995 a_n158_271626# VSUBS 0.576721f
C2996 a_n100_271529# VSUBS 0.247431f
C2997 a_100_274262# VSUBS 0.576721f
C2998 a_n158_274262# VSUBS 0.576721f
C2999 a_n100_274165# VSUBS 0.247431f
C3000 a_100_276898# VSUBS 0.576721f
C3001 a_n158_276898# VSUBS 0.576721f
C3002 a_n100_276801# VSUBS 0.247431f
C3003 a_100_279534# VSUBS 0.576721f
C3004 a_n158_279534# VSUBS 0.576721f
C3005 a_n100_279437# VSUBS 0.247431f
C3006 a_100_282170# VSUBS 0.576721f
C3007 a_n158_282170# VSUBS 0.576721f
C3008 a_n100_282073# VSUBS 0.247431f
C3009 a_100_284806# VSUBS 0.576721f
C3010 a_n158_284806# VSUBS 0.576721f
C3011 a_n100_284709# VSUBS 0.247431f
C3012 a_100_287442# VSUBS 0.576721f
C3013 a_n158_287442# VSUBS 0.576721f
C3014 a_n100_287345# VSUBS 0.247431f
C3015 a_100_290078# VSUBS 0.576721f
C3016 a_n158_290078# VSUBS 0.576721f
C3017 a_n100_289981# VSUBS 0.247431f
C3018 a_100_292714# VSUBS 0.576721f
C3019 a_n158_292714# VSUBS 0.576721f
C3020 a_n100_292617# VSUBS 0.247431f
C3021 a_100_295350# VSUBS 0.576721f
C3022 a_n158_295350# VSUBS 0.576721f
C3023 a_n100_295253# VSUBS 0.247431f
C3024 a_100_297986# VSUBS 0.576721f
C3025 a_n158_297986# VSUBS 0.576721f
C3026 a_n100_297889# VSUBS 0.247431f
C3027 a_100_300622# VSUBS 0.576721f
C3028 a_n158_300622# VSUBS 0.576721f
C3029 a_n100_300525# VSUBS 0.247431f
C3030 a_100_303258# VSUBS 0.576721f
C3031 a_n158_303258# VSUBS 0.576721f
C3032 a_n100_303161# VSUBS 0.247431f
C3033 a_100_305894# VSUBS 0.576721f
C3034 a_n158_305894# VSUBS 0.576721f
C3035 a_n100_305797# VSUBS 0.247431f
C3036 a_100_308530# VSUBS 0.576721f
C3037 a_n158_308530# VSUBS 0.576721f
C3038 a_n100_308433# VSUBS 0.247431f
C3039 a_100_311166# VSUBS 0.576721f
C3040 a_n158_311166# VSUBS 0.576721f
C3041 a_n100_311069# VSUBS 0.247431f
C3042 a_100_313802# VSUBS 0.576721f
C3043 a_n158_313802# VSUBS 0.576721f
C3044 a_n100_313705# VSUBS 0.247431f
C3045 a_100_316438# VSUBS 0.576721f
C3046 a_n158_316438# VSUBS 0.576721f
C3047 a_n100_316341# VSUBS 0.247431f
C3048 a_100_319074# VSUBS 0.576721f
C3049 a_n158_319074# VSUBS 0.576721f
C3050 a_n100_318977# VSUBS 0.247431f
C3051 a_100_321710# VSUBS 0.576721f
C3052 a_n158_321710# VSUBS 0.576721f
C3053 a_n100_321613# VSUBS 0.247431f
C3054 a_100_324346# VSUBS 0.576721f
C3055 a_n158_324346# VSUBS 0.576721f
C3056 a_n100_324249# VSUBS 0.247431f
C3057 a_100_326982# VSUBS 0.576721f
C3058 a_n158_326982# VSUBS 0.576721f
C3059 a_n100_326885# VSUBS 0.247431f
C3060 a_100_329618# VSUBS 0.576721f
C3061 a_n158_329618# VSUBS 0.576721f
C3062 a_n100_329521# VSUBS 0.247431f
C3063 a_100_332254# VSUBS 0.576721f
C3064 a_n158_332254# VSUBS 0.576721f
C3065 a_n100_332157# VSUBS 0.247431f
C3066 a_100_334890# VSUBS 0.58217f
C3067 a_n158_334890# VSUBS 0.58217f
C3068 a_n100_334793# VSUBS 0.291162f
C3069 w_n358_n337587# VSUBS 1.79542p
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_GK83LR a_100_n4026# a_100_n74474# a_n100_74613#
+ a_100_88178# a_n158_21874# a_100_93358# a_100_49846# a_n100_n63175# a_n100_n19663#
+ a_n158_86106# a_100_n34070# a_n158_n45466# a_n100_4165# a_n100_113981# a_100_n11278#
+ a_n100_n24843# a_n100_11417# a_n158_n50646# a_n158_82998# a_n100_n109795# a_n158_n116950#
+ a_100_14622# a_100_n95194# a_n100_n114975# a_n100_95333# a_n158_42594# a_n158_n10242#
+ a_n100_n85967# a_100_115114# a_100_n56862# a_n100_115017# a_n158_n66186# a_100_75746#
+ a_n100_n45563# a_n100_32137# a_n158_n27854# a_n158_n71366# a_n158_7370# a_100_80926#
+ a_n158_n109698# a_n100_n50743# a_100_n106590# a_n158_105790# a_100_35342# a_n158_n114878#
+ a_100_n111770# a_n158_110970# a_100_40522# a_100_n7134# a_100_2190# a_n100_49749#
+ a_100_n77582# a_n158_n88978# a_n100_77721# a_n158_24982# a_n100_54929# a_100_n82762#
+ a_n100_82901# a_100_96466# a_n100_n66283# a_n100_n100471# a_n100_7273# a_n158_89214#
+ a_n158_n48574# a_n158_n92086# a_n158_n1954# a_100_n14386# a_n100_n27951# a_n100_n71463#
+ a_n100_14525# a_n158_5298# a_100_56062# a_n158_112006# a_n158_n53754# a_100_n132490#
+ a_100_61242# a_n158_131690# a_100_17730# a_n158_26018# a_n100_98441# a_n158_n13350#
+ a_100_22910# a_n100_75649# a_100_n59970# a_100_118222# a_n100_118125# a_n158_129618#
+ a_n158_50882# a_n100_n121191# a_n158_n100374# a_n100_80829# a_100_123402# a_n158_n69294#
+ a_100_78854# a_n100_n92183# a_n100_123305# a_n100_n48671# a_n100_35245# a_n100_n25879#
+ a_n158_n74474# a_100_n40286# a_n100_n53851# a_n100_n119119# a_n100_40425# a_100_38450#
+ a_n158_n117986# a_100_15658# a_n158_n34070# a_100_43630# a_n100_96369# a_n158_n11278#
+ a_100_20838# a_n100_n1015# a_100_n57898# a_n158_n121094# a_100_n85870# a_100_99574#
+ a_n100_n69391# a_n158_n95194# a_n100_n46599# a_n100_n74571# a_n100_61145# a_100_n17494#
+ a_100_8406# a_n100_17633# a_n158_97502# a_n158_n56862# a_100_59170# a_n158_115114#
+ a_n100_n51779# a_100_n22674# a_n100_22813# a_100_36378# a_100_64350# a_n158_29126#
+ a_100_41558# a_n100_n11375# a_n158_34306# a_n100_78757# a_n158_53990# a_100_n83798#
+ a_n158_n103482# a_n100_83937# a_100_126510# a_n100_126413# a_n100_n95291# a_n100_38353#
+ a_100_103718# a_n158_n77582# a_n100_n28987# a_n100_n72499# a_100_n43394# a_n100_43533#
+ a_100_57098# a_100_85070# a_n158_n82762# a_n100_n127407# a_100_18766# a_100_62278#
+ a_n100_n32095# a_100_90250# a_n158_55026# a_n100_99477# a_n158_n14386# a_100_23946#
+ a_n100_n4123# a_n158_60206# a_100_119258# a_n100_59073# a_100_124438# a_n100_108801#
+ a_n100_64253# a_n158_n59970# a_100_n119022# a_n158_118222# a_n100_n54887# a_n158_77818#
+ w_n358_n132787# a_100_n25782# a_n100_25921# a_100_39486# a_100_n124202# a_n158_123402#
+ a_100_n30962# a_100_44666# a_n100_n14483# a_n158_37414# a_n158_n40286# a_n158_n106590#
+ a_n158_n9206# a_n100_129521# a_100_106826# a_n158_n111770# a_n100_106729# a_n100_18669#
+ a_n100_90153# a_n158_98538# a_n100_46641# a_n158_n57898# a_n100_111909# a_n100_n80787#
+ a_n158_n85870# a_n100_23849# a_100_n51682# a_100_65386# a_n100_51821# a_n158_58134#
+ a_n158_n17494# a_100_70566# a_n100_n7231# a_n100_n40383# a_n158_63314# a_n158_19802#
+ a_n158_n22674# a_n158_2190# a_100_127546# a_n158_n132490# a_n100_127449# a_100_30162#
+ a_n100_39389# a_n100_67361# a_n100_n57995# a_n100_44569# a_n100_72541# a_100_n28890#
+ a_n158_n83798# a_100_n127310# a_n158_126510# a_100_47774# a_100_91286# a_n158_103718#
+ a_100_n104518# a_n100_n17591# a_n158_84034# a_n158_118# a_n100_2093# a_n100_n5159#
+ a_n158_n43394# a_100_n98302# a_100_52954# a_n100_n22771# a_n158_45702# a_n100_n116011#
+ a_n100_21# a_n100_88081# a_100_109934# a_n100_n87003# a_100_12550# a_n100_109837#
+ a_n100_65289# a_n100_93261# a_n158_119258# a_100_n35106# a_n100_n83895# a_n100_26957#
+ a_n100_70469# a_100_113042# a_100_n54790# a_100_n125238# a_100_68494# a_n158_124438#
+ a_100_n31998# a_100_73674# a_100_n130418# a_n100_n43491# a_n100_30065# a_n158_66422#
+ a_100_28090# a_n100_n20699# a_n158_n25782# a_n158_71602# a_100_33270# a_n158_n30962#
+ a_100_10478# a_100_n5062# a_n100_47677# a_n100_91189# a_100_n61006# a_n158_8406#
+ a_100_n80690# a_n100_52857# a_100_94394# a_100_n107626# a_n158_106826# a_n158_87142#
+ a_100_100610# a_n100_n8267# a_100_n112806# a_n100_100513# a_n100_12453# a_n158_92322#
+ a_100_3226# a_n158_48810# a_n158_n51682# a_100_n78618# a_100_31198# a_n100_68397#
+ a_n100_n67319# a_100_n38214# a_n100_n101507# a_n100_8309# a_n100_73577# a_100_116150#
+ a_100_n128346# a_n100_116053# a_n158_127546# a_100_76782# a_100_121330# a_n100_121233#
+ a_n100_33173# a_100_n99338# a_n158_69530# a_n158_n28890# a_n158_n119022# a_100_81962#
+ a_n158_46738# a_n100_n117047# a_n158_74710# a_n158_n124202# a_n100_n88039# a_100_13586#
+ a_n158_51918# a_n100_n122227# a_100_n8170# a_n100_94297# a_n100_n93219# a_n158_n98302#
+ a_n100_n49707# a_100_n64114# a_100_114078# a_n158_11514# a_n100_55965# a_n158_109934#
+ a_n158_n35106# a_100_n115914# a_n158_67458# a_n100_103621# a_n158_n2990# a_n100_15561#
+ a_n158_95430# a_100_6334# a_n158_113042# a_n158_n54790# a_n158_72638# a_n158_n31998#
+ a_n100_20741# a_100_n86906# a_n158_27054# a_100_n6098# a_n100_n104615# a_n158_32234#
+ a_n100_76685# a_n100_n75607# a_100_n90014# a_n100_119161# a_100_n46502# a_n100_81865#
+ a_n158_n4026# a_100_79890# a_n158_88178# a_n100_124341# a_n100_36281# a_100_101646#
+ a_n100_n35203# a_n100_101549# a_n100_13489# a_n158_93358# a_n158_n61006# a_n100_41461#
+ a_n158_49846# a_n158_n80690# a_n158_n127310# a_100_16694# a_n100_n125335# a_n158_n104518#
+ a_100_n101410# a_n158_100610# a_n100_n96327# a_100_n67222# a_n100_n130515# a_100_21874#
+ a_n100_n2051# a_n158_n78618# a_100_117186# a_n158_14622# a_n100_117089# a_100_n72402#
+ a_100_86106# a_100_122366# a_n100_122269# a_n158_n38214# a_n100_62181# a_n100_n61103#
+ a_100_9442# a_100_82998# a_n158_116150# a_n158_75746# a_n158_n125238# a_n158_121330#
+ a_100_n122130# a_n158_80926# a_n158_n130418# a_n100_n107723# a_100_42594# a_n158_n99338#
+ a_n158_35342# a_n100_79793# a_n100_n78715# a_100_n49610# a_100_n93122# a_n100_n112903#
+ a_n158_40522# a_n100_84973# a_n158_n7134# a_100_n26818# a_100_104754# a_n100_n38311#
+ a_n100_104657# a_n158_n64114# a_n100_16597# a_n158_96466# a_n100_n15519# a_n158_114078#
+ a_n100_21777# a_n100_n128443# a_100_n120058# a_n158_n107626# a_n158_56062# a_n100_n99435#
+ a_100_24982# a_n100_86009# a_n158_n112806# a_n158_61242# a_n158_17730# a_100_n47538#
+ a_100_n75510# a_100_89214# a_100_125474# a_n158_n86906# a_n158_22910# a_100_n52718#
+ a_n100_n59031# a_n100_125377# a_100_n1954# a_n100_n36239# a_100_130654# a_n100_n64211#
+ a_n100_130557# a_n100_42497# a_n158_n46502# a_n158_n90014# a_n100_5201# a_n158_78854#
+ a_n100_n41419# a_n158_n128346# a_100_n12314# a_100_26018# a_n158_3226# a_100_n102446#
+ a_n158_101646# a_100_n68258# a_n158_38450# a_n100_n3087# a_100_50882# a_100_n96230#
+ a_n158_15658# a_n158_43630# a_100_n29926# a_100_n73438# a_100_n918# a_n158_20838#
+ a_100_107862# a_n100_107765# a_n100_n62139# a_n158_n67222# a_n158_99574# a_n100_n18627#
+ a_n100_n90111# a_n158_117186# a_100_n33034# a_n100_3129# a_n100_112945# a_n100_24885#
+ a_n100_n23807# a_n158_n72402# a_n158_122366# a_100_n123166# a_n158_59170# a_n100_n108759#
+ a_n100_89117# a_n158_n115914# a_n158_36378# a_n158_64350# a_100_n94158# a_n100_n113939#
+ a_n158_41558# a_100_128582# a_n100_128485# a_100_n55826# a_100_97502# a_n100_n39347#
+ a_n100_n44527# a_n158_n49610# a_n158_n93122# a_100_n15422# a_n158_n26818# a_n158_6334#
+ a_100_29126# a_n100_n129479# a_n100_50785# a_100_n105554# a_n158_104754# a_100_n20602#
+ a_100_34306# a_n158_57098# a_n158_85070# a_n100_n6195# a_100_n110734# a_100_53990#
+ a_n158_62278# a_n100_10381# a_n158_18766# a_n158_90250# a_100_1154# a_100_n76546#
+ a_n158_23946# a_100_n81726# a_n158_n101410# a_n100_n65247# a_100_n36142# a_n158_n47538#
+ a_n100_6237# a_n158_n75510# a_n100_27993# a_n100_n26915# a_n100_n70427# a_100_n126274#
+ a_n158_125474# a_100_n41322# a_100_55026# a_n158_n52718# a_100_n131454# a_n158_130654#
+ a_n158_39486# a_100_60206# a_n100_n30023# a_100_n97266# a_n100_97405# a_n158_44666#
+ a_n158_n12314# a_100_n58934# a_n158_n122130# a_100_108898# a_n100_n120155# a_n100_29029#
+ a_n158_n68258# a_n100_57001# a_100_77818# a_n158_n96230# a_n100_n47635# a_n100_n91147#
+ a_n100_34209# a_100_n18530# a_100_n62042# a_n158_n29926# a_n158_n73438# a_n158_9442#
+ a_n100_53893# a_n100_n52815# a_100_n108662# a_n158_107862# a_100_n23710# a_100_37414#
+ a_n158_n33034# a_100_n113842# a_n158_65386# a_100_n9206# a_n100_n12411# a_100_n79654#
+ a_100_4262# a_n158_70566# a_n158_n120058# a_100_n84834# a_100_98538# a_n100_n68355#
+ a_100_n39250# a_n100_n102543# a_n100_9345# a_n158_n94158# a_n158_30162# a_n100_n73535#
+ a_n100_60109# a_100_n16458# a_100_n129382# a_n158_128582# a_100_n44430# a_100_58134#
+ a_n158_n55826# a_100_n21638# a_100_63314# a_100_19802# a_n100_n33131# a_n158_91286#
+ a_n158_n15422# a_n158_47774# a_n100_n10339# a_n100_n118083# a_n158_52954# a_n158_n20602#
+ a_n100_n89075# a_n100_n123263# a_n158_n102446# a_100_n37178# a_n100_n94255# a_n100_37317#
+ a_100_n65150# a_n158_n76546# a_n158_12550# a_100_n42358# a_n100_n55923# a_100_n70330#
+ a_100_84034# a_n158_n81726# a_100_120294# a_n100_120197# a_100_n116950# a_n100_n31059#
+ a_n158_n36142# a_100_45702# a_n158_68494# a_100_7370# a_n158_73674# a_n158_n41322#
+ a_n158_n123166# a_100_n87942# a_n158_28090# a_n158_n918# a_n100_58037# a_n158_n97266#
+ a_n100_n105651# a_n158_33270# a_100_n19566# a_100_n63078# a_n100_n76643# a_n100_63217#
+ a_100_n91050# a_n100_n110831# a_n100_19705# a_n158_n58934# a_n158_10478# a_100_n109698#
+ a_n158_108898# a_n158_n5062# a_100_n24746# a_n100_n81823# a_100_118# a_100_66422#
+ a_100_102682# a_100_n114878# a_n100_102585# a_n158_94394# a_n100_n13447# a_n158_n18530#
+ a_n158_n62042# a_100_5298# a_100_71602# a_n158_n23710# a_n100_n126371# a_n158_n105554#
+ a_n100_n97363# a_n100_n103579# a_n100_n131551# a_n158_n110734# a_n158_31198# a_n158_n79654#
+ a_100_n45466# a_n100_45605# a_100_87142# a_n158_n84834# a_100_n50646# a_100_92322#
+ a_n100_n34167# a_n158_n39250# a_100_48810# a_n158_n16458# a_n158_n44430# a_n158_76782#
+ a_n158_n126274# a_100_n10242# a_n158_n21638# a_n158_1154# a_n100_n124299# a_n158_81962#
+ a_n158_n131454# a_100_n100374# a_100_n66186# a_n100_n79751# a_n100_66325# a_n158_13586#
+ a_n100_n56959# a_n158_n8170# a_100_n71366# a_n100_n84931# a_n100_71505# a_100_n27854#
+ a_100_69530# a_100_105790# a_n158_n37178# a_100_n117986# a_100_46738# a_n100_105693#
+ a_n158_n65150# a_100_74710# a_n100_n16555# a_n100_n60067# a_100_110970# a_n100_1057#
+ a_n100_31101# a_n100_110873# a_n158_n42358# a_100_51918# a_n158_n70330# a_n100_n21735#
+ a_100_n88978# a_100_n121094# a_n158_n108662# a_n158_120294# a_n100_n106687# a_n100_87045#
+ a_n158_n113842# a_100_11514# a_n100_n77679# a_100_n48574# a_100_n92086# a_n100_n111867#
+ a_n100_92225# a_n100_48713# a_n158_n87942# a_n158_n6098# a_n100_n82859# a_100_n53754#
+ a_100_67458# a_100_112006# a_100_n2990# a_100_95430# a_n100_n37275# a_100_131690#
+ a_n100_131593# a_n158_n19566# a_n158_n63078# a_100_72638# a_n100_n42455# a_n158_n91050#
+ a_n158_79890# a_n100_n9303# a_n158_n129382# a_100_n13350# a_n158_4262# a_100_27054#
+ a_n158_n24746# a_n158_102682# a_100_129618# VSUBS a_100_n103482# a_100_32234# a_n100_n98399#
+ a_100_n69294# a_n100_n132587# a_n100_69433# a_n158_16694#
X0 a_100_n104518# a_n100_n104615# a_n158_n104518# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X1 a_100_n126274# a_n100_n126371# a_n158_n126274# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X2 a_100_n117986# a_n100_n118083# a_n158_n117986# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X3 a_100_n69294# a_n100_n69391# a_n158_n69294# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X4 a_100_119258# a_n100_119161# a_n158_119258# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X5 a_100_74710# a_n100_74613# a_n158_74710# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X6 a_100_n91050# a_n100_n91147# a_n158_n91050# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X7 a_100_50882# a_n100_50785# a_n158_50882# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X8 a_100_48810# a_n100_48713# a_n158_48810# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X9 a_100_11514# a_n100_11417# a_n158_11514# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X10 a_100_7370# a_n100_7273# a_n158_7370# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X11 a_100_n122130# a_n100_n122227# a_n158_n122130# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X12 a_100_n65150# a_n100_n65247# a_n158_n65150# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X13 a_100_24982# a_n100_24885# a_n158_24982# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X14 a_100_33270# a_n100_33173# a_n158_33270# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X15 a_100_n39250# a_n100_n39347# a_n158_n39250# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X16 a_100_92322# a_n100_92225# a_n158_92322# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X17 a_100_3226# a_n100_3129# a_n158_3226# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X18 a_100_n109698# a_n100_n109795# a_n158_n109698# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X19 a_100_20838# a_n100_20741# a_n158_20838# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X20 a_100_121330# a_n100_121233# a_n158_121330# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X21 a_100_66422# a_n100_66325# a_n158_66422# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X22 a_100_79890# a_n100_79793# a_n158_79890# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X23 a_100_42594# a_n100_42497# a_n158_42594# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X24 a_100_16694# a_n100_16597# a_n158_16694# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X25 a_100_n41322# a_n100_n41419# a_n158_n41322# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X26 a_100_130654# a_n100_130557# a_n158_130654# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X27 a_100_84034# a_n100_83937# a_n158_84034# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X28 a_100_75746# a_n100_75649# a_n158_75746# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X29 a_100_n15422# a_n100_n15519# a_n158_n15422# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X30 a_100_113042# a_n100_112945# a_n158_113042# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X31 a_100_104754# a_n100_104657# a_n158_104754# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X32 a_100_58134# a_n100_58037# a_n158_58134# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X33 a_100_49846# a_n100_49749# a_n158_49846# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X34 a_100_93358# a_n100_93261# a_n158_93358# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X35 a_100_n87942# a_n100_n88039# a_n158_n87942# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X36 a_100_n50646# a_n100_n50743# a_n158_n50646# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X37 a_100_n24746# a_n100_n24843# a_n158_n24746# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X38 a_100_122366# a_n100_122269# a_n158_122366# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X39 a_100_67458# a_n100_67361# a_n158_67458# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X40 a_100_n33034# a_n100_n33131# a_n158_n33034# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X41 a_100_n103482# a_n100_n103579# a_n158_n103482# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X42 a_100_n5062# a_n100_n5159# a_n158_n5062# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X43 a_100_118# a_n100_21# a_n158_118# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X44 a_100_n79654# a_n100_n79751# a_n158_n79654# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X45 a_100_n42358# a_n100_n42455# a_n158_n42358# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X46 a_100_129618# a_n100_129521# a_n158_129618# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X47 a_100_n16458# a_n100_n16555# a_n158_n16458# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X48 a_100_114078# a_n100_113981# a_n158_114078# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X49 a_100_n121094# a_n100_n121191# a_n158_n121094# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X50 a_100_n119022# a_n100_n119119# a_n158_n119022# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X51 a_100_n75510# a_n100_n75607# a_n158_n75510# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X52 a_100_43630# a_n100_43533# a_n158_43630# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X53 a_100_2190# a_n100_2093# a_n158_2190# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X54 a_100_n97266# a_n100_n97363# a_n158_n97266# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X55 a_100_n88978# a_n100_n89075# a_n158_n88978# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X56 a_100_n49610# a_n100_n49707# a_n158_n49610# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X57 a_100_17730# a_n100_17633# a_n158_17730# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X58 a_100_n34070# a_n100_n34167# a_n158_n34070# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X59 a_100_n128346# a_n100_n128443# a_n158_n128346# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X60 a_100_61242# a_n100_61145# a_n158_61242# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X61 a_100_52954# a_n100_52857# a_n158_52954# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X62 a_100_9442# a_n100_9345# a_n158_9442# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X63 a_100_n6098# a_n100_n6195# a_n158_n6098# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X64 a_100_35342# a_n100_35245# a_n158_35342# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X65 a_100_70566# a_n100_70469# a_n158_70566# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X66 a_100_123402# a_n100_123305# a_n158_123402# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X67 a_100_n10242# a_n100_n10339# a_n158_n10242# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X68 a_100_44666# a_n100_44569# a_n158_44666# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X69 a_100_27054# a_n100_26957# a_n158_27054# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X70 a_100_18766# a_n100_18669# a_n158_18766# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X71 a_100_n82762# a_n100_n82859# a_n158_n82762# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X72 a_100_86106# a_n100_86009# a_n158_86106# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X73 a_100_77818# a_n100_77721# a_n158_77818# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X74 a_100_62278# a_n100_62181# a_n158_62278# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X75 a_100_n113842# a_n100_n113939# a_n158_n113842# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X76 a_100_n56862# a_n100_n56959# a_n158_n56862# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X77 a_100_115114# a_n100_115017# a_n158_115114# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X78 a_100_106826# a_n100_106729# a_n158_106826# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X79 a_100_99574# a_n100_99477# a_n158_99574# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X80 a_100_36378# a_n100_36281# a_n158_36378# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X81 a_100_128582# a_n100_128485# a_n158_128582# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X82 a_100_n98302# a_n100_n98399# a_n158_n98302# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X83 a_100_n61006# a_n100_n61103# a_n158_n61006# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X84 a_100_n52718# a_n100_n52815# a_n158_n52718# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X85 a_100_n26818# a_n100_n26915# a_n158_n26818# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X86 a_100_n74474# a_n100_n74571# a_n158_n74474# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X87 a_100_124438# a_n100_124341# a_n158_124438# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X88 a_100_n131454# a_n100_n131551# a_n158_n131454# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X89 a_100_n35106# a_n100_n35203# a_n158_n35106# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X90 a_100_n11278# a_n100_n11375# a_n158_n11278# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X91 a_100_n105554# a_n100_n105651# a_n158_n105554# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X92 a_100_n48574# a_n100_n48671# a_n158_n48574# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X93 a_100_n7134# a_n100_n7231# a_n158_n7134# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X94 a_100_n70330# a_n100_n70427# a_n158_n70330# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X95 a_100_n83798# a_n100_n83895# a_n158_n83798# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X96 a_100_n101410# a_n100_n101507# a_n158_n101410# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X97 a_100_n92086# a_n100_n92183# a_n158_n92086# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X98 a_100_n44430# a_n100_n44527# a_n158_n44430# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X99 a_100_12550# a_n100_12453# a_n158_12550# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X100 a_100_n66186# a_n100_n66283# a_n158_n66186# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X101 a_100_n57898# a_n100_n57995# a_n158_n57898# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X102 a_100_n18530# a_n100_n18627# a_n158_n18530# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X103 a_100_n123166# a_n100_n123263# a_n158_n123166# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X104 a_100_n114878# a_n100_n114975# a_n158_n114878# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X105 a_100_71602# a_n100_71505# a_n158_71602# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X106 a_100_4262# a_n100_4165# a_n158_4262# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X107 a_100_100610# a_n100_100513# a_n158_100610# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X108 a_100_45702# a_n100_45605# a_n158_45702# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X109 a_100_n99338# a_n100_n99435# a_n158_n99338# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X110 a_100_30162# a_n100_30065# a_n158_30162# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X111 a_100_21874# a_n100_21777# a_n158_21874# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X112 a_100_19802# a_n100_19705# a_n158_19802# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X113 a_100_n132490# a_n100_n132587# a_n158_n132490# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X114 a_100_80926# a_n100_80829# a_n158_80926# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X115 a_100_n20602# a_n100_n20699# a_n158_n20602# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X116 a_100_n106590# a_n100_n106687# a_n158_n106590# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X117 a_100_63314# a_n100_63217# a_n158_63314# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X118 a_100_n8170# a_n100_n8267# a_n158_n8170# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X119 a_100_76782# a_n100_76685# a_n158_76782# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X120 a_100_131690# a_n100_131593# a_n158_131690# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X121 a_100_85070# a_n100_84973# a_n158_85070# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X122 a_100_37414# a_n100_37317# a_n158_37414# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X123 a_100_105790# a_n100_105693# a_n158_105790# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X124 a_100_59170# a_n100_59073# a_n158_59170# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X125 a_100_13586# a_n100_13489# a_n158_13586# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X126 a_100_72638# a_n100_72541# a_n158_72638# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X127 a_100_5298# a_n100_5201# a_n158_5298# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X128 a_100_n12314# a_n100_n12411# a_n158_n12314# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X129 a_100_n51682# a_n100_n51779# a_n158_n51682# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X130 a_100_101646# a_n100_101549# a_n158_101646# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X131 a_100_94394# a_n100_94297# a_n158_94394# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X132 a_100_55026# a_n100_54929# a_n158_55026# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X133 a_100_46738# a_n100_46641# a_n158_46738# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X134 a_100_n1954# a_n100_n2051# a_n158_n1954# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X135 a_100_31198# a_n100_31101# a_n158_31198# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X136 a_100_n25782# a_n100_n25879# a_n158_n25782# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X137 a_100_68494# a_n100_68397# a_n158_68494# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X138 a_100_29126# a_n100_29029# a_n158_29126# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X139 a_100_n93122# a_n100_n93219# a_n158_n93122# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X140 a_100_n84834# a_n100_n84931# a_n158_n84834# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X141 a_100_n21638# a_n100_n21735# a_n158_n21638# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X142 a_100_n115914# a_n100_n116011# a_n158_n115914# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X143 a_100_n67222# a_n100_n67319# a_n158_n67222# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X144 a_100_n58934# a_n100_n59031# a_n158_n58934# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X145 a_100_n124202# a_n100_n124299# a_n158_n124202# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X146 a_100_n43394# a_n100_n43491# a_n158_n43394# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X147 a_100_n100374# a_n100_n100471# a_n158_n100374# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X148 a_100_n17494# a_n100_n17591# a_n158_n17494# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X149 a_100_22910# a_n100_22813# a_n158_22910# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X150 a_100_n76546# a_n100_n76643# a_n158_n76546# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X151 a_100_n2990# a_n100_n3087# a_n158_n2990# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X152 a_100_n13350# a_n100_n13447# a_n158_n13350# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X153 a_100_n9206# a_n100_n9303# a_n158_n9206# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X154 a_100_n107626# a_n100_n107723# a_n158_n107626# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X155 a_100_n129382# a_n100_n129479# a_n158_n129382# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X156 a_100_40522# a_n100_40425# a_n158_40522# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X157 a_100_n94158# a_n100_n94255# a_n158_n94158# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X158 a_100_n85870# a_n100_n85967# a_n158_n85870# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X159 a_100_53990# a_n100_53893# a_n158_53990# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X160 a_100_n59970# a_n100_n60067# a_n158_n59970# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X161 a_100_14622# a_n100_14525# a_n158_14622# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X162 a_100_n125238# a_n100_n125335# a_n158_n125238# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X163 a_100_n116950# a_n100_n117047# a_n158_n116950# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X164 a_100_n68258# a_n100_n68355# a_n158_n68258# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X165 a_100_6334# a_n100_6237# a_n158_6334# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X166 a_100_95430# a_n100_95333# a_n158_95430# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X167 a_100_69530# a_n100_69433# a_n158_69530# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X168 a_100_32234# a_n100_32137# a_n158_32234# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X169 a_100_23946# a_n100_23849# a_n158_23946# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X170 a_100_28090# a_n100_27993# a_n158_28090# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X171 a_100_78854# a_n100_78757# a_n158_78854# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X172 a_100_41558# a_n100_41461# a_n158_41558# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X173 a_100_87142# a_n100_87045# a_n158_87142# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X174 a_100_15658# a_n100_15561# a_n158_15658# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X175 a_100_116150# a_n100_116053# a_n158_116150# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X176 a_100_107862# a_n100_107765# a_n158_107862# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X177 a_100_n62042# a_n100_n62139# a_n158_n62042# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X178 a_100_n53754# a_n100_n53851# a_n158_n53754# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X179 a_100_103718# a_n100_103621# a_n158_103718# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X180 a_100_96466# a_n100_96369# a_n158_96466# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X181 a_100_n110734# a_n100_n110831# a_n158_n110734# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X182 a_100_112006# a_n100_111909# a_n158_112006# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X183 a_100_n27854# a_n100_n27951# a_n158_n27854# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X184 a_100_n36142# a_n100_n36239# a_n158_n36142# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X185 a_100_125474# a_n100_125377# a_n158_125474# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X186 a_100_n918# a_n100_n1015# a_n158_n918# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X187 a_100_n86906# a_n100_n87003# a_n158_n86906# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X188 a_100_n23710# a_n100_n23807# a_n158_n23710# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X189 a_100_n71366# a_n100_n71463# a_n158_n71366# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X190 a_100_n45466# a_n100_n45563# a_n158_n45466# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X191 a_100_88178# a_n100_88081# a_n158_88178# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X192 a_100_n102446# a_n100_n102543# a_n158_n102446# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X193 a_100_n4026# a_n100_n4123# a_n158_n4026# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X194 a_100_n19566# a_n100_n19663# a_n158_n19566# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X195 a_100_117186# a_n100_117089# a_n158_117186# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X196 a_100_108898# a_n100_108801# a_n158_108898# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X197 a_100_n80690# a_n100_n80787# a_n158_n80690# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X198 a_100_n78618# a_n100_n78715# a_n158_n78618# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X199 a_100_n120058# a_n100_n120155# a_n158_n120058# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X200 a_100_n111770# a_n100_n111867# a_n158_n111770# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X201 a_100_n63078# a_n100_n63175# a_n158_n63078# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X202 a_100_n54790# a_n100_n54887# a_n158_n54790# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X203 a_100_n28890# a_n100_n28987# a_n158_n28890# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X204 a_100_1154# a_n100_1057# a_n158_1154# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X205 a_100_n37178# a_n100_n37275# a_n158_n37178# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X206 a_100_90250# a_n100_90153# a_n158_90250# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X207 a_100_81962# a_n100_81865# a_n158_81962# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X208 a_100_n96230# a_n100_n96327# a_n158_n96230# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X209 a_100_110970# a_n100_110873# a_n158_110970# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X210 a_100_64350# a_n100_64253# a_n158_64350# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X211 a_100_n127310# a_n100_n127407# a_n158_n127310# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X212 a_100_38450# a_n100_38353# a_n158_38450# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X213 a_100_60206# a_n100_60109# a_n158_60206# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X214 a_100_51918# a_n100_51821# a_n158_51918# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X215 a_100_8406# a_n100_8309# a_n158_8406# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X216 a_100_97502# a_n100_97405# a_n158_97502# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X217 a_100_n30962# a_n100_n31059# a_n158_n30962# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X218 a_100_73674# a_n100_73577# a_n158_73674# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X219 a_100_34306# a_n100_34209# a_n158_34306# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X220 a_100_126510# a_n100_126413# a_n158_126510# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X221 a_100_47774# a_n100_47677# a_n158_47774# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X222 a_100_10478# a_n100_10381# a_n158_10478# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X223 a_100_102682# a_n100_102585# a_n158_102682# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X224 a_100_56062# a_n100_55965# a_n158_56062# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X225 a_100_n72402# a_n100_n72499# a_n158_n72402# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X226 a_100_91286# a_n100_91189# a_n158_91286# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X227 a_100_82998# a_n100_82901# a_n158_82998# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X228 a_100_n46502# a_n100_n46599# a_n158_n46502# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X229 a_100_89214# a_n100_89117# a_n158_89214# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X230 a_100_n22674# a_n100_n22771# a_n158_n22674# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X231 a_100_120294# a_n100_120197# a_n158_120294# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X232 a_100_65386# a_n100_65289# a_n158_65386# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X233 a_100_26018# a_n100_25921# a_n158_26018# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X234 a_100_118222# a_n100_118125# a_n158_118222# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X235 a_100_109934# a_n100_109837# a_n158_109934# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X236 a_100_n90014# a_n100_n90111# a_n158_n90014# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X237 a_100_n81726# a_n100_n81823# a_n158_n81726# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X238 a_100_39486# a_n100_39389# a_n158_39486# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X239 a_100_n55826# a_n100_n55923# a_n158_n55826# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X240 a_100_98538# a_n100_98441# a_n158_98538# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X241 a_100_n31998# a_n100_n32095# a_n158_n31998# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X242 a_100_n112806# a_n100_n112903# a_n158_n112806# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X243 a_100_n64114# a_n100_n64211# a_n158_n64114# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X244 a_100_n29926# a_n100_n30023# a_n158_n29926# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X245 a_100_n77582# a_n100_n77679# a_n158_n77582# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X246 a_100_n40286# a_n100_n40383# a_n158_n40286# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X247 a_100_n38214# a_n100_n38311# a_n158_n38214# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X248 a_100_127546# a_n100_127449# a_n158_127546# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X249 a_100_n14386# a_n100_n14483# a_n158_n14386# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X250 a_100_57098# a_n100_57001# a_n158_57098# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X251 a_100_n108662# a_n100_n108759# a_n158_n108662# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X252 a_100_n130418# a_n100_n130515# a_n158_n130418# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X253 a_100_n73438# a_n100_n73535# a_n158_n73438# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X254 a_100_n95194# a_n100_n95291# a_n158_n95194# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X255 a_100_n47538# a_n100_n47635# a_n158_n47538# w_n358_n132787# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
C0 a_n100_n51779# a_n100_n50743# 0.205388f
C1 a_100_129618# a_n158_129618# 0.219309f
C2 a_n158_90250# a_n158_89214# 0.010536f
C3 a_n100_n64211# a_n100_n63175# 0.205388f
C4 a_100_n17494# a_100_n16458# 0.010536f
C5 a_n158_60206# a_n158_59170# 0.010536f
C6 a_n158_n101410# w_n358_n132787# 0.240254f
C7 a_n100_93261# a_n100_92225# 0.205388f
C8 a_100_18766# a_100_17730# 0.010536f
C9 a_n158_75746# w_n358_n132787# 0.240254f
C10 a_100_n110734# a_100_n111770# 0.010536f
C11 a_n100_n111867# a_n158_n111770# 0.090922f
C12 a_100_105790# a_100_104754# 0.010536f
C13 a_n158_n10242# a_n158_n11278# 0.010536f
C14 a_n100_34209# a_n100_33173# 0.205388f
C15 a_n158_n45466# a_100_n45466# 0.219309f
C16 a_100_96466# a_n100_96369# 0.090922f
C17 a_n158_n61006# w_n358_n132787# 0.240254f
C18 a_n158_118# w_n358_n132787# 0.240254f
C19 a_n100_n104615# a_n158_n104518# 0.090922f
C20 a_n100_n67319# a_n100_n66283# 0.205388f
C21 a_n158_n116950# a_100_n116950# 0.219309f
C22 a_n100_n117047# a_n100_n118083# 0.205388f
C23 a_100_n82762# a_n158_n82762# 0.219309f
C24 a_n100_n52815# a_100_n52718# 0.090922f
C25 a_100_23946# a_100_22910# 0.010536f
C26 a_n100_22813# a_n158_22910# 0.090922f
C27 a_n158_68494# w_n358_n132787# 0.240254f
C28 a_100_n46502# w_n358_n132787# 0.240254f
C29 a_100_116150# a_n158_116150# 0.219309f
C30 a_n100_51821# a_100_51918# 0.090922f
C31 a_n100_n40383# a_n100_n39347# 0.205388f
C32 a_n158_41558# a_100_41558# 0.219309f
C33 a_n100_49749# w_n358_n132787# 0.269531f
C34 a_100_124438# w_n358_n132787# 0.240254f
C35 a_100_59170# a_n100_59073# 0.090922f
C36 a_n158_62278# a_100_62278# 0.219309f
C37 a_100_n74474# a_n158_n74474# 0.219309f
C38 a_n158_70566# w_n358_n132787# 0.240254f
C39 a_n100_n48671# a_n100_n47635# 0.205388f
C40 a_100_31198# a_100_30162# 0.010536f
C41 a_n100_n8267# w_n358_n132787# 0.269531f
C42 a_100_57098# w_n358_n132787# 0.240254f
C43 a_n100_41461# w_n358_n132787# 0.269531f
C44 a_n158_n123166# a_100_n123166# 0.219309f
C45 a_n100_n123263# a_n100_n124299# 0.205388f
C46 a_n158_n84834# a_100_n84834# 0.219309f
C47 a_n158_19802# a_100_19802# 0.219309f
C48 a_n100_61145# w_n358_n132787# 0.269531f
C49 a_n100_42497# a_n158_42594# 0.090922f
C50 a_n158_n110734# w_n358_n132787# 0.240254f
C51 a_100_20838# w_n358_n132787# 0.240254f
C52 a_n100_n2051# a_n158_n1954# 0.090922f
C53 a_n100_n127407# a_100_n127310# 0.090922f
C54 a_n100_n73535# a_n100_n72499# 0.205388f
C55 a_100_61242# a_100_62278# 0.010536f
C56 a_n158_85070# a_n100_84973# 0.090922f
C57 a_n158_78854# a_n100_78757# 0.090922f
C58 a_100_n30962# w_n358_n132787# 0.240254f
C59 a_n100_11417# a_100_11514# 0.090922f
C60 a_100_n30962# a_100_n31998# 0.010536f
C61 a_n100_n30023# a_n158_n29926# 0.090922f
C62 a_n158_121330# a_n158_120294# 0.010536f
C63 a_n158_n127310# a_n158_n126274# 0.010536f
C64 a_n100_25921# a_100_26018# 0.090922f
C65 a_n100_n46599# w_n358_n132787# 0.269531f
C66 a_100_128582# a_100_129618# 0.010536f
C67 a_n158_4262# a_n158_3226# 0.010536f
C68 a_100_120294# w_n358_n132787# 0.240254f
C69 a_n158_n90014# a_n100_n90111# 0.090922f
C70 a_n158_n87942# a_n158_n86906# 0.010536f
C71 a_n100_16597# a_100_16694# 0.090922f
C72 a_100_89214# a_100_90250# 0.010536f
C73 a_n158_n71366# a_n158_n70330# 0.010536f
C74 a_n158_98538# a_100_98538# 0.219309f
C75 a_100_n66186# a_n158_n66186# 0.219309f
C76 a_n100_n57995# a_100_n57898# 0.090922f
C77 a_n158_58134# a_n158_59170# 0.010536f
C78 a_100_n73438# a_100_n74474# 0.010536f
C79 a_n100_n100471# w_n358_n132787# 0.269531f
C80 a_100_n35106# w_n358_n132787# 0.240254f
C81 a_n158_9442# a_n158_8406# 0.010536f
C82 a_n100_64253# w_n358_n132787# 0.269531f
C83 a_100_47774# w_n358_n132787# 0.240254f
C84 a_100_n129382# a_100_n130418# 0.010536f
C85 a_n100_n130515# a_n158_n130418# 0.090922f
C86 a_n158_90250# w_n358_n132787# 0.240254f
C87 a_100_n1954# w_n358_n132787# 0.240254f
C88 a_n100_n83895# a_n158_n83798# 0.090922f
C89 a_n100_n35203# a_n100_n34167# 0.205388f
C90 a_100_22910# a_100_21874# 0.010536f
C91 a_n158_n12314# w_n358_n132787# 0.240254f
C92 a_n100_110873# a_100_110970# 0.090922f
C93 a_n158_n108662# a_n158_n107626# 0.010536f
C94 a_n158_88178# a_n158_89214# 0.010536f
C95 a_n100_91189# a_100_91286# 0.090922f
C96 a_n100_95333# a_n100_94297# 0.205388f
C97 a_100_40522# a_100_39486# 0.010536f
C98 a_n100_39389# a_n158_39486# 0.090922f
C99 a_100_127546# a_100_128582# 0.010536f
C100 a_100_n100374# w_n358_n132787# 0.240254f
C101 a_n158_121330# a_100_121330# 0.219309f
C102 a_n158_125474# a_n158_126510# 0.010536f
C103 w_n358_n132787# a_100_n122130# 0.240254f
C104 a_n100_126413# a_n100_125377# 0.205388f
C105 a_100_n48574# a_100_n49610# 0.010536f
C106 a_n100_n18627# a_n100_n17591# 0.205388f
C107 a_100_n65150# a_n100_n65247# 0.090922f
C108 a_100_n72402# a_100_n71366# 0.010536f
C109 a_n100_38353# w_n358_n132787# 0.269531f
C110 a_n100_n39347# w_n358_n132787# 0.269531f
C111 a_100_80926# a_n100_80829# 0.090922f
C112 a_n158_65386# a_n100_65289# 0.090922f
C113 a_n158_n94158# a_100_n94158# 0.219309f
C114 a_100_63314# a_n100_63217# 0.090922f
C115 a_n100_18669# a_100_18766# 0.090922f
C116 a_n158_123402# a_n100_123305# 0.090922f
C117 a_100_58134# a_100_57098# 0.010536f
C118 a_n100_17633# w_n358_n132787# 0.269531f
C119 a_100_36378# a_100_35342# 0.010536f
C120 a_n100_122269# w_n358_n132787# 0.269531f
C121 a_100_52954# a_n100_52857# 0.090922f
C122 a_n158_n129382# w_n358_n132787# 0.240254f
C123 a_n100_n44527# a_100_n44430# 0.090922f
C124 a_n158_n7134# a_n158_n8170# 0.010536f
C125 a_n100_n35203# w_n358_n132787# 0.269531f
C126 a_100_n30962# a_100_n29926# 0.010536f
C127 a_n100_10381# a_100_10478# 0.090922f
C128 a_n100_n32095# a_n100_n33131# 0.205388f
C129 a_n100_117089# a_100_117186# 0.090922f
C130 a_100_52954# a_100_53990# 0.010536f
C131 a_n158_48810# a_n158_47774# 0.010536f
C132 a_100_n18530# a_100_n19566# 0.010536f
C133 a_n100_2093# a_n158_2190# 0.090922f
C134 a_100_n39250# a_n158_n39250# 0.219309f
C135 a_100_n82762# w_n358_n132787# 0.240254f
C136 a_100_43630# w_n358_n132787# 0.240254f
C137 a_n158_128582# a_n158_129618# 0.010536f
C138 a_100_n25782# a_100_n26818# 0.010536f
C139 a_n158_12550# w_n358_n132787# 0.240254f
C140 a_n158_66422# a_n158_65386# 0.010536f
C141 a_n100_125377# w_n358_n132787# 0.269531f
C142 a_100_78854# a_n100_78757# 0.090922f
C143 a_n100_n15519# a_n100_n14483# 0.205388f
C144 a_100_n47538# a_n158_n47538# 0.219309f
C145 a_100_123402# w_n358_n132787# 0.240254f
C146 a_100_n59970# w_n358_n132787# 0.240254f
C147 a_100_n34070# a_n158_n34070# 0.219309f
C148 a_n100_n120155# a_n158_n120058# 0.090922f
C149 a_n100_n23807# a_100_n23710# 0.090922f
C150 a_n100_20741# a_100_20838# 0.090922f
C151 a_100_91286# w_n358_n132787# 0.240254f
C152 a_100_n55826# a_100_n56862# 0.010536f
C153 a_n100_n53851# w_n358_n132787# 0.269531f
C154 a_100_n71366# a_100_n70330# 0.010536f
C155 a_n158_n93122# w_n358_n132787# 0.240254f
C156 a_n100_n106687# w_n358_n132787# 0.269531f
C157 a_n100_n27951# w_n358_n132787# 0.269531f
C158 a_100_72638# a_n100_72541# 0.090922f
C159 a_100_94394# w_n358_n132787# 0.240254f
C160 a_n158_58134# a_n100_58037# 0.090922f
C161 a_n158_92322# a_n158_91286# 0.010536f
C162 a_n100_n49707# a_100_n49610# 0.090922f
C163 a_n158_28090# a_n158_27054# 0.010536f
C164 a_100_n43394# w_n358_n132787# 0.240254f
C165 a_100_n17494# a_n158_n17494# 0.219309f
C166 a_100_n68258# a_n100_n68355# 0.090922f
C167 a_100_87142# w_n358_n132787# 0.240254f
C168 a_100_36378# w_n358_n132787# 0.240254f
C169 a_n158_5298# a_n158_4262# 0.010536f
C170 a_n100_n119119# w_n358_n132787# 0.269531f
C171 a_n100_46641# a_n158_46738# 0.090922f
C172 a_n158_n91050# w_n358_n132787# 0.240254f
C173 a_n158_17730# a_100_17730# 0.219309f
C174 a_n158_88178# w_n358_n132787# 0.240254f
C175 a_n158_96466# a_n100_96369# 0.090922f
C176 a_n100_n81823# a_100_n81726# 0.090922f
C177 a_n158_101646# a_n158_102682# 0.010536f
C178 a_n158_15658# w_n358_n132787# 0.240254f
C179 a_n100_76685# w_n358_n132787# 0.269531f
C180 a_n158_109934# a_100_109934# 0.219309f
C181 a_n158_n109698# w_n358_n132787# 0.240254f
C182 a_100_62278# w_n358_n132787# 0.240254f
C183 a_n158_n30962# a_n100_n31059# 0.090922f
C184 a_n100_n1015# w_n358_n132787# 0.269531f
C185 a_n100_n9303# w_n358_n132787# 0.269531f
C186 a_n158_59170# w_n358_n132787# 0.240254f
C187 a_n158_57098# a_n158_56062# 0.010536f
C188 w_n358_n132787# a_100_n71366# 0.240254f
C189 a_n158_n73438# a_n100_n73535# 0.090922f
C190 a_100_n50646# w_n358_n132787# 0.240254f
C191 a_n100_72541# w_n358_n132787# 0.269531f
C192 a_100_n126274# a_n100_n126371# 0.090922f
C193 a_100_n106590# w_n358_n132787# 0.240254f
C194 a_n100_n24843# w_n358_n132787# 0.269531f
C195 a_n158_116150# w_n358_n132787# 0.240254f
C196 a_n100_14525# a_n100_13489# 0.205388f
C197 a_n100_n89075# w_n358_n132787# 0.269531f
C198 a_100_108898# a_100_109934# 0.010536f
C199 a_n158_128582# a_100_128582# 0.219309f
C200 a_n158_n62042# w_n358_n132787# 0.240254f
C201 a_n158_30162# a_100_30162# 0.219309f
C202 a_100_n61006# a_n158_n61006# 0.219309f
C203 a_n158_n87942# a_n100_n88039# 0.090922f
C204 a_100_81962# a_n158_81962# 0.219309f
C205 a_n158_56062# a_n158_55026# 0.010536f
C206 a_n158_n125238# a_n158_n126274# 0.010536f
C207 a_n158_n5062# w_n358_n132787# 0.240254f
C208 a_n100_n16555# w_n358_n132787# 0.269531f
C209 a_n100_n91147# w_n358_n132787# 0.269531f
C210 a_100_n109698# a_100_n110734# 0.010536f
C211 a_n100_n110831# a_n158_n110734# 0.090922f
C212 a_100_n56862# w_n358_n132787# 0.240254f
C213 a_100_n20602# a_100_n21638# 0.010536f
C214 a_n100_n2051# a_n100_n3087# 0.205388f
C215 a_n100_19705# w_n358_n132787# 0.269531f
C216 a_100_127546# a_n158_127546# 0.219309f
C217 a_n100_90153# a_100_90250# 0.090922f
C218 a_n100_101549# a_n100_100513# 0.205388f
C219 a_n100_n104615# w_n358_n132787# 0.269531f
C220 a_100_n62042# w_n358_n132787# 0.240254f
C221 a_n158_72638# a_100_72638# 0.219309f
C222 a_n100_n98399# a_100_n98302# 0.090922f
C223 a_n100_n104615# a_n100_n103579# 0.205388f
C224 a_n100_n17591# a_n158_n17494# 0.090922f
C225 a_n100_50785# w_n358_n132787# 0.269531f
C226 a_n158_26018# a_100_26018# 0.219309f
C227 w_n358_n132787# a_100_n121094# 0.240254f
C228 a_n158_99574# a_n100_99477# 0.090922f
C229 a_n100_53893# w_n358_n132787# 0.269531f
C230 a_n100_n24843# a_n100_n25879# 0.205388f
C231 a_n158_100610# w_n358_n132787# 0.240254f
C232 a_n158_n26818# a_n158_n25782# 0.010536f
C233 a_n100_n106687# a_n158_n106590# 0.090922f
C234 a_n158_n79654# a_n100_n79751# 0.090922f
C235 a_n158_16694# a_100_16694# 0.219309f
C236 a_n100_16597# a_n100_15561# 0.205388f
C237 a_n158_116150# a_n100_116053# 0.090922f
C238 a_n158_n113842# a_100_n113842# 0.219309f
C239 a_n100_n113939# a_n100_n114975# 0.205388f
C240 a_n158_n4026# a_n158_n5062# 0.010536f
C241 a_100_115114# a_n158_115114# 0.219309f
C242 a_n158_62278# a_n158_63314# 0.010536f
C243 a_n100_121233# w_n358_n132787# 0.269531f
C244 a_n158_48810# a_n158_49846# 0.010536f
C245 a_n158_n132490# a_100_n132490# 0.219309f
C246 a_n158_n36142# w_n358_n132787# 0.240254f
C247 a_n100_8309# a_n158_8406# 0.090922f
C248 a_n100_55965# a_n100_54929# 0.205388f
C249 a_100_n81726# a_n158_n81726# 0.219309f
C250 a_n100_n33131# a_n158_n33034# 0.090922f
C251 a_n158_94394# w_n358_n132787# 0.240254f
C252 a_n158_n128346# w_n358_n132787# 0.240254f
C253 a_n100_21777# a_n158_21874# 0.090922f
C254 a_100_74710# w_n358_n132787# 0.240254f
C255 a_n100_77721# w_n358_n132787# 0.269531f
C256 a_100_24982# w_n358_n132787# 0.240254f
C257 a_n100_21# a_n158_118# 0.090922f
C258 a_n100_39389# a_100_39486# 0.090922f
C259 a_n158_n8170# a_100_n8170# 0.219309f
C260 a_n100_122269# a_n158_122366# 0.090922f
C261 a_n158_85070# w_n358_n132787# 0.240254f
C262 a_n158_72638# w_n358_n132787# 0.240254f
C263 a_100_115114# a_n100_115017# 0.090922f
C264 a_100_n64114# a_n100_n64211# 0.090922f
C265 a_n100_n116011# a_n100_n114975# 0.205388f
C266 a_n158_117186# a_100_117186# 0.219309f
C267 a_100_n42358# w_n358_n132787# 0.240254f
C268 a_n158_6334# a_n158_5298# 0.010536f
C269 a_n100_n78715# a_n100_n77679# 0.205388f
C270 a_100_92322# a_100_91286# 0.010536f
C271 a_n100_58037# w_n358_n132787# 0.269531f
C272 a_n100_n66283# w_n358_n132787# 0.269531f
C273 a_100_n103482# w_n358_n132787# 0.240254f
C274 a_n158_18766# a_100_18766# 0.219309f
C275 a_100_n103482# a_n100_n103579# 0.090922f
C276 a_n158_n59970# w_n358_n132787# 0.240254f
C277 a_n158_n78618# a_100_n78618# 0.219309f
C278 a_100_n105554# w_n358_n132787# 0.240254f
C279 a_100_n106590# a_n158_n106590# 0.219309f
C280 a_100_117186# a_100_118222# 0.010536f
C281 a_n100_35245# a_100_35342# 0.090922f
C282 a_n158_n35106# w_n358_n132787# 0.240254f
C283 a_n100_120197# w_n358_n132787# 0.269531f
C284 a_n100_10381# a_n100_9345# 0.205388f
C285 a_n158_n115914# a_100_n115914# 0.219309f
C286 a_n100_n116011# a_n100_n117047# 0.205388f
C287 a_n100_n98399# a_n158_n98302# 0.090922f
C288 a_100_n83798# w_n358_n132787# 0.240254f
C289 a_100_50882# w_n358_n132787# 0.240254f
C290 a_n100_n19663# a_100_n19566# 0.090922f
C291 a_n158_45702# a_n158_46738# 0.010536f
C292 a_n100_30065# w_n358_n132787# 0.269531f
C293 a_100_n37178# a_100_n38214# 0.010536f
C294 a_n158_n40286# a_n158_n39250# 0.010536f
C295 a_100_65386# w_n358_n132787# 0.240254f
C296 a_n158_119258# a_n158_118222# 0.010536f
C297 a_100_n84834# w_n358_n132787# 0.240254f
C298 a_n100_42497# w_n358_n132787# 0.269531f
C299 a_n100_n77679# w_n358_n132787# 0.269531f
C300 a_n100_n10339# a_n158_n10242# 0.090922f
C301 a_100_59170# a_n158_59170# 0.219309f
C302 a_n100_14525# a_n158_14622# 0.090922f
C303 a_n100_n118083# w_n358_n132787# 0.269531f
C304 a_n100_11417# w_n358_n132787# 0.269531f
C305 a_100_n45466# a_100_n46502# 0.010536f
C306 a_100_n69294# a_n158_n69294# 0.219309f
C307 a_n100_n70427# a_n100_n69391# 0.205388f
C308 a_n158_n13350# a_100_n13350# 0.219309f
C309 a_n158_57098# a_n158_58134# 0.010536f
C310 a_n158_n122130# a_100_n122130# 0.219309f
C311 a_n100_n122227# a_n100_n123263# 0.205388f
C312 a_n100_20741# a_n100_19705# 0.205388f
C313 a_n158_n94158# w_n358_n132787# 0.240254f
C314 a_n100_130557# a_n158_130654# 0.090922f
C315 a_n100_n119119# a_100_n119022# 0.090922f
C316 a_100_120294# a_n158_120294# 0.219309f
C317 a_100_38450# a_100_37414# 0.010536f
C318 a_n158_108898# w_n358_n132787# 0.240254f
C319 a_n158_n43394# a_n158_n44430# 0.010536f
C320 a_100_13586# a_100_12550# 0.010536f
C321 a_n158_80926# w_n358_n132787# 0.240254f
C322 a_100_n97266# a_n158_n97266# 0.219309f
C323 a_100_n59970# a_100_n61006# 0.010536f
C324 a_100_72638# a_100_73674# 0.010536f
C325 a_100_6334# w_n358_n132787# 0.240254f
C326 a_n100_124341# a_n158_124438# 0.090922f
C327 a_n158_n77582# a_n100_n77679# 0.090922f
C328 a_n158_n51682# a_n158_n50646# 0.010536f
C329 a_n158_128582# a_n158_127546# 0.010536f
C330 a_n100_26957# a_n158_27054# 0.090922f
C331 a_n100_n51779# a_100_n51682# 0.090922f
C332 a_n100_n49707# a_n100_n50743# 0.205388f
C333 a_n158_98538# w_n358_n132787# 0.240254f
C334 a_100_n17494# a_100_n18530# 0.010536f
C335 a_n100_n44527# w_n358_n132787# 0.269531f
C336 a_n100_75649# w_n358_n132787# 0.269531f
C337 a_n158_82998# a_100_82998# 0.219309f
C338 a_n100_35245# w_n358_n132787# 0.269531f
C339 a_100_75746# w_n358_n132787# 0.240254f
C340 a_n100_46641# a_100_46738# 0.090922f
C341 a_n158_77818# w_n358_n132787# 0.240254f
C342 a_n158_n57898# w_n358_n132787# 0.240254f
C343 a_n100_n125335# a_100_n125238# 0.090922f
C344 a_100_15658# w_n358_n132787# 0.240254f
C345 a_n158_34306# a_n158_33270# 0.010536f
C346 a_100_n128346# a_100_n129382# 0.010536f
C347 a_n100_n129479# a_n158_n129382# 0.090922f
C348 a_100_58134# a_n100_58037# 0.090922f
C349 a_100_120294# a_100_121330# 0.010536f
C350 a_n158_n918# w_n358_n132787# 0.240254f
C351 a_n158_n9206# w_n358_n132787# 0.240254f
C352 a_n158_n105554# a_n100_n105651# 0.090922f
C353 a_100_n6098# a_n158_n6098# 0.219309f
C354 a_n158_22910# a_100_22910# 0.219309f
C355 a_100_n97266# w_n358_n132787# 0.240254f
C356 w_n358_n132787# a_n158_n107626# 0.240254f
C357 a_100_28090# w_n358_n132787# 0.240254f
C358 a_n158_n38214# a_100_n38214# 0.219309f
C359 a_n100_73577# a_n100_72541# 0.205388f
C360 a_100_119258# w_n358_n132787# 0.240254f
C361 a_n100_n85967# w_n358_n132787# 0.269531f
C362 a_100_n71366# a_n100_n71463# 0.090922f
C363 a_100_73674# w_n358_n132787# 0.240254f
C364 a_n100_81865# w_n358_n132787# 0.269531f
C365 a_100_97502# a_n158_97502# 0.219309f
C366 w_n358_n132787# a_100_n120058# 0.240254f
C367 a_100_n58934# a_100_n59970# 0.010536f
C368 a_n100_n43491# w_n358_n132787# 0.269531f
C369 a_n100_n81823# a_n158_n81726# 0.090922f
C370 a_n158_106826# a_n158_107862# 0.010536f
C371 a_100_n103482# a_100_n102446# 0.010536f
C372 a_n100_47677# a_n158_47774# 0.090922f
C373 a_n158_n94158# a_n100_n94255# 0.090922f
C374 a_n100_67361# a_n158_67458# 0.090922f
C375 a_n100_n56959# a_n100_n57995# 0.205388f
C376 a_n100_97405# w_n358_n132787# 0.269531f
C377 a_n100_n21735# a_100_n21638# 0.090922f
C378 a_n100_n23807# a_n100_n24843# 0.205388f
C379 a_n158_n127310# w_n358_n132787# 0.240254f
C380 a_n100_36281# a_100_36378# 0.090922f
C381 a_n158_123402# w_n358_n132787# 0.240254f
C382 a_100_57098# a_100_56062# 0.010536f
C383 a_n158_63314# w_n358_n132787# 0.240254f
C384 a_n100_n32095# w_n358_n132787# 0.269531f
C385 a_n100_n32095# a_100_n31998# 0.090922f
C386 a_n158_93358# a_n158_92322# 0.010536f
C387 a_n100_119161# a_n100_120197# 0.205388f
C388 a_n100_3129# w_n358_n132787# 0.269531f
C389 a_n158_n49610# a_100_n49610# 0.219309f
C390 w_n358_n132787# a_n158_n126274# 0.240254f
C391 a_n100_3129# a_100_3226# 0.090922f
C392 a_n158_n65150# a_n158_n64114# 0.010536f
C393 a_100_n20602# w_n358_n132787# 0.240254f
C394 a_100_94394# a_n100_94297# 0.090922f
C395 a_n100_n26915# a_n100_n27951# 0.205388f
C396 a_100_n62042# a_100_n61006# 0.010536f
C397 a_100_n36142# w_n358_n132787# 0.240254f
C398 a_n158_n15422# a_n158_n14386# 0.010536f
C399 a_n158_50882# a_n100_50785# 0.090922f
C400 a_n100_n33131# a_n100_n34167# 0.205388f
C401 a_n100_n114975# w_n358_n132787# 0.269531f
C402 a_n100_62181# a_n100_63217# 0.205388f
C403 a_100_n97266# a_100_n96230# 0.010536f
C404 a_n158_n2990# w_n358_n132787# 0.240254f
C405 a_n158_69530# a_n158_68494# 0.010536f
C406 a_n100_21777# a_100_21874# 0.090922f
C407 a_n158_n80690# a_100_n80690# 0.219309f
C408 a_n158_n50646# w_n358_n132787# 0.240254f
C409 a_n100_n74571# a_n158_n74474# 0.090922f
C410 a_n100_51821# a_n100_52857# 0.205388f
C411 a_n100_21# a_n100_n1015# 0.205388f
C412 a_n158_112006# a_100_112006# 0.219309f
C413 a_100_n5062# w_n358_n132787# 0.240254f
C414 a_n158_57098# w_n358_n132787# 0.240254f
C415 a_100_n95194# a_n100_n95291# 0.090922f
C416 a_100_n24746# w_n358_n132787# 0.240254f
C417 a_n100_13489# a_n158_13586# 0.090922f
C418 a_n100_129521# w_n358_n132787# 0.269531f
C419 a_n158_69530# a_n158_70566# 0.010536f
C420 a_n158_29126# a_n158_28090# 0.010536f
C421 a_n100_n16555# a_100_n16458# 0.090922f
C422 a_n100_n117047# w_n358_n132787# 0.269531f
C423 a_n100_n95291# w_n358_n132787# 0.269531f
C424 a_100_109934# a_n100_109837# 0.090922f
C425 a_n100_115017# a_n100_113981# 0.205388f
C426 a_n100_n81823# a_n100_n82859# 0.205388f
C427 a_n100_n99435# a_n100_n100471# 0.205388f
C428 a_n158_n106590# a_n158_n107626# 0.010536f
C429 a_n100_123305# w_n358_n132787# 0.269531f
C430 a_n158_55026# w_n358_n132787# 0.240254f
C431 a_n158_18766# a_n158_17730# 0.010536f
C432 a_n100_n8267# a_100_n8170# 0.090922f
C433 a_n158_n2990# a_n158_n4026# 0.010536f
C434 w_n358_n132787# a_n100_n69391# 0.269531f
C435 a_n158_n108662# w_n358_n132787# 0.240254f
C436 a_n100_n33131# w_n358_n132787# 0.269531f
C437 a_n158_n117986# a_n158_n119022# 0.010536f
C438 a_n100_110873# a_n100_111909# 0.205388f
C439 a_n158_110970# w_n358_n132787# 0.240254f
C440 a_100_98538# w_n358_n132787# 0.240254f
C441 a_n100_23849# a_100_23946# 0.090922f
C442 a_n158_113042# a_n158_112006# 0.010536f
C443 a_n158_84034# a_n158_85070# 0.010536f
C444 a_n100_108801# a_n158_108898# 0.090922f
C445 a_n100_n67319# w_n358_n132787# 0.269531f
C446 a_n100_n38311# a_100_n38214# 0.090922f
C447 a_n158_n84834# w_n358_n132787# 0.240254f
C448 a_n100_14525# a_100_14622# 0.090922f
C449 a_n158_42594# w_n358_n132787# 0.240254f
C450 a_n100_119161# a_100_119258# 0.090922f
C451 a_100_127546# a_n100_127449# 0.090922f
C452 a_n100_n67319# a_100_n67222# 0.090922f
C453 a_100_11514# w_n358_n132787# 0.240254f
C454 a_n100_31101# a_n158_31198# 0.090922f
C455 a_n100_70469# w_n358_n132787# 0.269531f
C456 a_n158_50882# a_100_50882# 0.219309f
C457 a_n158_n124202# a_n158_n125238# 0.010536f
C458 a_n100_101549# a_100_101646# 0.090922f
C459 a_100_86106# w_n358_n132787# 0.240254f
C460 a_100_n101410# a_n100_n101507# 0.090922f
C461 a_n158_n13350# w_n358_n132787# 0.240254f
C462 a_n158_20838# a_100_20838# 0.219309f
C463 a_n158_56062# w_n358_n132787# 0.240254f
C464 a_n100_n54887# w_n358_n132787# 0.269531f
C465 a_n100_43533# a_100_43630# 0.090922f
C466 a_n100_37317# a_100_37414# 0.090922f
C467 a_100_n72402# a_n158_n72402# 0.219309f
C468 a_100_n42358# a_n100_n42455# 0.090922f
C469 a_n100_12453# a_n158_12550# 0.090922f
C470 a_100_48810# a_100_49846# 0.010536f
C471 a_100_n87942# w_n358_n132787# 0.240254f
C472 a_n158_94394# a_n100_94297# 0.090922f
C473 a_n158_n64114# w_n358_n132787# 0.240254f
C474 a_100_n95194# a_100_n94158# 0.010536f
C475 a_n100_5201# w_n358_n132787# 0.269531f
C476 a_100_n84834# a_100_n85870# 0.010536f
C477 a_n100_26957# a_100_27054# 0.090922f
C478 a_100_n44430# w_n358_n132787# 0.240254f
C479 a_100_5298# a_100_4262# 0.010536f
C480 a_n158_46738# a_100_46738# 0.219309f
C481 a_n100_46641# a_n100_45605# 0.205388f
C482 a_n100_n95291# a_n100_n94255# 0.205388f
C483 a_n158_17730# a_n158_16694# 0.010536f
C484 a_100_n94158# w_n358_n132787# 0.240254f
C485 a_n158_n19566# w_n358_n132787# 0.240254f
C486 a_n100_n59031# w_n358_n132787# 0.269531f
C487 a_n158_n80690# w_n358_n132787# 0.240254f
C488 a_n158_n112806# a_100_n112806# 0.219309f
C489 a_n100_n112903# a_n100_n113939# 0.205388f
C490 a_n100_84973# w_n358_n132787# 0.269531f
C491 a_n158_n131454# a_100_n131454# 0.219309f
C492 a_n100_n131551# a_n100_n132587# 0.205388f
C493 a_n158_117186# a_n158_118222# 0.010536f
C494 a_100_130654# a_100_131690# 0.010536f
C495 a_n158_n104518# w_n358_n132787# 0.240254f
C496 a_100_10478# a_100_9442# 0.010536f
C497 a_n158_n33034# w_n358_n132787# 0.240254f
C498 a_100_n119022# a_100_n120058# 0.010536f
C499 a_100_n10242# w_n358_n132787# 0.240254f
C500 a_n158_106826# a_100_106826# 0.219309f
C501 a_n100_79793# a_100_79890# 0.090922f
C502 a_n158_118222# a_100_118222# 0.219309f
C503 a_100_84034# w_n358_n132787# 0.240254f
C504 a_100_41558# a_100_40522# 0.010536f
C505 a_n100_40425# a_n158_40522# 0.090922f
C506 a_n158_106826# a_n158_105790# 0.010536f
C507 a_n158_123402# a_n158_122366# 0.010536f
C508 a_n100_121233# a_100_121330# 0.090922f
C509 a_100_n21638# w_n358_n132787# 0.240254f
C510 a_n100_73577# a_100_73674# 0.090922f
C511 a_n100_n75607# w_n358_n132787# 0.269531f
C512 a_n158_14622# a_n158_13586# 0.010536f
C513 w_n358_n132787# a_n158_n125238# 0.240254f
C514 a_100_n99338# a_100_n98302# 0.010536f
C515 a_n158_60206# w_n358_n132787# 0.240254f
C516 a_n158_79890# a_n158_80926# 0.010536f
C517 a_n100_n107723# a_100_n107626# 0.090922f
C518 a_n158_30162# a_n158_29126# 0.010536f
C519 a_n100_78757# a_n100_77721# 0.205388f
C520 a_n100_95333# a_n158_95430# 0.090922f
C521 a_n100_120197# a_n158_120294# 0.090922f
C522 a_n100_40425# w_n358_n132787# 0.269531f
C523 a_100_89214# a_n100_89117# 0.090922f
C524 a_100_7370# a_100_6334# 0.010536f
C525 a_n158_n102446# w_n358_n132787# 0.240254f
C526 a_n100_n70427# a_100_n70330# 0.090922f
C527 a_n158_47774# a_100_47774# 0.219309f
C528 a_n100_n54887# a_100_n54790# 0.090922f
C529 a_100_n13350# w_n358_n132787# 0.240254f
C530 a_n100_n113939# w_n358_n132787# 0.269531f
C531 a_n158_n54790# a_n158_n55826# 0.010536f
C532 a_100_116150# w_n358_n132787# 0.240254f
C533 a_100_114078# w_n358_n132787# 0.240254f
C534 a_n158_19802# a_n158_18766# 0.010536f
C535 a_n100_n132587# w_n358_n132787# 0.349164f
C536 a_100_n22674# a_100_n21638# 0.010536f
C537 a_n158_n1954# a_100_n1954# 0.219309f
C538 a_100_n90014# a_100_n91050# 0.010536f
C539 a_n100_n12411# a_100_n12314# 0.090922f
C540 a_n100_36281# a_n100_35245# 0.205388f
C541 a_100_69530# w_n358_n132787# 0.240254f
C542 a_n158_n75510# a_n100_n75607# 0.090922f
C543 a_n158_113042# a_n158_114078# 0.010536f
C544 a_100_n30962# a_n158_n30962# 0.219309f
C545 a_100_43630# a_100_42594# 0.010536f
C546 a_n100_n85967# a_100_n85870# 0.090922f
C547 a_n158_32234# w_n358_n132787# 0.240254f
C548 a_n100_3129# a_n100_2093# 0.205388f
C549 a_n158_104754# w_n358_n132787# 0.240254f
C550 a_100_45702# w_n358_n132787# 0.240254f
C551 a_n100_n7231# a_n100_n6195# 0.205388f
C552 a_n100_n94255# a_100_n94158# 0.090922f
C553 a_n100_n21735# w_n358_n132787# 0.269531f
C554 a_100_64350# a_100_63314# 0.010536f
C555 a_n158_62278# w_n358_n132787# 0.240254f
C556 a_n100_n116011# w_n358_n132787# 0.269531f
C557 a_n100_n5159# a_n158_n5062# 0.090922f
C558 a_100_87142# a_n158_87142# 0.219309f
C559 a_100_76782# a_n158_76782# 0.219309f
C560 a_100_101646# a_n158_101646# 0.219309f
C561 a_100_55026# a_n158_55026# 0.219309f
C562 a_100_102682# w_n358_n132787# 0.240254f
C563 a_100_n47538# a_100_n48574# 0.010536f
C564 a_n158_n72402# w_n358_n132787# 0.240254f
C565 a_n100_n13447# a_n100_n14483# 0.205388f
C566 a_n100_n37275# w_n358_n132787# 0.269531f
C567 a_n158_87142# a_n158_88178# 0.010536f
C568 w_n358_n132787# a_n100_n70427# 0.269531f
C569 a_100_9442# a_100_8406# 0.010536f
C570 a_n158_n35106# a_n158_n34070# 0.010536f
C571 a_n158_n121094# a_100_n121094# 0.219309f
C572 a_n100_n121191# a_n100_n122227# 0.205388f
C573 a_n100_n4123# w_n358_n132787# 0.269531f
C574 a_100_61242# w_n358_n132787# 0.240254f
C575 a_n158_21874# a_100_21874# 0.219309f
C576 w_n358_n132787# a_100_131690# 0.244798f
C577 a_n100_131593# a_n158_131690# 0.090922f
C578 a_n158_23946# w_n358_n132787# 0.240254f
C579 a_100_116150# a_n100_116053# 0.090922f
C580 a_n100_n118083# a_100_n117986# 0.090922f
C581 a_n100_n85967# a_n158_n85870# 0.090922f
C582 a_n100_n43491# a_n100_n42455# 0.205388f
C583 a_n158_118# a_100_118# 0.219309f
C584 a_n100_107765# a_100_107862# 0.090922f
C585 a_100_100610# a_100_99574# 0.010536f
C586 a_n158_n100374# w_n358_n132787# 0.240254f
C587 a_n100_13489# a_100_13586# 0.090922f
C588 a_100_n27854# a_100_n28890# 0.010536f
C589 a_100_125474# a_100_124438# 0.010536f
C590 a_n100_129521# a_n100_128485# 0.205388f
C591 a_n158_58134# w_n358_n132787# 0.240254f
C592 a_n158_37414# w_n358_n132787# 0.240254f
C593 a_n158_n82762# w_n358_n132787# 0.240254f
C594 a_n100_49749# a_n158_49846# 0.090922f
C595 a_n100_n124299# a_100_n124202# 0.090922f
C596 a_n158_n23710# a_n158_n24746# 0.010536f
C597 a_100_n109698# a_100_n108662# 0.010536f
C598 a_n158_n109698# a_n100_n109795# 0.090922f
C599 a_n100_n4123# a_n158_n4026# 0.090922f
C600 a_n158_n44430# a_n158_n45466# 0.010536f
C601 a_100_n127310# a_100_n128346# 0.010536f
C602 a_n100_n128443# a_n158_n128346# 0.090922f
C603 a_100_n4026# a_100_n5062# 0.010536f
C604 a_n100_1057# w_n358_n132787# 0.269531f
C605 a_n158_n65150# w_n358_n132787# 0.240254f
C606 a_n158_n51682# w_n358_n132787# 0.240254f
C607 a_n100_n38311# a_n100_n39347# 0.205388f
C608 a_n158_2190# a_100_2190# 0.219309f
C609 a_100_n72402# w_n358_n132787# 0.240254f
C610 a_100_n80690# w_n358_n132787# 0.240254f
C611 a_n158_45702# a_n100_45605# 0.090922f
C612 a_n158_89214# w_n358_n132787# 0.240254f
C613 a_n158_14622# a_100_14622# 0.219309f
C614 a_n158_n102446# a_100_n102446# 0.219309f
C615 a_n100_n85967# a_n100_n87003# 0.205388f
C616 a_n158_n24746# a_n158_n25782# 0.010536f
C617 a_n100_n46599# a_n100_n47635# 0.205388f
C618 a_100_60206# a_n100_60109# 0.090922f
C619 a_n100_n6195# w_n358_n132787# 0.269531f
C620 a_n100_31101# a_100_31198# 0.090922f
C621 a_n100_n40383# w_n358_n132787# 0.269531f
C622 a_n100_104657# a_n158_104754# 0.090922f
C623 a_n158_85070# a_100_85070# 0.219309f
C624 a_n100_95333# a_100_95430# 0.090922f
C625 a_100_93358# a_n100_93261# 0.090922f
C626 a_n158_99574# a_100_99574# 0.219309f
C627 a_n100_n7231# w_n358_n132787# 0.269531f
C628 a_100_n63078# a_100_n62042# 0.010536f
C629 a_100_102682# a_100_103718# 0.010536f
C630 a_n158_80926# a_100_80926# 0.219309f
C631 a_100_67458# w_n358_n132787# 0.240254f
C632 a_n158_43630# a_100_43630# 0.219309f
C633 a_n100_43533# a_n100_42497# 0.205388f
C634 a_100_130654# w_n358_n132787# 0.240254f
C635 a_100_n55826# w_n358_n132787# 0.240254f
C636 a_n100_99477# a_100_99574# 0.090922f
C637 a_n158_n83798# a_100_n83798# 0.219309f
C638 a_100_n42358# a_n158_n42358# 0.219309f
C639 a_n158_70566# a_n158_71602# 0.010536f
C640 a_n100_n89075# a_n100_n90111# 0.205388f
C641 a_n100_n11375# a_n158_n11278# 0.090922f
C642 a_n100_100513# a_n158_100610# 0.090922f
C643 a_n100_98441# a_n100_99477# 0.205388f
C644 a_n100_91189# w_n358_n132787# 0.269531f
C645 a_n100_12453# a_n100_11417# 0.205388f
C646 a_n158_93358# a_100_93358# 0.219309f
C647 a_n100_n51779# a_n100_n52815# 0.205388f
C648 a_n158_27054# a_100_27054# 0.219309f
C649 w_n358_n132787# a_n158_n124202# 0.240254f
C650 a_100_n50646# a_100_n49610# 0.010536f
C651 a_n158_51918# a_n158_52954# 0.010536f
C652 a_n158_76782# a_n158_75746# 0.010536f
C653 a_100_35342# w_n358_n132787# 0.240254f
C654 a_n100_n80787# a_n100_n79751# 0.205388f
C655 a_n158_52954# w_n358_n132787# 0.240254f
C656 a_n100_84973# a_n100_83937# 0.205388f
C657 a_n100_n83895# a_n100_n84931# 0.205388f
C658 a_n100_n91147# a_n100_n90111# 0.205388f
C659 a_n158_n99338# a_n158_n100374# 0.010536f
C660 a_100_58134# a_n158_58134# 0.219309f
C661 a_n100_126413# w_n358_n132787# 0.269531f
C662 a_n100_n112903# w_n358_n132787# 0.269531f
C663 a_100_34306# a_100_33270# 0.010536f
C664 a_n100_9345# a_100_9442# 0.090922f
C665 a_100_72638# w_n358_n132787# 0.240254f
C666 a_n100_n34167# w_n358_n132787# 0.269531f
C667 a_n100_n131551# w_n358_n132787# 0.269531f
C668 w_n358_n132787# a_100_n70330# 0.240254f
C669 a_n100_112945# w_n358_n132787# 0.269531f
C670 a_100_84034# a_n100_83937# 0.090922f
C671 a_n158_n97266# w_n358_n132787# 0.240254f
C672 a_n100_n20699# a_100_n20602# 0.090922f
C673 a_100_n90014# a_n158_n90014# 0.219309f
C674 a_n100_1057# a_100_1154# 0.090922f
C675 a_n100_90153# a_n100_89117# 0.205388f
C676 a_100_105790# a_100_106826# 0.010536f
C677 a_n158_n84834# a_n158_n85870# 0.010536f
C678 a_n100_n78715# w_n358_n132787# 0.269531f
C679 a_n158_n40286# a_n158_n41322# 0.010536f
C680 a_100_105790# a_n158_105790# 0.219309f
C681 a_n100_105693# w_n358_n132787# 0.269531f
C682 a_n158_90250# a_100_90250# 0.219309f
C683 a_n100_n102543# a_n158_n102446# 0.090922f
C684 a_100_125474# a_n100_125377# 0.090922f
C685 a_n158_40522# w_n358_n132787# 0.240254f
C686 a_100_n95194# w_n358_n132787# 0.240254f
C687 a_n100_6237# a_100_6334# 0.090922f
C688 a_n158_109934# a_n100_109837# 0.090922f
C689 a_n100_n105651# a_n100_n106687# 0.205388f
C690 a_n100_n111867# a_n100_n112903# 0.205388f
C691 a_100_n55826# a_100_n54790# 0.010536f
C692 a_n100_69433# a_n100_68397# 0.205388f
C693 a_n158_51918# w_n358_n132787# 0.240254f
C694 a_n158_36378# a_100_36378# 0.219309f
C695 a_n158_n12314# a_100_n12314# 0.219309f
C696 a_100_n31998# w_n358_n132787# 0.240254f
C697 a_100_n68258# a_100_n69294# 0.010536f
C698 a_n158_n116950# a_n158_n117986# 0.010536f
C699 a_n158_n66186# a_n100_n66283# 0.090922f
C700 a_n100_n103579# w_n358_n132787# 0.269531f
C701 a_n100_71505# a_n100_72541# 0.205388f
C702 a_100_3226# w_n358_n132787# 0.240254f
C703 a_100_53990# a_n158_53990# 0.219309f
C704 a_n100_64253# a_n100_65289# 0.205388f
C705 a_n100_42497# a_100_42594# 0.090922f
C706 a_100_n67222# w_n358_n132787# 0.240254f
C707 a_n158_93358# a_n100_93261# 0.090922f
C708 a_n100_n62139# a_n100_n61103# 0.205388f
C709 a_n158_84034# a_100_84034# 0.219309f
C710 a_n100_24885# a_100_24982# 0.090922f
C711 a_n158_n48574# w_n358_n132787# 0.240254f
C712 a_100_126510# a_n100_126413# 0.090922f
C713 a_100_n58934# a_n100_n59031# 0.090922f
C714 a_100_n22674# w_n358_n132787# 0.240254f
C715 a_n158_44666# w_n358_n132787# 0.240254f
C716 a_100_16694# a_100_15658# 0.010536f
C717 a_n100_15561# a_n158_15658# 0.090922f
C718 a_n100_47677# a_n100_46641# 0.205388f
C719 a_n158_32234# a_100_32234# 0.219309f
C720 a_n158_n75510# w_n358_n132787# 0.240254f
C721 a_n100_n48671# a_100_n48574# 0.090922f
C722 a_n100_n15519# a_n100_n16555# 0.205388f
C723 a_n158_n123166# a_n158_n124202# 0.010536f
C724 a_100_n14386# a_100_n13350# 0.010536f
C725 a_n158_8406# a_100_8406# 0.219309f
C726 a_n158_n77582# w_n358_n132787# 0.240254f
C727 a_n100_n35203# a_n100_n36239# 0.205388f
C728 a_n158_n4026# w_n358_n132787# 0.240254f
C729 a_100_71602# a_100_72638# 0.010536f
C730 a_n100_n111867# w_n358_n132787# 0.269531f
C731 a_n100_n70427# a_n100_n71463# 0.205388f
C732 a_n100_38353# a_n158_38450# 0.090922f
C733 a_n100_n41419# a_n158_n41322# 0.090922f
C734 a_n158_114078# a_n100_113981# 0.090922f
C735 a_n158_13586# a_100_13586# 0.219309f
C736 a_n100_n25879# w_n358_n132787# 0.269531f
C737 a_n100_116053# w_n358_n132787# 0.269531f
C738 a_n158_7370# w_n358_n132787# 0.240254f
C739 a_n100_n28987# a_100_n28890# 0.090922f
C740 a_100_n96230# a_100_n95194# 0.010536f
C741 a_100_114078# a_100_113042# 0.010536f
C742 a_n100_n89075# a_n100_n88039# 0.205388f
C743 a_n100_57001# a_n100_55965# 0.205388f
C744 a_100_90250# a_100_91286# 0.010536f
C745 a_100_n90014# a_100_n88978# 0.010536f
C746 a_n100_27993# a_100_28090# 0.090922f
C747 a_n158_n101410# a_n100_n101507# 0.090922f
C748 a_n100_49749# a_100_49846# 0.090922f
C749 a_100_126510# w_n358_n132787# 0.240254f
C750 a_100_n36142# a_100_n37178# 0.010536f
C751 a_n100_104657# a_n100_105693# 0.205388f
C752 a_n158_n111770# a_100_n111770# 0.219309f
C753 a_n100_17633# a_n158_17730# 0.090922f
C754 a_100_n96230# w_n358_n132787# 0.240254f
C755 a_n100_n4123# a_100_n4026# 0.090922f
C756 a_n100_n104615# a_n100_n105651# 0.205388f
C757 a_n158_n130418# a_100_n130418# 0.219309f
C758 a_n100_n130515# a_n100_n131551# 0.205388f
C759 a_n158_n10242# a_n158_n9206# 0.010536f
C760 a_100_n54790# w_n358_n132787# 0.240254f
C761 a_n100_n94255# w_n358_n132787# 0.269531f
C762 a_n158_35342# a_n158_34306# 0.010536f
C763 a_100_n44430# a_100_n45466# 0.010536f
C764 a_100_n29926# w_n358_n132787# 0.240254f
C765 a_100_71602# w_n358_n132787# 0.240254f
C766 a_n100_n5159# a_100_n5062# 0.090922f
C767 a_100_1154# w_n358_n132787# 0.240254f
C768 a_100_n108662# a_100_n107626# 0.010536f
C769 a_n158_n108662# a_n100_n108759# 0.090922f
C770 a_100_103718# w_n358_n132787# 0.240254f
C771 a_100_58134# w_n358_n132787# 0.240254f
C772 a_n100_41461# a_n158_41558# 0.090922f
C773 a_100_n80690# a_100_n79654# 0.010536f
C774 a_n100_2093# a_n100_1057# 0.205388f
C775 a_n100_44569# a_n100_45605# 0.205388f
C776 a_n100_104657# w_n358_n132787# 0.269531f
C777 w_n358_n132787# a_n158_n123166# 0.240254f
C778 a_n158_n99338# w_n358_n132787# 0.240254f
C779 a_n100_103621# w_n358_n132787# 0.269531f
C780 a_n158_n22674# w_n358_n132787# 0.240254f
C781 a_n158_73674# a_n158_74710# 0.010536f
C782 a_n158_n106590# w_n358_n132787# 0.240254f
C783 a_n158_n46502# a_n158_n47538# 0.010536f
C784 a_n100_n48671# a_n100_n49707# 0.205388f
C785 a_n100_n114975# a_100_n114878# 0.090922f
C786 a_n158_n68258# w_n358_n132787# 0.240254f
C787 a_100_62278# a_100_63314# 0.010536f
C788 a_n158_n79654# a_n158_n78618# 0.010536f
C789 a_100_78854# a_100_79890# 0.010536f
C790 a_n100_87045# a_n100_88081# 0.205388f
C791 a_n158_n33034# a_n158_n34070# 0.010536f
C792 a_100_n102446# w_n358_n132787# 0.240254f
C793 a_n100_48713# a_n158_48810# 0.090922f
C794 a_100_n22674# a_n158_n22674# 0.219309f
C795 a_n100_n130515# w_n358_n132787# 0.269531f
C796 a_n158_n92086# a_100_n92086# 0.219309f
C797 a_n100_110873# a_n100_109837# 0.205388f
C798 a_n100_20741# w_n358_n132787# 0.269531f
C799 a_n158_n918# a_n158_n1954# 0.010536f
C800 a_n158_n76546# w_n358_n132787# 0.240254f
C801 a_100_n100374# a_100_n99338# 0.010536f
C802 a_n158_n41322# a_100_n41322# 0.219309f
C803 a_100_n10242# a_100_n11278# 0.010536f
C804 a_n158_n28890# w_n358_n132787# 0.240254f
C805 a_n100_119161# w_n358_n132787# 0.269531f
C806 a_n158_12550# a_100_12550# 0.219309f
C807 a_n158_56062# a_100_56062# 0.219309f
C808 a_n158_n84834# a_n158_n83798# 0.010536f
C809 a_100_n50646# a_n100_n50743# 0.090922f
C810 a_100_59170# w_n358_n132787# 0.240254f
C811 a_n158_n51682# a_n158_n52718# 0.010536f
C812 a_n100_106729# a_n100_105693# 0.205388f
C813 a_n100_101549# a_n100_102585# 0.205388f
C814 a_n158_112006# a_n100_111909# 0.090922f
C815 a_n100_4165# a_n100_3129# 0.205388f
C816 a_n100_n105651# a_100_n105554# 0.090922f
C817 a_n100_n83895# a_n100_n82859# 0.205388f
C818 a_n100_76685# a_n158_76782# 0.090922f
C819 a_100_92322# w_n358_n132787# 0.240254f
C820 a_100_n97266# a_n100_n97363# 0.090922f
C821 a_n100_n101507# a_n100_n100471# 0.205388f
C822 a_n158_n76546# a_n158_n75510# 0.010536f
C823 a_n158_n120058# a_100_n120058# 0.219309f
C824 a_n100_n120155# a_n100_n121191# 0.205388f
C825 a_100_86106# a_n100_86009# 0.090922f
C826 a_100_55026# w_n358_n132787# 0.240254f
C827 a_n158_n77582# a_n158_n76546# 0.010536f
C828 a_n100_n53851# a_n158_n53754# 0.090922f
C829 a_100_102682# a_n158_102682# 0.219309f
C830 a_n158_22910# a_n158_21874# 0.010536f
C831 a_n100_106729# w_n358_n132787# 0.269531f
C832 a_n100_n117047# a_100_n116950# 0.090922f
C833 a_n100_n20699# a_n100_n21735# 0.205388f
C834 a_n100_25921# w_n358_n132787# 0.269531f
C835 a_100_86106# a_100_85070# 0.010536f
C836 a_n100_1057# a_n100_21# 0.205388f
C837 a_n158_n39250# a_n100_n39347# 0.090922f
C838 a_n100_108801# w_n358_n132787# 0.269531f
C839 a_n158_122366# w_n358_n132787# 0.240254f
C840 a_100_14622# a_100_13586# 0.010536f
C841 a_n100_n27951# a_n158_n27854# 0.090922f
C842 a_n100_n92183# a_n158_n92086# 0.090922f
C843 a_n158_9442# w_n358_n132787# 0.240254f
C844 a_100_30162# a_100_29126# 0.010536f
C845 a_n100_29029# a_n158_29126# 0.090922f
C846 a_100_n119022# w_n358_n132787# 0.240254f
C847 a_100_n76546# w_n358_n132787# 0.240254f
C848 a_100_50882# a_100_51918# 0.010536f
C849 a_n100_129521# a_n158_129618# 0.090922f
C850 a_100_78854# a_100_77818# 0.010536f
C851 a_100_103718# a_n100_103621# 0.090922f
C852 a_n100_6237# a_n100_5201# 0.205388f
C853 a_n100_n36239# a_n158_n36142# 0.090922f
C854 a_n100_104657# a_n100_103621# 0.205388f
C855 a_100_n9206# a_n100_n9303# 0.090922f
C856 a_n158_85070# a_n158_86106# 0.010536f
C857 a_n100_n56959# a_n100_n55923# 0.205388f
C858 a_n100_83937# w_n358_n132787# 0.269531f
C859 a_n100_n102543# w_n358_n132787# 0.269531f
C860 a_n100_n123263# a_100_n123166# 0.090922f
C861 a_n158_124438# a_100_124438# 0.219309f
C862 a_n158_72638# a_n158_71602# 0.010536f
C863 a_n158_n90014# a_n158_n88978# 0.010536f
C864 a_n158_n1954# a_n158_n2990# 0.010536f
C865 a_100_n126274# a_100_n127310# 0.010536f
C866 a_n100_n127407# a_n158_n127310# 0.090922f
C867 a_n100_n102543# a_n100_n103579# 0.205388f
C868 a_100_n79654# w_n358_n132787# 0.240254f
C869 a_n100_n110831# w_n358_n132787# 0.269531f
C870 a_n100_86009# a_n100_84973# 0.205388f
C871 a_n100_73577# w_n358_n132787# 0.269531f
C872 a_n100_n12411# a_n100_n13447# 0.205388f
C873 a_n158_n29926# w_n358_n132787# 0.240254f
C874 a_n158_42594# a_100_42594# 0.219309f
C875 w_n358_n132787# a_n100_n71463# 0.269531f
C876 a_n100_2093# w_n358_n132787# 0.269531f
C877 a_n100_84973# a_100_85070# 0.090922f
C878 a_n100_128485# w_n358_n132787# 0.269531f
C879 a_n158_24982# a_100_24982# 0.219309f
C880 a_n100_n81823# a_n100_n80787# 0.205388f
C881 a_n158_51918# a_n158_50882# 0.010536f
C882 a_100_32234# w_n358_n132787# 0.240254f
C883 a_n100_48713# a_100_48810# 0.090922f
C884 a_100_n39250# a_100_n40286# 0.010536f
C885 a_n100_n23807# w_n358_n132787# 0.269531f
C886 a_n100_n73535# a_n100_n74571# 0.205388f
C887 a_100_n61006# w_n358_n132787# 0.240254f
C888 a_n100_15561# a_100_15658# 0.090922f
C889 a_n158_50882# w_n358_n132787# 0.240254f
C890 a_100_59170# a_100_58134# 0.010536f
C891 a_n100_n7231# a_n158_n7134# 0.090922f
C892 a_100_113042# a_n100_112945# 0.090922f
C893 a_100_84034# a_100_85070# 0.010536f
C894 a_n100_n126371# a_n158_n126274# 0.090922f
C895 a_n100_32137# a_n100_31101# 0.205388f
C896 a_n158_n87942# a_n158_n88978# 0.010536f
C897 a_100_n34070# a_100_n33034# 0.010536f
C898 a_n158_n110734# a_100_n110734# 0.219309f
C899 a_n100_n110831# a_n100_n111867# 0.205388f
C900 a_100_n4026# w_n358_n132787# 0.240254f
C901 a_100_n85870# w_n358_n132787# 0.240254f
C902 a_100_122366# a_n100_122269# 0.090922f
C903 a_100_n14386# w_n358_n132787# 0.240254f
C904 a_n158_84034# w_n358_n132787# 0.240254f
C905 a_n158_n52718# w_n358_n132787# 0.240254f
C906 a_n100_22813# w_n358_n132787# 0.269531f
C907 a_n100_44569# a_100_44666# 0.090922f
C908 a_n100_38353# a_100_38450# 0.090922f
C909 a_n100_n41419# a_100_n41322# 0.090922f
C910 a_n100_89117# a_n100_88081# 0.205388f
C911 a_n158_125474# a_n100_125377# 0.090922f
C912 a_n158_79890# w_n358_n132787# 0.240254f
C913 a_n158_68494# a_n158_67458# 0.010536f
C914 a_n100_n28987# a_n100_n30023# 0.205388f
C915 a_100_77818# a_100_76782# 0.010536f
C916 a_100_7370# w_n358_n132787# 0.240254f
C917 a_100_n92086# a_100_n91050# 0.010536f
C918 w_n358_n132787# a_n158_n122130# 0.240254f
C919 a_n100_36281# w_n358_n132787# 0.269531f
C920 a_n158_5298# a_100_5298# 0.219309f
C921 a_n100_5201# a_n100_4165# 0.205388f
C922 a_100_113042# w_n358_n132787# 0.240254f
C923 a_n100_n42455# w_n358_n132787# 0.269531f
C924 a_100_n65150# a_n158_n65150# 0.219309f
C925 a_n100_n37275# a_100_n37178# 0.090922f
C926 a_100_65386# a_n100_65289# 0.090922f
C927 a_n158_94394# a_n158_95430# 0.010536f
C928 a_100_n16458# w_n358_n132787# 0.240254f
C929 a_n158_n85870# w_n358_n132787# 0.240254f
C930 a_n158_n113842# a_n158_n114878# 0.010536f
C931 a_100_n58934# w_n358_n132787# 0.240254f
C932 a_n158_n4026# a_100_n4026# 0.219309f
C933 a_n100_n4123# a_n100_n5159# 0.205388f
C934 a_n158_n10242# a_100_n10242# 0.219309f
C935 a_n100_n10339# a_n100_n11375# 0.205388f
C936 a_100_122366# a_100_123402# 0.010536f
C937 a_n100_74613# a_n158_74710# 0.090922f
C938 a_100_69530# a_n158_69530# 0.219309f
C939 a_n100_34209# a_n158_34306# 0.090922f
C940 a_n100_n45563# a_n158_n45466# 0.090922f
C941 a_n100_n129479# w_n358_n132787# 0.269531f
C942 a_100_94394# a_100_95430# 0.010536f
C943 a_n158_n29926# a_100_n29926# 0.219309f
C944 a_n100_21# w_n358_n132787# 0.269531f
C945 a_100_n88978# a_n158_n88978# 0.219309f
C946 a_n158_115114# a_n100_115017# 0.090922f
C947 a_100_107862# a_n158_107862# 0.219309f
C948 a_100_70566# a_n158_70566# 0.219309f
C949 a_n100_n93219# a_100_n93122# 0.090922f
C950 a_n100_41461# a_100_41558# 0.090922f
C951 a_n100_94297# w_n358_n132787# 0.269531f
C952 a_100_n39250# a_100_n38214# 0.010536f
C953 a_n158_n115914# a_n158_n114878# 0.010536f
C954 a_n158_n83798# a_n158_n82762# 0.010536f
C955 a_n100_n26915# w_n358_n132787# 0.269531f
C956 a_100_n47538# a_100_n46502# 0.010536f
C957 a_n158_120294# w_n358_n132787# 0.240254f
C958 a_n158_64350# a_n158_65386# 0.010536f
C959 a_n158_n76546# a_100_n76546# 0.219309f
C960 a_n158_n14386# a_n100_n14483# 0.090922f
C961 a_n100_62181# a_n100_61145# 0.205388f
C962 a_n158_7370# a_100_7370# 0.219309f
C963 a_n100_n102543# a_100_n102446# 0.090922f
C964 a_n158_n96230# a_n158_n97266# 0.010536f
C965 a_n100_n34167# a_n158_n34070# 0.090922f
C966 a_n158_n7134# w_n358_n132787# 0.240254f
C967 a_100_20838# a_100_19802# 0.010536f
C968 a_n100_19705# a_n158_19802# 0.090922f
C969 a_n100_n18627# w_n358_n132787# 0.269531f
C970 a_n158_43630# a_n158_42594# 0.010536f
C971 a_100_n82762# a_100_n81726# 0.010536f
C972 a_n158_n115914# a_n158_n116950# 0.010536f
C973 a_n100_n11375# a_n100_n12411# 0.205388f
C974 a_n158_12550# a_n158_11514# 0.010536f
C975 a_n158_n28890# a_n158_n29926# 0.010536f
C976 a_n100_n87003# w_n358_n132787# 0.269531f
C977 a_n158_102682# w_n358_n132787# 0.240254f
C978 a_n158_76782# a_n158_77818# 0.010536f
C979 a_n100_71505# a_n100_70469# 0.205388f
C980 a_100_n45466# w_n358_n132787# 0.240254f
C981 a_n100_78757# w_n358_n132787# 0.269531f
C982 a_100_96466# w_n358_n132787# 0.240254f
C983 a_100_n117986# w_n358_n132787# 0.240254f
C984 a_n158_n96230# w_n358_n132787# 0.240254f
C985 a_n100_n20699# w_n358_n132787# 0.269531f
C986 a_n100_80829# a_n100_79793# 0.205388f
C987 a_100_121330# w_n358_n132787# 0.240254f
C988 a_n100_n5159# a_n100_n6195# 0.205388f
C989 a_n158_n69294# a_n100_n69391# 0.090922f
C990 a_n100_n24843# a_n158_n24746# 0.090922f
C991 a_n100_n26915# a_n100_n25879# 0.205388f
C992 a_n158_n122130# a_n158_n123166# 0.010536f
C993 a_n158_n34070# w_n358_n132787# 0.240254f
C994 a_n158_63314# a_100_63314# 0.219309f
C995 a_n100_n53851# a_100_n53754# 0.090922f
C996 a_100_n11278# w_n358_n132787# 0.240254f
C997 a_100_n77582# a_n100_n77679# 0.090922f
C998 a_n100_n74571# a_100_n74474# 0.090922f
C999 a_n158_26018# w_n358_n132787# 0.240254f
C1000 a_n158_40522# a_n158_39486# 0.010536f
C1001 a_100_89214# a_100_88178# 0.010536f
C1002 a_n158_119258# a_100_119258# 0.219309f
C1003 a_n158_110970# a_100_110970# 0.219309f
C1004 a_100_n65150# w_n358_n132787# 0.240254f
C1005 a_n100_118125# w_n358_n132787# 0.269531f
C1006 a_100_n75510# a_n100_n75607# 0.090922f
C1007 a_n100_n27951# a_100_n27854# 0.090922f
C1008 a_100_n126274# a_100_n125238# 0.010536f
C1009 a_n100_8309# w_n358_n132787# 0.269531f
C1010 a_100_108898# a_100_107862# 0.010536f
C1011 a_n158_104754# a_100_104754# 0.219309f
C1012 a_100_49846# a_100_50882# 0.010536f
C1013 a_n100_29029# a_100_29126# 0.090922f
C1014 a_n158_6334# a_100_6334# 0.219309f
C1015 a_n158_39486# w_n358_n132787# 0.240254f
C1016 a_n100_n16555# a_n158_n16458# 0.090922f
C1017 a_n158_n67222# a_n100_n67319# 0.090922f
C1018 a_n100_n36239# a_100_n36142# 0.090922f
C1019 a_100_80926# w_n358_n132787# 0.240254f
C1020 a_100_n9206# a_n158_n9206# 0.219309f
C1021 a_n100_18669# a_n158_18766# 0.090922f
C1022 a_100_n1954# a_100_n2990# 0.010536f
C1023 a_n100_n3087# a_n158_n2990# 0.090922f
C1024 a_n158_n129382# a_100_n129382# 0.219309f
C1025 a_n100_n129479# a_n100_n130515# 0.205388f
C1026 a_n158_n21638# a_100_n21638# 0.219309f
C1027 a_n158_90250# a_n158_91286# 0.010536f
C1028 a_100_81962# a_100_82998# 0.010536f
C1029 w_n358_n132787# a_n100_n108759# 0.269531f
C1030 a_n100_n63175# w_n358_n132787# 0.269531f
C1031 a_100_n87942# a_n100_n88039# 0.090922f
C1032 a_100_n92086# a_100_n93122# 0.010536f
C1033 a_n100_n50743# a_n158_n50646# 0.090922f
C1034 a_n100_66325# w_n358_n132787# 0.269531f
C1035 a_100_n96230# a_n158_n96230# 0.219309f
C1036 a_n158_48810# a_100_48810# 0.219309f
C1037 a_n100_48713# a_n100_47677# 0.205388f
C1038 a_100_56062# w_n358_n132787# 0.240254f
C1039 a_n158_3226# a_n158_2190# 0.010536f
C1040 a_n100_n104615# a_100_n104518# 0.090922f
C1041 a_n158_n40286# a_100_n40286# 0.219309f
C1042 a_n100_n95291# a_n100_n96327# 0.205388f
C1043 w_n358_n132787# a_n158_n121094# 0.240254f
C1044 a_n100_67361# a_n100_68397# 0.205388f
C1045 a_n100_43533# w_n358_n132787# 0.269531f
C1046 a_n158_n66186# a_n158_n65150# 0.010536f
C1047 a_100_n25782# a_n158_n25782# 0.219309f
C1048 a_n100_n7231# a_100_n7134# 0.090922f
C1049 a_n100_12453# w_n358_n132787# 0.269531f
C1050 a_n158_32234# a_n158_31198# 0.010536f
C1051 a_n100_n113939# a_100_n113842# 0.090922f
C1052 a_n158_n83798# w_n358_n132787# 0.240254f
C1053 a_n158_84034# a_n100_83937# 0.090922f
C1054 a_n100_n132587# a_100_n132490# 0.090922f
C1055 a_100_n37178# w_n358_n132787# 0.240254f
C1056 a_n158_117186# a_n158_116150# 0.010536f
C1057 a_n100_n5159# w_n358_n132787# 0.269531f
C1058 a_n158_80926# a_n158_81962# 0.010536f
C1059 a_n100_n128443# w_n358_n132787# 0.269531f
C1060 a_n100_n99435# w_n358_n132787# 0.269531f
C1061 a_n100_n56959# a_n158_n56862# 0.090922f
C1062 a_100_n52718# w_n358_n132787# 0.240254f
C1063 a_n100_n21735# a_n158_n21638# 0.090922f
C1064 a_n100_38353# a_n100_37317# 0.205388f
C1065 a_n100_86009# w_n358_n132787# 0.269531f
C1066 a_100_86106# a_n158_86106# 0.219309f
C1067 a_n100_6237# w_n358_n132787# 0.269531f
C1068 a_100_n64114# a_n158_n64114# 0.219309f
C1069 a_n100_n65247# a_n100_n64211# 0.205388f
C1070 a_n158_28090# a_100_28090# 0.219309f
C1071 a_100_85070# w_n358_n132787# 0.240254f
C1072 a_n158_n18530# a_n158_n19566# 0.010536f
C1073 a_n158_n42358# w_n358_n132787# 0.240254f
C1074 a_n158_82998# w_n358_n132787# 0.240254f
C1075 a_n100_n37275# a_n100_n38311# 0.205388f
C1076 a_n158_n55826# a_n100_n55923# 0.090922f
C1077 a_100_n56862# a_100_n57898# 0.010536f
C1078 a_n158_n17494# w_n358_n132787# 0.240254f
C1079 a_100_107862# a_100_106826# 0.010536f
C1080 a_100_n114878# w_n358_n132787# 0.240254f
C1081 a_100_16694# w_n358_n132787# 0.240254f
C1082 a_100_68494# a_n100_68397# 0.090922f
C1083 a_n100_62181# a_100_62278# 0.090922f
C1084 a_n100_34209# a_100_34306# 0.090922f
C1085 a_n158_69530# w_n358_n132787# 0.240254f
C1086 a_n158_91286# a_100_91286# 0.219309f
C1087 a_100_n103482# a_100_n104518# 0.010536f
C1088 a_n100_81865# a_n158_81962# 0.090922f
C1089 a_100_n6098# a_100_n5062# 0.010536f
C1090 a_100_n8170# w_n358_n132787# 0.240254f
C1091 a_100_n104518# a_100_n105554# 0.010536f
C1092 a_n100_n116011# a_100_n115914# 0.090922f
C1093 a_n158_87142# w_n358_n132787# 0.240254f
C1094 a_n158_2190# a_n158_1154# 0.010536f
C1095 a_n100_82901# a_100_82998# 0.090922f
C1096 a_n158_97502# a_n158_98538# 0.010536f
C1097 a_100_100610# a_n158_100610# 0.219309f
C1098 a_n100_27993# w_n358_n132787# 0.269531f
C1099 a_100_n39250# a_n100_n39347# 0.090922f
C1100 a_n158_n26818# w_n358_n132787# 0.240254f
C1101 a_n100_91189# a_n100_92225# 0.205388f
C1102 a_n158_10478# w_n358_n132787# 0.240254f
C1103 a_n100_118125# a_n100_119161# 0.205388f
C1104 a_n100_87045# a_100_87142# 0.090922f
C1105 a_100_n116950# w_n358_n132787# 0.240254f
C1106 a_n100_100513# w_n358_n132787# 0.269531f
C1107 a_n100_30065# a_n158_30162# 0.090922f
C1108 a_100_115114# a_100_116150# 0.010536f
C1109 a_100_115114# a_100_114078# 0.010536f
C1110 a_n158_n10242# w_n358_n132787# 0.240254f
C1111 a_100_n63078# w_n358_n132787# 0.240254f
C1112 a_n158_n38214# w_n358_n132787# 0.240254f
C1113 a_n100_n98399# w_n358_n132787# 0.269531f
C1114 a_100_n85870# a_n158_n85870# 0.219309f
C1115 a_100_42594# w_n358_n132787# 0.240254f
C1116 a_100_n7134# w_n358_n132787# 0.240254f
C1117 a_n100_19705# a_100_19802# 0.090922f
C1118 a_n100_n122227# a_100_n122130# 0.090922f
C1119 a_n100_n109795# w_n358_n132787# 0.269531f
C1120 a_n158_20838# w_n358_n132787# 0.240254f
C1121 a_100_n918# a_100_n1954# 0.010536f
C1122 a_n158_n86906# w_n358_n132787# 0.240254f
C1123 a_n158_37414# a_n158_36378# 0.010536f
C1124 a_100_n117986# a_100_n119022# 0.010536f
C1125 a_n100_n119119# a_n158_n119022# 0.090922f
C1126 a_n158_96466# w_n358_n132787# 0.240254f
C1127 a_100_12550# a_100_11514# 0.010536f
C1128 a_n100_11417# a_n158_11514# 0.090922f
C1129 a_n158_n92086# a_n158_n93122# 0.010536f
C1130 a_n158_n66186# w_n358_n132787# 0.240254f
C1131 a_n100_124341# a_100_124438# 0.090922f
C1132 a_n100_4165# w_n358_n132787# 0.269531f
C1133 a_100_27054# a_100_26018# 0.010536f
C1134 a_n100_25921# a_n158_26018# 0.090922f
C1135 a_100_n50646# a_100_n51682# 0.010536f
C1136 a_n158_129618# w_n358_n132787# 0.240254f
C1137 a_n100_33173# w_n358_n132787# 0.269531f
C1138 a_n100_n99435# a_n158_n99338# 0.090922f
C1139 a_n100_n106687# a_n100_n107723# 0.205388f
C1140 a_n158_n92086# a_n158_n91050# 0.010536f
C1141 a_n100_n57995# a_n158_n57898# 0.090922f
C1142 a_n100_n76643# a_n100_n77679# 0.205388f
C1143 a_n100_16597# a_n158_16694# 0.090922f
C1144 a_n158_97502# a_n100_97405# 0.090922f
C1145 a_n158_99574# a_n158_100610# 0.010536f
C1146 a_100_65386# a_100_66422# 0.010536f
C1147 a_n158_33270# a_n158_32234# 0.010536f
C1148 a_100_n124202# a_100_n125238# 0.010536f
C1149 a_n100_n125335# a_n158_n125238# 0.090922f
C1150 a_n100_n90111# w_n358_n132787# 0.269531f
C1151 a_n100_48713# a_n100_49749# 0.205388f
C1152 a_n158_n97266# a_n100_n97363# 0.090922f
C1153 a_100_n12314# a_100_n13350# 0.010536f
C1154 a_n158_47774# w_n358_n132787# 0.240254f
C1155 a_n158_n109698# a_100_n109698# 0.219309f
C1156 a_n158_n1954# w_n358_n132787# 0.240254f
C1157 a_100_104754# w_n358_n132787# 0.240254f
C1158 a_n158_n20602# a_100_n20602# 0.219309f
C1159 a_100_68494# a_n158_68494# 0.219309f
C1160 a_n158_75746# a_n158_74710# 0.010536f
C1161 a_n100_24885# w_n358_n132787# 0.269531f
C1162 a_n158_1154# a_n158_118# 0.010536f
C1163 a_100_n49610# w_n358_n132787# 0.240254f
C1164 a_100_55026# a_100_56062# 0.010536f
C1165 a_100_n40286# a_100_n41322# 0.010536f
C1166 a_n100_92225# w_n358_n132787# 0.269531f
C1167 a_100_n71366# a_n158_n71366# 0.219309f
C1168 a_n100_n27951# a_n100_n28987# 0.205388f
C1169 w_n358_n132787# a_n158_n120058# 0.240254f
C1170 a_n158_29126# a_100_29126# 0.219309f
C1171 a_n100_n97363# w_n358_n132787# 0.269531f
C1172 a_100_39486# w_n358_n132787# 0.240254f
C1173 a_n100_n36239# a_n100_n37275# 0.205388f
C1174 a_100_n72402# a_100_n73438# 0.010536f
C1175 a_n158_n112806# a_n158_n113842# 0.010536f
C1176 a_100_n9206# a_100_n10242# 0.010536f
C1177 a_n158_n131454# a_n158_n132490# 0.010536f
C1178 a_100_18766# w_n358_n132787# 0.240254f
C1179 a_100_130654# a_n158_130654# 0.219309f
C1180 a_n100_64253# a_n100_63217# 0.205388f
C1181 a_n100_53893# a_n100_52857# 0.205388f
C1182 a_n100_n3087# a_n100_n4123# 0.205388f
C1183 a_100_n75510# w_n358_n132787# 0.240254f
C1184 a_n100_n44527# a_n158_n44430# 0.090922f
C1185 a_n158_n30962# w_n358_n132787# 0.240254f
C1186 a_n100_n127407# w_n358_n132787# 0.269531f
C1187 a_100_11514# a_100_10478# 0.010536f
C1188 a_n158_n62042# a_n100_n62139# 0.090922f
C1189 a_n100_53893# a_100_53990# 0.090922f
C1190 a_n158_42594# a_n158_41558# 0.010536f
C1191 a_n100_n30023# a_n100_n31059# 0.205388f
C1192 a_n158_24982# a_n158_23946# 0.010536f
C1193 a_n100_n19663# a_n158_n19566# 0.090922f
C1194 a_100_128582# w_n358_n132787# 0.240254f
C1195 a_n158_31198# w_n358_n132787# 0.240254f
C1196 w_n358_n132787# a_n100_n126371# 0.269531f
C1197 a_n100_n92183# a_n100_n93219# 0.205388f
C1198 a_n158_n21638# w_n358_n132787# 0.240254f
C1199 a_n158_15658# a_n158_14622# 0.010536f
C1200 a_n158_43630# w_n358_n132787# 0.240254f
C1201 a_n158_n57898# a_100_n57898# 0.219309f
C1202 a_n158_123402# a_n158_124438# 0.010536f
C1203 a_n100_95333# a_n100_96369# 0.205388f
C1204 a_n158_n24746# a_100_n24746# 0.219309f
C1205 a_100_47774# a_100_46738# 0.010536f
C1206 a_100_n75510# a_n158_n75510# 0.219309f
C1207 a_n100_69433# a_n100_70469# 0.205388f
C1208 a_100_n62042# a_n100_n62139# 0.090922f
C1209 a_n100_71505# w_n358_n132787# 0.269531f
C1210 a_n100_n38311# w_n358_n132787# 0.269531f
C1211 a_100_n113842# w_n358_n132787# 0.240254f
C1212 a_n100_n84931# a_100_n84834# 0.090922f
C1213 a_100_101646# a_100_102682# 0.010536f
C1214 a_n100_n15519# w_n358_n132787# 0.269531f
C1215 a_100_n132490# w_n358_n132787# 0.244798f
C1216 a_100_n82762# a_n100_n82859# 0.090922f
C1217 a_100_21874# a_100_20838# 0.010536f
C1218 a_n100_20741# a_n158_20838# 0.090922f
C1219 a_n100_n54887# a_n158_n54790# 0.090922f
C1220 a_100_112006# w_n358_n132787# 0.240254f
C1221 a_n158_44666# a_n158_43630# 0.010536f
C1222 a_n100_n1015# a_100_n918# 0.090922f
C1223 a_100_22910# w_n358_n132787# 0.240254f
C1224 a_n158_38450# a_n158_37414# 0.010536f
C1225 a_100_119258# a_100_118222# 0.010536f
C1226 a_n158_n43394# a_100_n43394# 0.219309f
C1227 a_100_n26818# w_n358_n132787# 0.240254f
C1228 a_n100_n72499# a_n158_n72402# 0.090922f
C1229 a_n158_13586# a_n158_12550# 0.010536f
C1230 a_n158_113042# a_n100_112945# 0.090922f
C1231 a_n158_n74474# w_n358_n132787# 0.240254f
C1232 a_100_103718# a_100_104754# 0.010536f
C1233 a_n100_104657# a_100_104754# 0.090922f
C1234 a_n100_n49707# a_n158_n49610# 0.090922f
C1235 a_100_n17494# a_n100_n17591# 0.090922f
C1236 a_n158_36378# w_n358_n132787# 0.240254f
C1237 a_n100_124341# a_n100_125377# 0.205388f
C1238 a_100_77818# a_n100_77721# 0.090922f
C1239 a_n158_99574# a_n158_98538# 0.010536f
C1240 a_100_94394# a_100_93358# 0.010536f
C1241 a_100_n115914# w_n358_n132787# 0.240254f
C1242 a_n100_n105651# w_n358_n132787# 0.269531f
C1243 a_100_n18530# w_n358_n132787# 0.240254f
C1244 a_n100_17633# a_100_17730# 0.090922f
C1245 a_n158_114078# a_n158_115114# 0.010536f
C1246 w_n358_n132787# a_n158_n69294# 0.240254f
C1247 a_100_78854# a_n158_78854# 0.219309f
C1248 a_n100_15561# w_n358_n132787# 0.269531f
C1249 a_n158_34306# a_100_34306# 0.219309f
C1250 a_n158_n121094# a_n158_n122130# 0.010536f
C1251 a_n100_n45563# a_n100_n46599# 0.205388f
C1252 a_n158_131690# a_100_131690# 0.219309f
C1253 w_n358_n132787# a_n158_130654# 0.240254f
C1254 a_n100_131593# a_n100_130557# 0.205388f
C1255 a_n158_n75510# a_n158_n74474# 0.010536f
C1256 a_100_125474# w_n358_n132787# 0.240254f
C1257 a_n158_n103482# a_100_n103482# 0.219309f
C1258 a_n158_10478# a_n158_9442# 0.010536f
C1259 a_n100_n88039# w_n358_n132787# 0.269531f
C1260 a_n100_n68355# a_n100_n69391# 0.205388f
C1261 a_100_118# w_n358_n132787# 0.240254f
C1262 a_n158_n19566# a_n158_n20602# 0.010536f
C1263 a_n158_n91050# a_100_n91050# 0.219309f
C1264 a_n158_113042# w_n358_n132787# 0.240254f
C1265 a_n158_n52718# a_100_n52718# 0.219309f
C1266 a_n100_n47635# w_n358_n132787# 0.269531f
C1267 a_n100_n70427# a_n158_n70330# 0.090922f
C1268 a_100_110970# w_n358_n132787# 0.240254f
C1269 a_n158_51918# a_100_51918# 0.219309f
C1270 a_n158_n67222# w_n358_n132787# 0.240254f
C1271 a_n158_49846# w_n358_n132787# 0.240254f
C1272 a_100_51918# w_n358_n132787# 0.240254f
C1273 a_100_n78618# a_n100_n78715# 0.090922f
C1274 a_100_n73438# w_n358_n132787# 0.240254f
C1275 a_n100_53893# a_n100_54929# 0.205388f
C1276 a_n158_n67222# a_100_n67222# 0.219309f
C1277 a_n100_n67319# a_n100_n68355# 0.205388f
C1278 a_n100_n60067# a_n100_n61103# 0.205388f
C1279 a_n100_30065# a_100_30162# 0.090922f
C1280 a_n158_84034# a_n158_82998# 0.010536f
C1281 a_n100_n72499# a_100_n72402# 0.090922f
C1282 a_n100_n85967# a_n100_n84931# 0.205388f
C1283 a_100_71602# a_n100_71505# 0.090922f
C1284 a_n158_n56862# a_n158_n55826# 0.010536f
C1285 a_n158_n18530# w_n358_n132787# 0.240254f
C1286 a_100_115114# w_n358_n132787# 0.240254f
C1287 a_n100_n110831# a_n100_n109795# 0.205388f
C1288 a_n158_n21638# a_n158_n22674# 0.010536f
C1289 a_n158_n128346# a_100_n128346# 0.219309f
C1290 a_n100_n128443# a_n100_n129479# 0.205388f
C1291 a_100_n98302# a_n158_n98302# 0.219309f
C1292 a_n158_56062# a_n100_55965# 0.090922f
C1293 a_n100_n2051# a_100_n1954# 0.090922f
C1294 a_n158_108898# a_n158_107862# 0.010536f
C1295 a_n158_n11278# a_n158_n12314# 0.010536f
C1296 a_n100_69433# a_100_69530# 0.090922f
C1297 a_n100_n42455# a_n158_n42358# 0.090922f
C1298 a_100_37414# a_100_36378# 0.010536f
C1299 a_100_n78618# w_n358_n132787# 0.240254f
C1300 a_100_92322# a_n100_92225# 0.090922f
C1301 a_n158_11514# a_100_11514# 0.219309f
C1302 a_n100_11417# a_n100_10381# 0.205388f
C1303 a_100_114078# a_n100_113981# 0.090922f
C1304 a_100_n64114# w_n358_n132787# 0.240254f
C1305 a_n100_51821# a_n100_50785# 0.205388f
C1306 a_n158_4262# w_n358_n132787# 0.240254f
C1307 a_n100_n92183# a_100_n92086# 0.090922f
C1308 a_n100_25921# a_n100_24885# 0.205388f
C1309 a_n158_86106# w_n358_n132787# 0.240254f
C1310 a_n158_33270# w_n358_n132787# 0.240254f
C1311 a_n100_n91147# a_100_n91050# 0.090922f
C1312 a_100_90250# w_n358_n132787# 0.240254f
C1313 a_100_n6098# a_n100_n6195# 0.090922f
C1314 a_n100_n57995# a_n100_n59031# 0.205388f
C1315 a_n158_60206# a_100_60206# 0.219309f
C1316 a_100_125474# a_100_126510# 0.010536f
C1317 a_n158_90250# a_n100_90153# 0.090922f
C1318 a_n158_71602# w_n358_n132787# 0.240254f
C1319 a_n100_n112903# a_100_n112806# 0.090922f
C1320 a_100_63314# w_n358_n132787# 0.240254f
C1321 a_n158_n45466# a_n158_n46502# 0.010536f
C1322 a_n100_n96327# w_n358_n132787# 0.269531f
C1323 a_n100_n36239# w_n358_n132787# 0.269531f
C1324 a_n100_n131551# a_100_n131454# 0.090922f
C1325 a_n100_107765# w_n358_n132787# 0.269531f
C1326 a_n100_n3087# w_n358_n132787# 0.269531f
C1327 a_100_n12314# w_n358_n132787# 0.240254f
C1328 a_n100_101549# a_n158_101646# 0.090922f
C1329 a_n100_n50743# w_n358_n132787# 0.269531f
C1330 a_100_77818# a_n158_77818# 0.219309f
C1331 a_n158_n104518# a_100_n104518# 0.219309f
C1332 a_100_1154# a_100_118# 0.010536f
C1333 a_n158_24982# w_n358_n132787# 0.240254f
C1334 a_n158_127546# w_n358_n132787# 0.240254f
C1335 a_n100_65289# w_n358_n132787# 0.269531f
C1336 w_n358_n132787# a_n100_n125335# 0.269531f
C1337 a_100_n75510# a_100_n76546# 0.010536f
C1338 a_100_n101410# a_n158_n101410# 0.219309f
C1339 a_100_n106590# a_100_n107626# 0.010536f
C1340 a_n100_n107723# a_n158_n107626# 0.090922f
C1341 a_n158_n68258# a_n158_n69294# 0.010536f
C1342 a_n158_109934# a_n158_108898# 0.010536f
C1343 a_n158_38450# w_n358_n132787# 0.240254f
C1344 a_n158_n36142# a_n158_n37178# 0.010536f
C1345 a_n158_n63078# a_n158_n62042# 0.010536f
C1346 a_n158_n86906# a_n158_n85870# 0.010536f
C1347 a_n158_n61006# a_n100_n61103# 0.090922f
C1348 a_n100_n26915# a_n158_n26818# 0.090922f
C1349 a_n158_76782# w_n358_n132787# 0.240254f
C1350 a_n100_18669# a_n100_17633# 0.205388f
C1351 a_n158_17730# w_n358_n132787# 0.240254f
C1352 a_n158_n2990# a_100_n2990# 0.219309f
C1353 a_100_n112806# w_n358_n132787# 0.240254f
C1354 a_n100_35245# a_n158_35342# 0.090922f
C1355 a_n158_n44430# a_100_n44430# 0.219309f
C1356 a_100_n131454# w_n358_n132787# 0.240254f
C1357 a_n158_119258# w_n358_n132787# 0.240254f
C1358 a_n158_n29926# a_n158_n30962# 0.010536f
C1359 a_n158_n67222# a_n158_n68258# 0.010536f
C1360 a_100_n30962# a_n100_n31059# 0.090922f
C1361 a_100_2190# w_n358_n132787# 0.240254f
C1362 a_100_24982# a_100_23946# 0.010536f
C1363 a_100_108898# a_n158_108898# 0.219309f
C1364 a_100_61242# a_100_60206# 0.010536f
C1365 a_100_101646# w_n358_n132787# 0.240254f
C1366 a_n158_66422# w_n358_n132787# 0.240254f
C1367 a_100_3226# a_100_2190# 0.010536f
C1368 a_100_70566# a_n100_70469# 0.090922f
C1369 a_100_n70330# a_n158_n70330# 0.219309f
C1370 a_100_31198# w_n358_n132787# 0.240254f
C1371 a_n158_n73438# a_n158_n72402# 0.010536f
C1372 a_n100_n72499# w_n358_n132787# 0.269531f
C1373 a_n100_59073# a_n100_60109# 0.205388f
C1374 a_n100_n76643# a_n100_n75607# 0.205388f
C1375 a_n158_n93122# a_100_n93122# 0.219309f
C1376 a_100_n96230# a_n100_n96327# 0.090922f
C1377 a_n158_n7134# a_100_n7134# 0.219309f
C1378 a_100_71602# a_n158_71602# 0.219309f
C1379 a_100_65386# a_n158_65386# 0.219309f
C1380 a_100_12550# w_n358_n132787# 0.240254f
C1381 a_100_128582# a_n100_128485# 0.090922f
C1382 a_100_n9206# w_n358_n132787# 0.240254f
C1383 a_n158_95430# w_n358_n132787# 0.240254f
C1384 a_n158_n15422# w_n358_n132787# 0.240254f
C1385 a_n100_n121191# a_100_n121094# 0.090922f
C1386 a_100_n6098# w_n358_n132787# 0.240254f
C1387 a_100_88178# a_n100_88081# 0.090922f
C1388 a_n158_61242# a_n100_61145# 0.090922f
C1389 a_n100_n56959# a_100_n56862# 0.090922f
C1390 a_n158_n84834# a_n100_n84931# 0.090922f
C1391 a_n158_n23710# a_100_n23710# 0.219309f
C1392 w_n358_n132787# a_n158_131690# 0.244798f
C1393 a_n158_n53754# w_n358_n132787# 0.240254f
C1394 a_n158_n918# a_100_n918# 0.219309f
C1395 a_n100_n1015# a_n100_n2051# 0.205388f
C1396 a_100_n116950# a_100_n117986# 0.010536f
C1397 a_n100_n118083# a_n158_n117986# 0.090922f
C1398 a_n158_n27854# w_n358_n132787# 0.240254f
C1399 a_n100_n87003# a_n158_n86906# 0.090922f
C1400 a_n158_n91050# a_n158_n90014# 0.010536f
C1401 a_n158_6334# w_n358_n132787# 0.240254f
C1402 w_n358_n132787# a_n158_n70330# 0.240254f
C1403 a_100_74710# a_n158_74710# 0.219309f
C1404 a_n158_96466# a_100_96466# 0.219309f
C1405 a_100_n77582# w_n358_n132787# 0.240254f
C1406 a_n100_n19663# w_n358_n132787# 0.269531f
C1407 a_n100_17633# a_n100_16597# 0.205388f
C1408 a_100_n123166# a_100_n124202# 0.010536f
C1409 a_n100_n124299# a_n158_n124202# 0.090922f
C1410 a_n100_n78715# a_n100_n79751# 0.205388f
C1411 a_n100_n13447# a_n158_n13350# 0.090922f
C1412 a_100_n99338# w_n358_n132787# 0.240254f
C1413 a_n158_94394# a_n158_93358# 0.010536f
C1414 a_n100_117089# w_n358_n132787# 0.269531f
C1415 a_100_52954# a_n158_52954# 0.219309f
C1416 a_n100_22813# a_100_22910# 0.090922f
C1417 a_100_64350# a_n158_64350# 0.219309f
C1418 a_n100_n52815# a_n100_n53851# 0.205388f
C1419 a_100_n101410# a_100_n100374# 0.010536f
C1420 a_n158_28090# w_n358_n132787# 0.240254f
C1421 a_n158_n94158# a_n158_n95194# 0.010536f
C1422 a_100_2190# a_100_1154# 0.010536f
C1423 a_n158_41558# a_n158_40522# 0.010536f
C1424 a_n100_n43491# a_n158_n43394# 0.090922f
C1425 a_100_49846# w_n358_n132787# 0.240254f
C1426 a_n100_113981# a_n100_112945# 0.205388f
C1427 a_n158_n77582# a_100_n77582# 0.219309f
C1428 a_100_81962# a_n100_81865# 0.090922f
C1429 a_100_10478# w_n358_n132787# 0.240254f
C1430 a_100_113042# a_100_112006# 0.010536f
C1431 a_n100_n79751# w_n358_n132787# 0.269531f
C1432 a_n100_30065# a_n100_29029# 0.205388f
C1433 a_n158_n39250# w_n358_n132787# 0.240254f
C1434 a_n158_81962# w_n358_n132787# 0.240254f
C1435 a_n158_7370# a_n158_6334# 0.010536f
C1436 a_n100_n89075# a_n158_n88978# 0.090922f
C1437 a_100_70566# a_100_69530# 0.010536f
C1438 a_n158_41558# w_n358_n132787# 0.240254f
C1439 a_100_48810# a_100_47774# 0.010536f
C1440 a_n158_n111770# a_n158_n112806# 0.010536f
C1441 a_n100_19705# a_n100_18669# 0.205388f
C1442 a_n158_n130418# a_n158_n131454# 0.010536f
C1443 a_100_n81726# a_100_n80690# 0.010536f
C1444 a_n158_49846# a_n158_50882# 0.010536f
C1445 a_100_n63078# a_n100_n63175# 0.090922f
C1446 a_n158_n54790# w_n358_n132787# 0.240254f
C1447 a_n158_19802# w_n358_n132787# 0.240254f
C1448 a_n100_107765# a_n100_106729# 0.205388f
C1449 a_n100_n119119# a_n100_n120155# 0.205388f
C1450 a_n100_69433# w_n358_n132787# 0.269531f
C1451 a_n100_n101507# w_n358_n132787# 0.269531f
C1452 a_n100_36281# a_n158_36378# 0.090922f
C1453 a_n100_107765# a_n100_108801# 0.205388f
C1454 a_n100_n109795# a_n100_n108759# 0.205388f
C1455 a_100_n78618# a_100_n79654# 0.010536f
C1456 a_n100_n32095# a_n158_n31998# 0.090922f
C1457 a_n158_115114# a_n158_116150# 0.010536f
C1458 a_n100_117089# a_n100_116053# 0.205388f
C1459 a_n100_119161# a_n158_119258# 0.090922f
C1460 a_100_4262# w_n358_n132787# 0.240254f
C1461 a_n100_113981# w_n358_n132787# 0.269531f
C1462 w_n358_n132787# a_n100_n124299# 0.269531f
C1463 a_100_33270# w_n358_n132787# 0.240254f
C1464 a_n100_62181# a_n158_62278# 0.090922f
C1465 a_100_109934# w_n358_n132787# 0.240254f
C1466 a_100_4262# a_100_3226# 0.010536f
C1467 a_n100_3129# a_n158_3226# 0.090922f
C1468 a_n100_54929# a_n158_55026# 0.090922f
C1469 a_n158_n20602# w_n358_n132787# 0.240254f
C1470 a_n158_110970# a_n158_109934# 0.010536f
C1471 a_100_52954# w_n358_n132787# 0.240254f
C1472 a_n158_125474# w_n358_n132787# 0.240254f
C1473 a_n158_n59970# a_n158_n58934# 0.010536f
C1474 a_n100_n26915# a_100_n26818# 0.090922f
C1475 a_n100_n99435# a_n100_n98399# 0.205388f
C1476 a_n158_113042# a_100_113042# 0.219309f
C1477 a_100_95430# w_n358_n132787# 0.240254f
C1478 a_n100_32137# a_n158_32234# 0.090922f
C1479 a_n100_n13447# a_100_n13350# 0.090922f
C1480 a_n158_97502# w_n358_n132787# 0.240254f
C1481 a_100_n111770# w_n358_n132787# 0.240254f
C1482 a_n100_n33131# a_100_n33034# 0.090922f
C1483 a_100_n130418# w_n358_n132787# 0.240254f
C1484 a_100_122366# w_n358_n132787# 0.240254f
C1485 a_n158_n93122# a_n100_n93219# 0.090922f
C1486 a_n158_n5062# a_n158_n6098# 0.010536f
C1487 a_n158_45702# a_100_45702# 0.219309f
C1488 a_n158_n103482# a_n158_n104518# 0.010536f
C1489 a_n158_63314# a_n100_63217# 0.090922f
C1490 a_n100_21# a_100_118# 0.090922f
C1491 a_n158_72638# a_n158_73674# 0.010536f
C1492 a_100_60206# w_n358_n132787# 0.240254f
C1493 a_n158_39486# a_100_39486# 0.219309f
C1494 a_n100_39389# a_n100_38353# 0.205388f
C1495 a_100_66422# a_100_67458# 0.010536f
C1496 a_n158_n99338# a_100_n99338# 0.219309f
C1497 a_n100_60109# a_n100_61145# 0.205388f
C1498 a_n158_n24746# w_n358_n132787# 0.240254f
C1499 a_n158_n27854# a_n158_n28890# 0.010536f
C1500 a_n158_n107626# a_100_n107626# 0.219309f
C1501 a_100_8406# w_n358_n132787# 0.240254f
C1502 a_n100_n89075# a_100_n88978# 0.090922f
C1503 a_n100_n18627# a_100_n18530# 0.090922f
C1504 a_100_38450# w_n358_n132787# 0.240254f
C1505 a_n158_n73438# w_n358_n132787# 0.240254f
C1506 a_n100_81865# a_n100_82901# 0.205388f
C1507 a_n158_n54790# a_100_n54790# 0.219309f
C1508 a_n158_n16458# w_n358_n132787# 0.240254f
C1509 a_n100_n111867# a_100_n111770# 0.090922f
C1510 a_n100_46641# w_n358_n132787# 0.269531f
C1511 a_n158_n103482# a_n158_n102446# 0.010536f
C1512 a_n100_n8267# a_n158_n8170# 0.090922f
C1513 a_n100_n57995# w_n358_n132787# 0.269531f
C1514 a_n100_35245# a_n100_34209# 0.205388f
C1515 a_n158_n120058# a_n158_n121094# 0.010536f
C1516 a_n100_n44527# a_n100_n45563# 0.205388f
C1517 a_100_n7134# a_100_n8170# 0.010536f
C1518 a_n158_67458# a_100_67458# 0.219309f
C1519 a_n100_55965# w_n358_n132787# 0.269531f
C1520 a_n158_n80690# a_n158_n81726# 0.010536f
C1521 a_100_n66186# a_n100_n66283# 0.090922f
C1522 a_n100_23849# a_n158_23946# 0.090922f
C1523 a_n100_n87003# a_n100_n88039# 0.205388f
C1524 a_100_n104518# w_n358_n132787# 0.240254f
C1525 a_n100_n68355# w_n358_n132787# 0.269531f
C1526 a_n158_30162# w_n358_n132787# 0.240254f
C1527 a_n158_n47538# w_n358_n132787# 0.240254f
C1528 a_n100_127449# a_n100_126413# 0.205388f
C1529 a_n158_92322# w_n358_n132787# 0.240254f
C1530 a_n100_2093# a_100_2190# 0.090922f
C1531 a_n158_n57898# a_n158_n58934# 0.010536f
C1532 a_100_n81726# w_n358_n132787# 0.240254f
C1533 a_100_15658# a_100_14622# 0.010536f
C1534 a_n158_124438# w_n358_n132787# 0.240254f
C1535 a_n100_n72499# a_n100_n71463# 0.205388f
C1536 a_n158_11514# w_n358_n132787# 0.240254f
C1537 a_n100_123305# a_n100_124341# 0.205388f
C1538 a_n158_n48574# a_n158_n47538# 0.010536f
C1539 a_n100_n18627# a_n158_n18530# 0.090922f
C1540 a_100_32234# a_100_31198# 0.010536f
C1541 a_n158_n33034# a_100_n33034# 0.219309f
C1542 a_100_n34070# a_100_n35106# 0.010536f
C1543 a_100_117186# a_100_116150# 0.010536f
C1544 a_100_n110734# w_n358_n132787# 0.240254f
C1545 a_100_n15422# w_n358_n132787# 0.240254f
C1546 a_n158_n72402# a_n158_n71366# 0.010536f
C1547 a_n158_n127310# a_100_n127310# 0.219309f
C1548 a_n100_n127407# a_n100_n128443# 0.205388f
C1549 a_n158_n95194# a_n100_n95291# 0.090922f
C1550 a_n100_21777# w_n358_n132787# 0.269531f
C1551 a_100_n53754# w_n358_n132787# 0.240254f
C1552 a_100_44666# a_100_43630# 0.010536f
C1553 a_n100_43533# a_n158_43630# 0.090922f
C1554 a_n100_37317# a_n158_37414# 0.090922f
C1555 a_100_n42358# a_100_n41322# 0.010536f
C1556 a_100_n77582# a_100_n76546# 0.010536f
C1557 a_n100_n76643# w_n358_n132787# 0.269531f
C1558 a_100_n27854# w_n358_n132787# 0.240254f
C1559 a_n100_64253# a_n158_64350# 0.090922f
C1560 a_n158_n51682# a_100_n51682# 0.219309f
C1561 a_100_28090# a_100_27054# 0.010536f
C1562 a_100_66422# w_n358_n132787# 0.240254f
C1563 a_n158_n44430# w_n358_n132787# 0.240254f
C1564 a_100_97502# a_n100_97405# 0.090922f
C1565 a_n158_117186# w_n358_n132787# 0.240254f
C1566 a_n100_127449# w_n358_n132787# 0.269531f
C1567 a_n158_103718# a_n158_104754# 0.010536f
C1568 a_100_100610# w_n358_n132787# 0.240254f
C1569 a_100_102682# a_n100_102585# 0.090922f
C1570 a_n100_14525# w_n358_n132787# 0.269531f
C1571 a_100_n57898# w_n358_n132787# 0.240254f
C1572 a_n100_110873# a_n158_110970# 0.090922f
C1573 a_100_118222# w_n358_n132787# 0.240254f
C1574 a_n100_n130515# a_100_n130418# 0.090922f
C1575 a_n158_68494# a_n100_68397# 0.090922f
C1576 a_n158_n31998# a_n158_n33034# 0.010536f
C1577 a_n158_n52718# a_n158_n53754# 0.010536f
C1578 a_n100_57001# a_100_57098# 0.090922f
C1579 a_n158_67458# w_n358_n132787# 0.240254f
C1580 a_100_n19566# a_100_n20602# 0.010536f
C1581 a_n100_26957# w_n358_n132787# 0.269531f
C1582 a_n100_91189# a_n158_91286# 0.090922f
C1583 a_n100_53893# a_n158_53990# 0.090922f
C1584 a_n158_73674# a_100_73674# 0.219309f
C1585 a_n100_111909# a_n100_112945# 0.205388f
C1586 a_n100_n98399# a_n100_n97363# 0.205388f
C1587 a_n158_n96230# a_n100_n96327# 0.090922f
C1588 w_n358_n132787# a_n100_n123263# 0.269531f
C1589 a_n100_129521# a_100_129618# 0.090922f
C1590 a_100_n87942# a_100_n86906# 0.010536f
C1591 a_100_n65150# a_100_n64114# 0.010536f
C1592 a_n100_9345# w_n358_n132787# 0.269531f
C1593 a_100_n79654# a_n100_n79751# 0.090922f
C1594 a_n100_n51779# a_n158_n51682# 0.090922f
C1595 a_n158_n46502# a_100_n46502# 0.219309f
C1596 a_100_59170# a_100_60206# 0.010536f
C1597 a_100_41558# w_n358_n132787# 0.240254f
C1598 a_n158_119258# a_n158_120294# 0.010536f
C1599 a_n158_n79654# a_n158_n80690# 0.010536f
C1600 a_n158_126510# a_n100_126413# 0.090922f
C1601 a_100_70566# w_n358_n132787# 0.240254f
C1602 a_100_n113842# a_100_n114878# 0.010536f
C1603 a_n100_n114975# a_n158_n114878# 0.090922f
C1604 a_n100_47677# a_100_47774# 0.090922f
C1605 a_n158_52954# a_n100_52857# 0.090922f
C1606 a_n100_n102543# a_n100_n101507# 0.205388f
C1607 a_100_n53754# a_100_n54790# 0.010536f
C1608 a_n100_62181# w_n358_n132787# 0.269531f
C1609 a_n100_n21735# a_n100_n22771# 0.205388f
C1610 a_100_19802# w_n358_n132787# 0.240254f
C1611 a_100_n129382# w_n358_n132787# 0.240254f
C1612 a_n158_n82762# a_n158_n81726# 0.010536f
C1613 a_n158_n68258# a_n100_n68355# 0.090922f
C1614 a_100_n11278# a_100_n12314# 0.010536f
C1615 a_n100_n12411# a_n158_n12314# 0.090922f
C1616 a_n158_99574# w_n358_n132787# 0.240254f
C1617 a_n100_111909# w_n358_n132787# 0.269531f
C1618 a_n158_26018# a_n158_24982# 0.010536f
C1619 a_n100_88081# a_n158_88178# 0.090922f
C1620 a_100_n47538# w_n358_n132787# 0.240254f
C1621 a_n100_n83895# a_100_n83798# 0.090922f
C1622 a_100_122366# a_n158_122366# 0.219309f
C1623 a_n100_99477# w_n358_n132787# 0.269531f
C1624 a_100_n115914# a_100_n114878# 0.010536f
C1625 a_100_74710# a_n100_74613# 0.090922f
C1626 a_n100_32137# w_n358_n132787# 0.269531f
C1627 a_n158_n64114# a_n158_n63078# 0.010536f
C1628 a_n100_n38311# a_n158_n38214# 0.090922f
C1629 a_n100_n84931# w_n358_n132787# 0.269531f
C1630 a_n158_45702# w_n358_n132787# 0.240254f
C1631 a_n158_n26818# a_100_n26818# 0.219309f
C1632 a_100_79890# w_n358_n132787# 0.240254f
C1633 a_n158_16694# a_n158_15658# 0.010536f
C1634 a_100_n25782# a_100_n24746# 0.010536f
C1635 a_n100_13489# w_n358_n132787# 0.269531f
C1636 a_100_64350# a_n100_64253# 0.090922f
C1637 a_n100_n46599# a_n158_n46502# 0.090922f
C1638 a_100_33270# a_100_32234# 0.010536f
C1639 a_n158_n110734# a_n158_n111770# 0.010536f
C1640 a_100_97502# a_100_98538# 0.010536f
C1641 a_n158_126510# w_n358_n132787# 0.240254f
C1642 a_100_n2990# w_n358_n132787# 0.240254f
C1643 a_n100_n120155# a_100_n120058# 0.090922f
C1644 a_n100_21777# a_n100_20741# 0.205388f
C1645 a_n100_n13447# w_n358_n132787# 0.269531f
C1646 a_n100_87045# w_n358_n132787# 0.269531f
C1647 a_n158_91286# w_n358_n132787# 0.240254f
C1648 a_100_n51682# w_n358_n132787# 0.240254f
C1649 a_n158_45702# a_n158_44666# 0.010536f
C1650 a_n100_23849# w_n358_n132787# 0.269531f
C1651 a_n100_n76643# a_n158_n76546# 0.090922f
C1652 a_n100_98441# a_n158_98538# 0.090922f
C1653 a_n158_92322# a_100_92322# 0.219309f
C1654 a_100_n115914# a_100_n116950# 0.010536f
C1655 a_n100_n117047# a_n158_n116950# 0.090922f
C1656 a_n100_n81823# w_n358_n132787# 0.269531f
C1657 a_n158_39486# a_n158_38450# 0.010536f
C1658 a_n100_52857# w_n358_n132787# 0.269531f
C1659 a_100_n68258# w_n358_n132787# 0.240254f
C1660 a_n100_7273# w_n358_n132787# 0.269531f
C1661 a_n100_121233# a_n158_121330# 0.090922f
C1662 a_n158_n119022# w_n358_n132787# 0.240254f
C1663 a_n158_n18530# a_n158_n17494# 0.010536f
C1664 a_100_n68258# a_100_n67222# 0.010536f
C1665 a_n100_n16555# a_n100_n17591# 0.205388f
C1666 a_n100_n18627# a_n100_n19663# 0.205388f
C1667 a_n158_86106# a_n100_86009# 0.090922f
C1668 a_n100_66325# a_n100_65289# 0.205388f
C1669 a_n100_37317# w_n358_n132787# 0.269531f
C1670 a_100_6334# a_100_5298# 0.010536f
C1671 a_n100_5201# a_n158_5298# 0.090922f
C1672 a_100_53990# w_n358_n132787# 0.240254f
C1673 a_n100_n37275# a_n158_n37178# 0.090922f
C1674 a_100_71602# a_100_70566# 0.010536f
C1675 a_n158_46738# w_n358_n132787# 0.240254f
C1676 a_100_n122130# a_100_n123166# 0.010536f
C1677 a_n100_n123263# a_n158_n123166# 0.090922f
C1678 a_n100_n10339# a_n100_n9303# 0.205388f
C1679 a_n158_n108662# a_100_n108662# 0.219309f
C1680 a_n158_35342# a_100_35342# 0.219309f
C1681 a_100_n109698# w_n358_n132787# 0.240254f
C1682 a_n158_107862# w_n358_n132787# 0.240254f
C1683 a_100_68494# a_100_69530# 0.010536f
C1684 a_n100_89117# a_n158_89214# 0.090922f
C1685 a_n100_n66283# a_n100_n65247# 0.205388f
C1686 a_n158_n92086# w_n358_n132787# 0.240254f
C1687 a_n100_n32095# a_n100_n31059# 0.205388f
C1688 a_n158_105790# a_n158_104754# 0.010536f
C1689 a_n100_n82859# a_n158_n82762# 0.090922f
C1690 a_n158_n103482# w_n358_n132787# 0.240254f
C1691 w_n358_n132787# a_n158_n71366# 0.240254f
C1692 a_n158_23946# a_100_23946# 0.219309f
C1693 a_100_30162# w_n358_n132787# 0.240254f
C1694 a_n100_n51779# w_n358_n132787# 0.269531f
C1695 a_n158_n19566# a_100_n19566# 0.219309f
C1696 a_n100_n19663# a_n100_n20699# 0.205388f
C1697 a_n158_n105554# a_100_n105554# 0.219309f
C1698 a_n100_n91147# a_n100_n92183# 0.205388f
C1699 a_100_n126274# a_n158_n126274# 0.219309f
C1700 a_n100_n127407# a_n100_n126371# 0.205388f
C1701 a_n158_129618# a_n158_130654# 0.010536f
C1702 a_n158_n103482# a_n100_n103579# 0.090922f
C1703 a_100_45702# a_100_46738# 0.010536f
C1704 a_n100_n107723# w_n358_n132787# 0.269531f
C1705 a_n158_126510# a_100_126510# 0.219309f
C1706 a_100_77818# w_n358_n132787# 0.240254f
C1707 a_n100_n59031# a_n158_n58934# 0.090922f
C1708 a_n100_n62139# w_n358_n132787# 0.269531f
C1709 a_n100_10381# w_n358_n132787# 0.269531f
C1710 a_n158_86106# a_n158_87142# 0.010536f
C1711 a_n158_66422# a_n100_66325# 0.090922f
C1712 a_100_89214# a_n158_89214# 0.219309f
C1713 a_n158_n67222# a_n158_n66186# 0.010536f
C1714 a_n100_n76643# a_100_n76546# 0.090922f
C1715 a_n100_98441# a_n100_97405# 0.205388f
C1716 a_n100_n60067# a_100_n59970# 0.090922f
C1717 a_n100_n46599# a_100_n46502# 0.090922f
C1718 a_n100_n73535# w_n358_n132787# 0.269531f
C1719 a_100_76782# a_n100_76685# 0.090922f
C1720 a_100_87142# a_100_88178# 0.010536f
C1721 a_100_8406# a_100_7370# 0.010536f
C1722 a_n100_7273# a_n158_7370# 0.090922f
C1723 a_n158_106826# w_n358_n132787# 0.240254f
C1724 a_100_n39250# w_n358_n132787# 0.240254f
C1725 a_n100_n110831# a_100_n110734# 0.090922f
C1726 a_n100_74613# a_n100_75649# 0.205388f
C1727 a_100_n64114# a_100_n63078# 0.010536f
C1728 a_n158_n56862# a_100_n56862# 0.219309f
C1729 a_100_88178# a_n158_88178# 0.219309f
C1730 a_n158_n129382# a_n158_n130418# 0.010536f
C1731 a_n100_102585# w_n358_n132787# 0.269531f
C1732 a_100_n94158# a_100_n93122# 0.010536f
C1733 a_n158_21874# w_n358_n132787# 0.240254f
C1734 a_n158_37414# a_100_37414# 0.219309f
C1735 a_100_117186# w_n358_n132787# 0.240254f
C1736 a_n100_n28987# w_n358_n132787# 0.269531f
C1737 a_n158_80926# a_n100_80829# 0.090922f
C1738 a_n100_59073# a_n158_59170# 0.090922f
C1739 a_n100_12453# a_100_12550# 0.090922f
C1740 a_n158_103718# w_n358_n132787# 0.240254f
C1741 a_n100_118125# a_n100_117089# 0.205388f
C1742 a_n158_78854# a_n158_77818# 0.010536f
C1743 a_n100_96369# a_n100_97405# 0.205388f
C1744 a_n100_26957# a_n100_25921# 0.205388f
C1745 a_n158_n81726# w_n358_n132787# 0.240254f
C1746 a_n158_35342# w_n358_n132787# 0.240254f
C1747 w_n358_n132787# a_n100_n122227# 0.269531f
C1748 a_n158_n16458# a_100_n16458# 0.219309f
C1749 a_n158_109934# w_n358_n132787# 0.240254f
C1750 a_n100_4165# a_n158_4262# 0.090922f
C1751 a_n100_67361# a_100_67458# 0.090922f
C1752 a_n158_14622# w_n358_n132787# 0.240254f
C1753 a_n100_127449# a_n100_128485# 0.205388f
C1754 a_n158_n87942# a_100_n87942# 0.219309f
C1755 a_n100_54929# w_n358_n132787# 0.269531f
C1756 a_n100_33173# a_n158_33270# 0.090922f
C1757 a_100_n14386# a_100_n15422# 0.010536f
C1758 a_100_n33034# w_n358_n132787# 0.240254f
C1759 a_n100_9345# a_n158_9442# 0.090922f
C1760 a_100_n918# w_n358_n132787# 0.240254f
C1761 a_100_n31998# a_100_n33034# 0.010536f
C1762 a_100_n68258# a_n158_n68258# 0.219309f
C1763 a_100_n128346# w_n358_n132787# 0.240254f
C1764 a_n158_101646# a_n158_100610# 0.010536f
C1765 a_n100_n11375# w_n358_n132787# 0.269531f
C1766 a_n100_n20699# a_n158_n20602# 0.090922f
C1767 a_n100_22813# a_n100_21777# 0.205388f
C1768 a_100_108898# w_n358_n132787# 0.240254f
C1769 a_100_96466# a_100_95430# 0.010536f
C1770 a_n158_27054# w_n358_n132787# 0.240254f
C1771 a_n100_1057# a_n158_1154# 0.090922f
C1772 a_n100_40425# a_100_40522# 0.090922f
C1773 a_n100_81865# a_n100_80829# 0.205388f
C1774 a_n100_n22771# w_n358_n132787# 0.269531f
C1775 a_100_n90014# w_n358_n132787# 0.240254f
C1776 a_n158_n64114# a_n100_n64211# 0.090922f
C1777 a_n100_89117# w_n358_n132787# 0.269531f
C1778 a_100_n97266# a_100_n98302# 0.010536f
C1779 a_100_122366# a_100_121330# 0.010536f
C1780 a_n158_n43394# w_n358_n132787# 0.240254f
C1781 a_100_n15422# a_100_n16458# 0.010536f
C1782 a_n100_6237# a_n158_6334# 0.090922f
C1783 a_n100_51821# a_n158_51918# 0.090922f
C1784 a_100_n9206# a_100_n8170# 0.010536f
C1785 a_n100_n99435# a_100_n99338# 0.090922f
C1786 a_n100_n54887# a_n100_n55923# 0.205388f
C1787 a_100_99574# a_100_98538# 0.010536f
C1788 a_n100_98441# a_100_98538# 0.090922f
C1789 a_n100_51821# w_n358_n132787# 0.269531f
C1790 a_100_n22674# a_n100_n22771# 0.090922f
C1791 a_100_68494# a_100_67458# 0.010536f
C1792 a_100_n100374# a_n100_n100471# 0.090922f
C1793 a_100_81962# w_n358_n132787# 0.240254f
C1794 a_n158_n31998# w_n358_n132787# 0.240254f
C1795 a_100_89214# w_n358_n132787# 0.240254f
C1796 a_n158_3226# w_n358_n132787# 0.240254f
C1797 a_n158_n31998# a_100_n31998# 0.219309f
C1798 a_100_110970# a_100_112006# 0.010536f
C1799 a_100_n87942# a_100_n88978# 0.010536f
C1800 a_100_123402# a_100_124438# 0.010536f
C1801 a_n158_65386# w_n358_n132787# 0.240254f
C1802 a_n100_129521# a_n100_130557# 0.205388f
C1803 a_100_26018# a_100_24982# 0.010536f
C1804 a_n100_24885# a_n158_24982# 0.090922f
C1805 a_n100_n97363# a_n100_n96327# 0.205388f
C1806 a_n100_n48671# w_n358_n132787# 0.269531f
C1807 a_n158_3226# a_100_3226# 0.219309f
C1808 a_100_93358# w_n358_n132787# 0.240254f
C1809 a_n158_55026# a_n158_53990# 0.010536f
C1810 a_n158_103718# a_100_103718# 0.219309f
C1811 a_n100_102585# a_n100_103621# 0.205388f
C1812 a_n100_n40383# a_n158_n40286# 0.090922f
C1813 a_n100_n82859# w_n358_n132787# 0.269531f
C1814 a_n100_44569# w_n358_n132787# 0.269531f
C1815 a_100_55026# a_100_53990# 0.010536f
C1816 a_n158_n117986# w_n358_n132787# 0.240254f
C1817 a_100_n58934# a_100_n57898# 0.010536f
C1818 a_n158_n26818# a_n158_n27854# 0.010536f
C1819 a_100_n91050# w_n358_n132787# 0.240254f
C1820 a_100_n6098# a_100_n7134# 0.010536f
C1821 a_100_n69294# a_n100_n69391# 0.090922f
C1822 a_n158_13586# w_n358_n132787# 0.240254f
C1823 a_n158_103718# a_n100_103621# 0.090922f
C1824 a_n100_32137# a_100_32234# 0.090922f
C1825 a_n100_n48671# a_n158_n48574# 0.090922f
C1826 a_n100_67361# w_n358_n132787# 0.269531f
C1827 a_n158_n37178# w_n358_n132787# 0.240254f
C1828 a_n158_n13350# a_n158_n14386# 0.010536f
C1829 a_n158_96466# a_n158_95430# 0.010536f
C1830 a_n100_59073# a_n100_58037# 0.205388f
C1831 a_n100_n35203# a_100_n35106# 0.090922f
C1832 a_n100_124341# w_n358_n132787# 0.269531f
C1833 a_n100_8309# a_100_8406# 0.090922f
C1834 a_n158_n95194# a_100_n95194# 0.219309f
C1835 a_100_130654# a_100_129618# 0.010536f
C1836 a_n100_63217# w_n358_n132787# 0.269531f
C1837 a_n158_105790# a_n100_105693# 0.090922f
C1838 a_n158_n79654# w_n358_n132787# 0.240254f
C1839 a_n100_57001# a_n100_58037# 0.205388f
C1840 a_n100_44569# a_n158_44666# 0.090922f
C1841 a_100_23946# w_n358_n132787# 0.240254f
C1842 a_n158_n119022# a_100_n119022# 0.219309f
C1843 a_100_n86906# w_n358_n132787# 0.240254f
C1844 a_n158_n8170# a_n158_n9206# 0.010536f
C1845 a_100_n74474# w_n358_n132787# 0.240254f
C1846 a_n158_81962# a_n158_82998# 0.010536f
C1847 a_n158_n95194# w_n358_n132787# 0.240254f
C1848 a_n100_n28987# a_n158_n28890# 0.090922f
C1849 a_n100_71505# a_n158_71602# 0.090922f
C1850 a_100_106826# w_n358_n132787# 0.240254f
C1851 a_n100_48713# w_n358_n132787# 0.269531f
C1852 a_100_29126# a_100_28090# 0.010536f
C1853 a_n100_27993# a_n158_28090# 0.090922f
C1854 a_n158_n18530# a_100_n18530# 0.219309f
C1855 a_n158_n41322# w_n358_n132787# 0.240254f
C1856 a_100_37414# w_n358_n132787# 0.240254f
C1857 a_n100_5201# a_100_5298# 0.090922f
C1858 a_n158_n62042# a_n158_n61006# 0.010536f
C1859 a_n158_105790# w_n358_n132787# 0.240254f
C1860 a_n100_n60067# a_n158_n59970# 0.090922f
C1861 a_n158_n56862# a_n158_n57898# 0.010536f
C1862 a_n158_n22674# a_n100_n22771# 0.090922f
C1863 a_n100_110873# w_n358_n132787# 0.269531f
C1864 a_100_46738# w_n358_n132787# 0.240254f
C1865 a_n158_n125238# a_100_n125238# 0.219309f
C1866 a_n100_n125335# a_n100_n126371# 0.205388f
C1867 a_n158_79890# a_100_79890# 0.219309f
C1868 a_100_17730# w_n358_n132787# 0.240254f
C1869 a_n158_106826# a_n100_106729# 0.090922f
C1870 a_n100_n8267# a_n100_n9303# 0.205388f
C1871 a_100_n2990# a_100_n4026# 0.010536f
C1872 a_n100_69433# a_n158_69530# 0.090922f
C1873 a_n100_n129479# a_100_n129382# 0.090922f
C1874 a_n158_n109698# a_n158_n110734# 0.010536f
C1875 a_100_68494# w_n358_n132787# 0.240254f
C1876 a_n158_10478# a_100_10478# 0.219309f
C1877 a_n158_1154# w_n358_n132787# 0.240254f
C1878 a_100_64350# a_100_65386# 0.010536f
C1879 a_100_105790# a_n100_105693# 0.090922f
C1880 w_n358_n132787# a_100_n107626# 0.240254f
C1881 a_n158_n63078# w_n358_n132787# 0.240254f
C1882 a_n100_23849# a_n100_22813# 0.205388f
C1883 a_n100_29029# w_n358_n132787# 0.269531f
C1884 a_n100_n40383# a_n100_n41419# 0.205388f
C1885 a_100_45702# a_n100_45605# 0.090922f
C1886 a_n100_82901# w_n358_n132787# 0.269531f
C1887 a_n100_93261# w_n358_n132787# 0.269531f
C1888 a_n158_n38214# a_n158_n39250# 0.010536f
C1889 a_n158_n71366# a_n100_n71463# 0.090922f
C1890 a_n100_55965# a_100_56062# 0.090922f
C1891 a_n158_74710# w_n358_n132787# 0.240254f
C1892 w_n358_n132787# a_n100_n121191# 0.269531f
C1893 a_100_76782# a_100_75746# 0.010536f
C1894 a_n158_60206# a_n158_61242# 0.010536f
C1895 a_n158_63314# a_n158_64350# 0.010536f
C1896 a_n100_49749# a_n100_50785# 0.205388f
C1897 a_n158_31198# a_100_31198# 0.219309f
C1898 a_n100_31101# a_n100_30065# 0.205388f
C1899 a_n100_7273# a_100_7370# 0.090922f
C1900 a_100_n112806# a_100_n113842# 0.010536f
C1901 a_n100_n113939# a_n158_n113842# 0.090922f
C1902 a_100_55026# a_n100_54929# 0.090922f
C1903 a_100_105790# w_n358_n132787# 0.240254f
C1904 a_n158_n40286# w_n358_n132787# 0.240254f
C1905 a_100_n131454# a_100_n132490# 0.010536f
C1906 a_n100_n132587# a_n158_n132490# 0.090922f
C1907 a_n100_91189# a_n100_90153# 0.205388f
C1908 a_n158_93358# w_n358_n132787# 0.240254f
C1909 a_n158_20838# a_n158_19802# 0.010536f
C1910 a_100_21874# w_n358_n132787# 0.240254f
C1911 a_n100_n56959# w_n358_n132787# 0.269531f
C1912 a_100_n127310# w_n358_n132787# 0.240254f
C1913 a_100_129618# w_n358_n132787# 0.240254f
C1914 a_n100_37317# a_n100_36281# 0.205388f
C1915 a_n100_118125# a_100_118222# 0.090922f
C1916 a_n158_5298# w_n358_n132787# 0.240254f
C1917 a_100_108898# a_n100_108801# 0.090922f
C1918 a_n100_34209# w_n358_n132787# 0.269531f
C1919 a_n158_n16458# a_n158_n17494# 0.010536f
C1920 a_n100_n45563# w_n358_n132787# 0.269531f
C1921 a_n100_4165# a_100_4262# 0.090922f
C1922 a_n158_62278# a_n158_61242# 0.010536f
C1923 a_n100_79793# w_n358_n132787# 0.269531f
C1924 a_100_66422# a_n100_66325# 0.090922f
C1925 a_100_97502# w_n358_n132787# 0.240254f
C1926 a_100_n19566# w_n358_n132787# 0.240254f
C1927 a_100_14622# w_n358_n132787# 0.240254f
C1928 a_n158_n58934# w_n358_n132787# 0.240254f
C1929 a_n158_n114878# w_n358_n132787# 0.240254f
C1930 a_n158_n59970# a_n158_n61006# 0.010536f
C1931 a_n100_n15519# a_n158_n15422# 0.090922f
C1932 a_n100_33173# a_100_33270# 0.090922f
C1933 a_100_127546# w_n358_n132787# 0.240254f
C1934 a_n100_9345# a_n100_8309# 0.205388f
C1935 a_n158_n6098# a_n100_n6195# 0.090922f
C1936 a_n100_n2051# w_n358_n132787# 0.269531f
C1937 a_n158_96466# a_n158_97502# 0.010536f
C1938 a_100_n52718# a_100_n53754# 0.010536f
C1939 a_n158_n11278# w_n358_n132787# 0.240254f
C1940 a_100_61242# a_n158_61242# 0.219309f
C1941 a_n100_n116011# a_n158_n115914# 0.090922f
C1942 a_n158_1154# a_100_1154# 0.219309f
C1943 a_100_93358# a_100_92322# 0.010536f
C1944 a_100_27054# w_n358_n132787# 0.240254f
C1945 a_n158_40522# a_100_40522# 0.219309f
C1946 a_n100_40425# a_n100_39389# 0.205388f
C1947 a_n158_n104518# a_n158_n105554# 0.010536f
C1948 a_100_n25782# w_n358_n132787# 0.240254f
C1949 a_100_n93122# w_n358_n132787# 0.240254f
C1950 a_n158_n116950# w_n358_n132787# 0.240254f
C1951 a_100_40522# w_n358_n132787# 0.240254f
C1952 a_n100_n41419# w_n358_n132787# 0.269531f
C1953 a_n100_90153# w_n358_n132787# 0.269531f
C1954 a_n158_n90014# w_n358_n132787# 0.240254f
C1955 a_n100_n14483# w_n358_n132787# 0.269531f
C1956 a_100_n55826# a_n100_n55923# 0.090922f
C1957 a_n100_n23807# a_n100_n22771# 0.205388f
C1958 a_n100_18669# w_n358_n132787# 0.269531f
C1959 a_100_n121094# a_100_n122130# 0.010536f
C1960 a_n100_n122227# a_n158_n122130# 0.090922f
C1961 a_100_n108662# w_n358_n132787# 0.240254f
C1962 a_n158_73674# w_n358_n132787# 0.240254f
C1963 a_n158_131690# a_n158_130654# 0.010536f
C1964 a_n158_11514# a_n158_10478# 0.010536f
C1965 a_100_80926# a_100_79890# 0.010536f
C1966 a_n100_42497# a_n100_41461# 0.205388f
C1967 a_n100_75649# a_n158_75746# 0.090922f
C1968 a_100_75746# a_n158_75746# 0.219309f
C1969 a_n158_n88978# w_n358_n132787# 0.240254f
C1970 a_n158_112006# a_n158_110970# 0.010536f
C1971 a_n158_n49610# a_n158_n50646# 0.010536f
C1972 a_n158_n69294# a_n158_n70330# 0.010536f
C1973 a_100_n66186# w_n358_n132787# 0.240254f
C1974 a_100_n48574# w_n358_n132787# 0.240254f
C1975 a_n158_118222# w_n358_n132787# 0.240254f
C1976 a_n100_n106687# a_100_n106590# 0.090922f
C1977 a_n100_120197# a_100_120294# 0.090922f
C1978 a_100_106826# a_n100_106729# 0.090922f
C1979 a_100_127546# a_100_126510# 0.010536f
C1980 a_n158_57098# a_n100_57001# 0.090922f
C1981 a_n158_n87942# w_n358_n132787# 0.240254f
C1982 a_100_n66186# a_100_n67222# 0.010536f
C1983 a_100_n25782# a_n100_n25879# 0.090922f
C1984 a_100_13586# w_n358_n132787# 0.240254f
C1985 a_n158_n48574# a_100_n48574# 0.219309f
C1986 a_n100_121233# a_n100_122269# 0.205388f
C1987 a_n158_60206# a_n100_60109# 0.090922f
C1988 a_n100_8309# a_n100_7273# 0.205388f
C1989 a_n158_n35106# a_100_n35106# 0.219309f
C1990 a_n158_115114# w_n358_n132787# 0.240254f
C1991 a_n158_n128346# a_n158_n129382# 0.010536f
C1992 a_n158_n78618# a_n100_n78715# 0.090922f
C1993 a_n158_n79654# a_100_n79654# 0.219309f
C1994 a_100_45702# a_100_44666# 0.010536f
C1995 a_n100_n52815# w_n358_n132787# 0.269531f
C1996 a_n158_n20602# a_n158_n21638# 0.010536f
C1997 a_n158_118# a_n158_n918# 0.010536f
C1998 a_100_39486# a_100_38450# 0.010536f
C1999 a_n100_n64211# w_n358_n132787# 0.269531f
C2000 a_100_100610# a_n100_100513# 0.090922f
C2001 a_n100_13489# a_n100_12453# 0.205388f
C2002 a_n158_102682# a_n100_102585# 0.090922f
C2003 a_n100_109837# w_n358_n132787# 0.269531f
C2004 a_n158_n6098# w_n358_n132787# 0.240254f
C2005 a_n100_n91147# a_n158_n91050# 0.090922f
C2006 a_n100_115017# w_n358_n132787# 0.269531f
C2007 a_n158_48810# w_n358_n132787# 0.240254f
C2008 a_n100_27993# a_n100_26957# 0.205388f
C2009 w_n358_n132787# a_n100_n120155# 0.269531f
C2010 a_100_n41322# w_n358_n132787# 0.240254f
C2011 a_n158_103718# a_n158_102682# 0.010536f
C2012 a_n158_49846# a_100_49846# 0.219309f
C2013 a_n158_92322# a_n100_92225# 0.090922f
C2014 a_100_n78618# a_100_n77582# 0.010536f
C2015 a_n100_45605# w_n358_n132787# 0.269531f
C2016 a_100_n23710# a_100_n24746# 0.010536f
C2017 a_n158_n78618# w_n358_n132787# 0.240254f
C2018 a_n100_n10339# a_100_n10242# 0.090922f
C2019 a_n100_n55923# w_n358_n132787# 0.269531f
C2020 a_n100_16597# w_n358_n132787# 0.269531f
C2021 a_100_130654# a_n100_130557# 0.090922f
C2022 a_n100_n31059# w_n358_n132787# 0.269531f
C2023 a_100_n126274# w_n358_n132787# 0.240254f
C2024 a_n100_n35203# a_n158_n35106# 0.090922f
C2025 a_100_n88978# w_n358_n132787# 0.240254f
C2026 a_n100_82901# a_n100_83937# 0.205388f
C2027 a_n158_52954# a_n158_53990# 0.010536f
C2028 a_100_n86906# a_100_n85870# 0.010536f
C2029 a_n158_128582# w_n358_n132787# 0.240254f
C2030 a_n100_87045# a_n100_86009# 0.205388f
C2031 a_n158_94394# a_100_94394# 0.219309f
C2032 a_100_n51682# a_100_n52718# 0.010536f
C2033 a_n158_23946# a_n158_22910# 0.010536f
C2034 a_n100_n74571# a_n100_n75607# 0.205388f
C2035 a_n100_n49707# w_n358_n132787# 0.269531f
C2036 a_n158_29126# w_n358_n132787# 0.240254f
C2037 a_100_42594# a_100_41558# 0.010536f
C2038 w_n358_n132787# a_100_n125238# 0.240254f
C2039 a_n158_n65150# a_n100_n65247# 0.090922f
C2040 a_n158_31198# a_n158_30162# 0.010536f
C2041 a_100_99574# w_n358_n132787# 0.240254f
C2042 a_n158_n78618# a_n158_n77582# 0.010536f
C2043 a_n158_n59970# a_100_n59970# 0.219309f
C2044 a_n100_n107723# a_n100_n108759# 0.205388f
C2045 a_n158_125474# a_100_125474# 0.219309f
C2046 a_n158_n80690# a_n100_n80787# 0.090922f
C2047 a_n100_115017# a_n100_116053# 0.205388f
C2048 a_100_n62042# a_n158_n62042# 0.219309f
C2049 a_n100_n63175# a_n100_n62139# 0.205388f
C2050 a_n100_7273# a_n100_6237# 0.205388f
C2051 a_n100_98441# w_n358_n132787# 0.269531f
C2052 w_n358_n132787# a_n100_n61103# 0.269531f
C2053 a_100_n82762# a_100_n83798# 0.010536f
C2054 a_100_109934# a_100_110970# 0.010536f
C2055 a_100_n69294# a_100_n70330# 0.010536f
C2056 a_100_120294# a_100_119258# 0.010536f
C2057 a_n100_n93219# w_n358_n132787# 0.269531f
C2058 a_n158_n73438# a_n158_n74474# 0.010536f
C2059 a_n158_n14386# w_n358_n132787# 0.240254f
C2060 a_100_n55826# a_n158_n55826# 0.219309f
C2061 a_n100_76685# a_n100_77721# 0.205388f
C2062 a_n158_n113842# w_n358_n132787# 0.240254f
C2063 a_100_n101410# w_n358_n132787# 0.240254f
C2064 a_n158_n132490# w_n358_n132787# 0.244798f
C2065 a_n100_99477# a_n100_100513# 0.205388f
C2066 a_n158_61242# w_n358_n132787# 0.240254f
C2067 a_100_52954# a_100_51918# 0.010536f
C2068 a_100_n42358# a_100_n43394# 0.010536f
C2069 a_100_n28890# w_n358_n132787# 0.240254f
C2070 a_n100_87045# a_n158_87142# 0.090922f
C2071 a_n100_n11375# a_100_n11278# 0.090922f
C2072 a_n100_n83895# w_n358_n132787# 0.269531f
C2073 a_100_5298# w_n358_n132787# 0.240254f
C2074 a_n158_27054# a_n158_26018# 0.010536f
C2075 a_n158_n45466# w_n358_n132787# 0.240254f
C2076 a_n158_34306# w_n358_n132787# 0.240254f
C2077 a_n100_96369# w_n358_n132787# 0.269531f
C2078 a_n158_4262# a_100_4262# 0.219309f
C2079 a_n158_72638# a_n100_72541# 0.090922f
C2080 a_n158_n115914# w_n358_n132787# 0.240254f
C2081 a_n158_53990# w_n358_n132787# 0.240254f
C2082 a_n100_n60067# a_n100_n59031# 0.205388f
C2083 a_n158_33270# a_100_33270# 0.219309f
C2084 a_n100_33173# a_n100_32137# 0.205388f
C2085 w_n358_n132787# a_100_n69294# 0.240254f
C2086 a_n100_n15519# a_100_n15422# 0.090922f
C2087 a_100_48810# w_n358_n132787# 0.240254f
C2088 w_n358_n132787# a_n100_130557# 0.269531f
C2089 a_n100_131593# a_100_131690# 0.090922f
C2090 a_n158_57098# a_100_57098# 0.219309f
C2091 a_n158_n117986# a_100_n117986# 0.219309f
C2092 a_n100_n118083# a_n100_n119119# 0.205388f
C2093 a_n158_n73438# a_100_n73438# 0.219309f
C2094 a_n158_n94158# a_n158_n93122# 0.010536f
C2095 a_100_n105554# a_100_n106590# 0.010536f
C2096 a_100_84034# a_100_82998# 0.010536f
C2097 a_n100_n87003# a_100_n86906# 0.090922f
C2098 a_n100_74613# w_n358_n132787# 0.269531f
C2099 a_100_n26818# a_100_n27854# 0.010536f
C2100 a_100_9442# w_n358_n132787# 0.240254f
C2101 a_n158_n47538# a_n100_n47635# 0.090922f
C2102 a_n100_94297# a_n100_93261# 0.205388f
C2103 a_100_81962# a_100_80926# 0.010536f
C2104 a_n100_39389# w_n358_n132787# 0.269531f
C2105 a_n158_78854# w_n358_n132787# 0.240254f
C2106 a_100_n35106# a_100_n36142# 0.010536f
C2107 a_100_n17494# w_n358_n132787# 0.240254f
C2108 a_n100_n94255# a_n100_n93219# 0.205388f
C2109 a_n158_n124202# a_100_n124202# 0.219309f
C2110 a_n100_n124299# a_n100_n125335# 0.205388f
C2111 a_100_n109698# a_n100_n109795# 0.090922f
C2112 a_100_19802# a_100_18766# 0.010536f
C2113 a_n158_79890# a_n100_79793# 0.090922f
C2114 a_n158_n96230# a_n158_n95194# 0.010536f
C2115 a_n158_18766# w_n358_n132787# 0.240254f
C2116 a_n158_n55826# w_n358_n132787# 0.240254f
C2117 a_n100_80829# w_n358_n132787# 0.269531f
C2118 a_n100_n128443# a_100_n128346# 0.090922f
C2119 a_n100_73577# a_n158_73674# 0.090922f
C2120 a_n100_10381# a_n158_10478# 0.090922f
C2121 a_100_n28890# a_100_n29926# 0.010536f
C2122 a_n100_70469# a_n158_70566# 0.090922f
C2123 a_n100_24885# a_n100_23849# 0.205388f
C2124 a_n100_n65247# w_n358_n132787# 0.269531f
C2125 a_n158_n105554# w_n358_n132787# 0.240254f
C2126 a_n100_75649# a_n100_76685# 0.205388f
C2127 a_n100_n40383# a_100_n40286# 0.090922f
C2128 a_100_n98302# w_n358_n132787# 0.240254f
C2129 a_n158_15658# a_100_15658# 0.219309f
C2130 a_n100_15561# a_n100_14525# 0.205388f
C2131 a_100_44666# w_n358_n132787# 0.240254f
C2132 a_n158_n23710# w_n358_n132787# 0.240254f
C2133 a_n100_108801# a_n100_109837# 0.205388f
C2134 a_n100_50785# a_100_50882# 0.090922f
C2135 a_100_n58934# a_n158_n58934# 0.219309f
C2136 a_n100_101549# w_n358_n132787# 0.269531f
C2137 a_n158_47774# a_n158_46738# 0.010536f
C2138 a_n158_121330# w_n358_n132787# 0.240254f
C2139 a_100_n14386# a_n100_n14483# 0.090922f
C2140 a_100_n101410# a_100_n102446# 0.010536f
C2141 a_n100_120197# a_n100_121233# 0.205388f
C2142 a_n158_123402# a_100_123402# 0.219309f
C2143 a_100_n111770# a_100_n112806# 0.010536f
C2144 a_n100_n112903# a_n158_n112806# 0.090922f
C2145 a_n158_114078# a_100_114078# 0.219309f
C2146 a_100_n130418# a_100_n131454# 0.010536f
C2147 a_n100_n131551# a_n158_n131454# 0.090922f
C2148 a_n158_n35106# a_n158_n36142# 0.010536f
C2149 a_100_n34070# a_n100_n34167# 0.090922f
C2150 a_100_n92086# w_n358_n132787# 0.240254f
C2151 a_n100_67361# a_n100_66325# 0.205388f
C2152 a_n158_n119022# a_n158_n120058# 0.010536f
C2153 a_n158_21874# a_n158_20838# 0.010536f
C2154 a_n158_n53754# a_n158_n54790# 0.010536f
C2155 a_n158_44666# a_100_44666# 0.219309f
C2156 a_n100_44569# a_n100_43533# 0.205388f
C2157 a_n158_22910# w_n358_n132787# 0.240254f
C2158 a_n158_n43394# a_n158_n42358# 0.010536f
C2159 a_n100_n43491# a_100_n43394# 0.090922f
C2160 a_n158_38450# a_100_38450# 0.219309f
C2161 a_n100_n41419# a_n100_n42455# 0.205388f
C2162 a_n100_n1015# a_n158_n918# 0.090922f
C2163 a_n100_n9303# a_n158_n9206# 0.090922f
C2164 a_n158_n102446# a_n158_n101410# 0.010536f
C2165 a_n158_n25782# w_n358_n132787# 0.240254f
C2166 a_n100_111909# a_100_112006# 0.090922f
C2167 a_n158_n28890# a_100_n28890# 0.219309f
C2168 a_n100_n80787# a_100_n80690# 0.090922f
C2169 a_100_95430# a_n158_95430# 0.219309f
C2170 a_n100_60109# w_n358_n132787# 0.269531f
C2171 w_n358_n132787# a_100_n124202# 0.240254f
C2172 a_n158_n97266# a_n158_n98302# 0.010536f
C2173 a_n158_n37178# a_100_n37178# 0.219309f
C2174 a_n100_88081# w_n358_n132787# 0.269531f
C2175 a_n100_n17591# w_n358_n132787# 0.269531f
C2176 a_n100_123305# a_n100_122269# 0.205388f
C2177 a_n158_16694# w_n358_n132787# 0.240254f
C2178 a_n158_n131454# w_n358_n132787# 0.240254f
C2179 a_n100_n45563# a_100_n45466# 0.090922f
C2180 a_n158_n112806# w_n358_n132787# 0.240254f
C2181 a_100_35342# a_100_34306# 0.010536f
C2182 a_n100_95333# w_n358_n132787# 0.269531f
C2183 a_n158_n12314# a_n158_n13350# 0.010536f
C2184 a_100_n34070# w_n358_n132787# 0.240254f
C2185 a_100_97502# a_100_96466# 0.010536f
C2186 a_n100_78757# a_n100_79793# 0.205388f
C2187 a_100_78854# w_n358_n132787# 0.240254f
C2188 a_n158_n8170# w_n358_n132787# 0.240254f
C2189 a_n100_n52815# a_n158_n52718# 0.090922f
C2190 a_100_29126# w_n358_n132787# 0.240254f
C2191 a_n158_64350# w_n358_n132787# 0.240254f
C2192 a_n100_41461# a_n100_40425# 0.205388f
C2193 a_n158_n63078# a_n100_n63175# 0.090922f
C2194 a_n100_n92183# w_n358_n132787# 0.269531f
C2195 a_n158_n98302# w_n358_n132787# 0.240254f
C2196 a_n158_128582# a_n100_128485# 0.090922f
C2197 a_n100_123305# a_100_123402# 0.090922f
C2198 a_n100_n25879# a_n158_n25782# 0.090922f
C2199 a_100_n83798# a_100_n84834# 0.010536f
C2200 a_100_n47538# a_n100_n47635# 0.090922f
C2201 a_100_74710# a_100_75746# 0.010536f
C2202 a_n158_n15422# a_n158_n16458# 0.010536f
C2203 a_100_n40286# w_n358_n132787# 0.240254f
C2204 a_n100_77721# a_n158_77818# 0.090922f
C2205 a_n100_n10339# w_n358_n132787# 0.269531f
C2206 a_n100_127449# a_n158_127546# 0.090922f
C2207 a_n158_n101410# a_n158_n100374# 0.010536f
C2208 a_n100_n74571# w_n358_n132787# 0.269531f
C2209 a_n158_n105554# a_n158_n106590# 0.010536f
C2210 a_n158_n23710# a_n158_n22674# 0.010536f
C2211 a_100_n120058# a_100_n121094# 0.010536f
C2212 a_n100_n121191# a_n158_n121094# 0.090922f
C2213 a_n158_n56862# w_n358_n132787# 0.240254f
C2214 w_n358_n132787# a_n100_131593# 0.349164f
C2215 a_n158_n41322# a_n158_n42358# 0.010536f
C2216 a_n158_n11278# a_100_n11278# 0.219309f
C2217 a_100_n90014# a_n100_n90111# 0.090922f
C2218 a_n158_112006# w_n358_n132787# 0.240254f
C2219 a_n100_n30023# w_n358_n132787# 0.269531f
C2220 a_100_n61006# a_n100_n61103# 0.090922f
C2221 a_100_n50646# a_n158_n50646# 0.219309f
C2222 a_100_74710# a_100_73674# 0.010536f
C2223 a_100_34306# w_n358_n132787# 0.240254f
C2224 a_n158_101646# w_n358_n132787# 0.240254f
C2225 a_n158_n37178# a_n158_n38214# 0.010536f
C2226 a_100_17730# a_100_16694# 0.010536f
C2227 a_n158_66422# a_100_66422# 0.219309f
C2228 a_n100_n24843# a_100_n24746# 0.090922f
C2229 a_n158_n109698# a_n158_n108662# 0.010536f
C2230 a_n158_n15422# a_100_n15422# 0.219309f
C2231 a_100_100610# a_100_101646# 0.010536f
C2232 a_100_n14386# a_n158_n14386# 0.219309f
C2233 a_100_76782# w_n358_n132787# 0.240254f
C2234 a_100_61242# a_n100_61145# 0.090922f
C2235 a_n158_9442# a_100_9442# 0.219309f
C2236 a_n100_82901# a_n158_82998# 0.090922f
C2237 a_n100_47677# w_n358_n132787# 0.269531f
C2238 a_n100_n80787# w_n358_n132787# 0.269531f
C2239 a_n158_n127310# a_n158_n128346# 0.010536f
C2240 a_n158_n5062# a_100_n5062# 0.219309f
C2241 a_n158_n53754# a_100_n53754# 0.219309f
C2242 a_n100_n53851# a_n100_n54887# 0.205388f
C2243 a_n100_n12411# w_n358_n132787# 0.269531f
C2244 a_n158_n7134# a_n158_n6098# 0.010536f
C2245 a_n100_59073# w_n358_n132787# 0.269531f
C2246 a_100_26018# w_n358_n132787# 0.240254f
C2247 a_n158_n49610# w_n358_n132787# 0.240254f
C2248 a_100_86106# a_100_87142# 0.010536f
C2249 a_100_88178# w_n358_n132787# 0.240254f
C2250 a_100_n86906# a_n158_n86906# 0.219309f
C2251 a_n100_57001# w_n358_n132787# 0.269531f
C2252 a_n100_73577# a_n100_74613# 0.205388f
C2253 a_n158_n27854# a_100_n27854# 0.219309f
C2254 a_n158_8406# w_n358_n132787# 0.240254f
C2255 a_n158_66422# a_n158_67458# 0.010536f
C2256 a_n158_n48574# a_n158_n49610# 0.010536f
C2257 a_n100_29029# a_n100_27993# 0.205388f
C2258 a_100_n66186# a_100_n65150# 0.010536f
C2259 a_100_n38214# w_n358_n132787# 0.240254f
C2260 a_n158_n36142# a_100_n36142# 0.219309f
C2261 a_n100_118125# a_n158_118222# 0.090922f
C2262 a_100_64350# w_n358_n132787# 0.240254f
C2263 a_n100_68397# w_n358_n132787# 0.269531f
C2264 a_n100_n3087# a_100_n2990# 0.090922f
C2265 a_n100_n60067# w_n358_n132787# 0.269531f
C2266 a_100_n63078# a_n158_n63078# 0.219309f
C2267 a_n158_n99338# a_n158_n98302# 0.010536f
C2268 a_n158_36378# a_n158_35342# 0.010536f
C2269 a_100_82998# w_n358_n132787# 0.240254f
C2270 a_100_n43394# a_100_n44430# 0.010536f
C2271 a_n100_n73535# a_100_n73438# 0.090922f
C2272 a_100_n108662# a_n100_n108759# 0.090922f
C2273 a_n100_n100471# a_n158_n100374# 0.090922f
C2274 a_n158_121330# a_n158_122366# 0.010536f
C2275 a_n158_126510# a_n158_127546# 0.010536f
C2276 a_n100_75649# a_100_75746# 0.090922f
C2277 a_n158_n31998# a_n158_n30962# 0.010536f
C2278 a_n100_n30023# a_100_n29926# 0.090922f
C2279 a_n158_2190# w_n358_n132787# 0.240254f
C2280 a_100_107862# w_n358_n132787# 0.240254f
C2281 a_n158_n46502# w_n358_n132787# 0.240254f
C2282 a_n100_31101# w_n358_n132787# 0.269531f
C2283 a_n100_117089# a_n158_117186# 0.090922f
C2284 w_n358_n132787# a_100_n123166# 0.240254f
C2285 a_100_n100374# a_n158_n100374# 0.219309f
C2286 a_100_n23710# w_n358_n132787# 0.240254f
C2287 a_n100_n7231# a_n100_n8267# 0.205388f
C2288 a_n158_n114878# a_100_n114878# 0.219309f
C2289 a_n100_107765# a_n158_107862# 0.090922f
C2290 a_n158_8406# a_n158_7370# 0.010536f
C2291 a_n158_n130418# w_n358_n132787# 0.240254f
C2292 a_n158_n111770# w_n358_n132787# 0.240254f
C2293 a_n158_79890# a_n158_78854# 0.010536f
C2294 a_n158_114078# w_n358_n132787# 0.240254f
C2295 a_n158_125474# a_n158_124438# 0.010536f
C2296 a_100_n22674# a_100_n23710# 0.010536f
C2297 a_n100_n23807# a_n158_n23710# 0.090922f
C2298 a_100_118# a_100_n918# 0.010536f
C2299 a_n100_n43491# a_n100_n44527# 0.205388f
C2300 a_100_n75510# a_100_n74474# 0.010536f
C2301 a_100_n132490# VSUBS 0.196066f
C2302 a_n158_n132490# VSUBS 0.196066f
C2303 a_n100_n132587# VSUBS 0.260213f
C2304 a_100_n131454# VSUBS 0.190616f
C2305 a_n158_n131454# VSUBS 0.190616f
C2306 a_n100_n131551# VSUBS 0.216482f
C2307 a_100_n130418# VSUBS 0.190616f
C2308 a_n158_n130418# VSUBS 0.190616f
C2309 a_n100_n130515# VSUBS 0.216482f
C2310 a_100_n129382# VSUBS 0.190616f
C2311 a_n158_n129382# VSUBS 0.190616f
C2312 a_n100_n129479# VSUBS 0.216482f
C2313 a_100_n128346# VSUBS 0.190616f
C2314 a_n158_n128346# VSUBS 0.190616f
C2315 a_n100_n128443# VSUBS 0.216482f
C2316 a_100_n127310# VSUBS 0.190616f
C2317 a_n158_n127310# VSUBS 0.190616f
C2318 a_n100_n127407# VSUBS 0.216482f
C2319 a_100_n126274# VSUBS 0.190616f
C2320 a_n158_n126274# VSUBS 0.190616f
C2321 a_n100_n126371# VSUBS 0.216482f
C2322 a_100_n125238# VSUBS 0.190616f
C2323 a_n158_n125238# VSUBS 0.190616f
C2324 a_n100_n125335# VSUBS 0.216482f
C2325 a_100_n124202# VSUBS 0.190616f
C2326 a_n158_n124202# VSUBS 0.190616f
C2327 a_n100_n124299# VSUBS 0.216482f
C2328 a_100_n123166# VSUBS 0.190616f
C2329 a_n158_n123166# VSUBS 0.190616f
C2330 a_n100_n123263# VSUBS 0.216482f
C2331 a_100_n122130# VSUBS 0.190616f
C2332 a_n158_n122130# VSUBS 0.190616f
C2333 a_n100_n122227# VSUBS 0.216482f
C2334 a_100_n121094# VSUBS 0.190616f
C2335 a_n158_n121094# VSUBS 0.190616f
C2336 a_n100_n121191# VSUBS 0.216482f
C2337 a_100_n120058# VSUBS 0.190616f
C2338 a_n158_n120058# VSUBS 0.190616f
C2339 a_n100_n120155# VSUBS 0.216482f
C2340 a_100_n119022# VSUBS 0.190616f
C2341 a_n158_n119022# VSUBS 0.190616f
C2342 a_n100_n119119# VSUBS 0.216482f
C2343 a_100_n117986# VSUBS 0.190616f
C2344 a_n158_n117986# VSUBS 0.190616f
C2345 a_n100_n118083# VSUBS 0.216482f
C2346 a_100_n116950# VSUBS 0.190616f
C2347 a_n158_n116950# VSUBS 0.190616f
C2348 a_n100_n117047# VSUBS 0.216482f
C2349 a_100_n115914# VSUBS 0.190616f
C2350 a_n158_n115914# VSUBS 0.190616f
C2351 a_n100_n116011# VSUBS 0.216482f
C2352 a_100_n114878# VSUBS 0.190616f
C2353 a_n158_n114878# VSUBS 0.190616f
C2354 a_n100_n114975# VSUBS 0.216482f
C2355 a_100_n113842# VSUBS 0.190616f
C2356 a_n158_n113842# VSUBS 0.190616f
C2357 a_n100_n113939# VSUBS 0.216482f
C2358 a_100_n112806# VSUBS 0.190616f
C2359 a_n158_n112806# VSUBS 0.190616f
C2360 a_n100_n112903# VSUBS 0.216482f
C2361 a_100_n111770# VSUBS 0.190616f
C2362 a_n158_n111770# VSUBS 0.190616f
C2363 a_n100_n111867# VSUBS 0.216482f
C2364 a_100_n110734# VSUBS 0.190616f
C2365 a_n158_n110734# VSUBS 0.190616f
C2366 a_n100_n110831# VSUBS 0.216482f
C2367 a_100_n109698# VSUBS 0.190616f
C2368 a_n158_n109698# VSUBS 0.190616f
C2369 a_n100_n109795# VSUBS 0.216482f
C2370 a_100_n108662# VSUBS 0.190616f
C2371 a_n158_n108662# VSUBS 0.190616f
C2372 a_n100_n108759# VSUBS 0.216482f
C2373 a_100_n107626# VSUBS 0.190616f
C2374 a_n158_n107626# VSUBS 0.190616f
C2375 a_n100_n107723# VSUBS 0.216482f
C2376 a_100_n106590# VSUBS 0.190616f
C2377 a_n158_n106590# VSUBS 0.190616f
C2378 a_n100_n106687# VSUBS 0.216482f
C2379 a_100_n105554# VSUBS 0.190616f
C2380 a_n158_n105554# VSUBS 0.190616f
C2381 a_n100_n105651# VSUBS 0.216482f
C2382 a_100_n104518# VSUBS 0.190616f
C2383 a_n158_n104518# VSUBS 0.190616f
C2384 a_n100_n104615# VSUBS 0.216482f
C2385 a_100_n103482# VSUBS 0.190616f
C2386 a_n158_n103482# VSUBS 0.190616f
C2387 a_n100_n103579# VSUBS 0.216482f
C2388 a_100_n102446# VSUBS 0.190616f
C2389 a_n158_n102446# VSUBS 0.190616f
C2390 a_n100_n102543# VSUBS 0.216482f
C2391 a_100_n101410# VSUBS 0.190616f
C2392 a_n158_n101410# VSUBS 0.190616f
C2393 a_n100_n101507# VSUBS 0.216482f
C2394 a_100_n100374# VSUBS 0.190616f
C2395 a_n158_n100374# VSUBS 0.190616f
C2396 a_n100_n100471# VSUBS 0.216482f
C2397 a_100_n99338# VSUBS 0.190616f
C2398 a_n158_n99338# VSUBS 0.190616f
C2399 a_n100_n99435# VSUBS 0.216482f
C2400 a_100_n98302# VSUBS 0.190616f
C2401 a_n158_n98302# VSUBS 0.190616f
C2402 a_n100_n98399# VSUBS 0.216482f
C2403 a_100_n97266# VSUBS 0.190616f
C2404 a_n158_n97266# VSUBS 0.190616f
C2405 a_n100_n97363# VSUBS 0.216482f
C2406 a_100_n96230# VSUBS 0.190616f
C2407 a_n158_n96230# VSUBS 0.190616f
C2408 a_n100_n96327# VSUBS 0.216482f
C2409 a_100_n95194# VSUBS 0.190616f
C2410 a_n158_n95194# VSUBS 0.190616f
C2411 a_n100_n95291# VSUBS 0.216482f
C2412 a_100_n94158# VSUBS 0.190616f
C2413 a_n158_n94158# VSUBS 0.190616f
C2414 a_n100_n94255# VSUBS 0.216482f
C2415 a_100_n93122# VSUBS 0.190616f
C2416 a_n158_n93122# VSUBS 0.190616f
C2417 a_n100_n93219# VSUBS 0.216482f
C2418 a_100_n92086# VSUBS 0.190616f
C2419 a_n158_n92086# VSUBS 0.190616f
C2420 a_n100_n92183# VSUBS 0.216482f
C2421 a_100_n91050# VSUBS 0.190616f
C2422 a_n158_n91050# VSUBS 0.190616f
C2423 a_n100_n91147# VSUBS 0.216482f
C2424 a_100_n90014# VSUBS 0.190616f
C2425 a_n158_n90014# VSUBS 0.190616f
C2426 a_n100_n90111# VSUBS 0.216482f
C2427 a_100_n88978# VSUBS 0.190616f
C2428 a_n158_n88978# VSUBS 0.190616f
C2429 a_n100_n89075# VSUBS 0.216482f
C2430 a_100_n87942# VSUBS 0.190616f
C2431 a_n158_n87942# VSUBS 0.190616f
C2432 a_n100_n88039# VSUBS 0.216482f
C2433 a_100_n86906# VSUBS 0.190616f
C2434 a_n158_n86906# VSUBS 0.190616f
C2435 a_n100_n87003# VSUBS 0.216482f
C2436 a_100_n85870# VSUBS 0.190616f
C2437 a_n158_n85870# VSUBS 0.190616f
C2438 a_n100_n85967# VSUBS 0.216482f
C2439 a_100_n84834# VSUBS 0.190616f
C2440 a_n158_n84834# VSUBS 0.190616f
C2441 a_n100_n84931# VSUBS 0.216482f
C2442 a_100_n83798# VSUBS 0.190616f
C2443 a_n158_n83798# VSUBS 0.190616f
C2444 a_n100_n83895# VSUBS 0.216482f
C2445 a_100_n82762# VSUBS 0.190616f
C2446 a_n158_n82762# VSUBS 0.190616f
C2447 a_n100_n82859# VSUBS 0.216482f
C2448 a_100_n81726# VSUBS 0.190616f
C2449 a_n158_n81726# VSUBS 0.190616f
C2450 a_n100_n81823# VSUBS 0.216482f
C2451 a_100_n80690# VSUBS 0.190616f
C2452 a_n158_n80690# VSUBS 0.190616f
C2453 a_n100_n80787# VSUBS 0.216482f
C2454 a_100_n79654# VSUBS 0.190616f
C2455 a_n158_n79654# VSUBS 0.190616f
C2456 a_n100_n79751# VSUBS 0.216482f
C2457 a_100_n78618# VSUBS 0.190616f
C2458 a_n158_n78618# VSUBS 0.190616f
C2459 a_n100_n78715# VSUBS 0.216482f
C2460 a_100_n77582# VSUBS 0.190616f
C2461 a_n158_n77582# VSUBS 0.190616f
C2462 a_n100_n77679# VSUBS 0.216482f
C2463 a_100_n76546# VSUBS 0.190616f
C2464 a_n158_n76546# VSUBS 0.190616f
C2465 a_n100_n76643# VSUBS 0.216482f
C2466 a_100_n75510# VSUBS 0.190616f
C2467 a_n158_n75510# VSUBS 0.190616f
C2468 a_n100_n75607# VSUBS 0.216482f
C2469 a_100_n74474# VSUBS 0.190616f
C2470 a_n158_n74474# VSUBS 0.190616f
C2471 a_n100_n74571# VSUBS 0.216482f
C2472 a_100_n73438# VSUBS 0.190616f
C2473 a_n158_n73438# VSUBS 0.190616f
C2474 a_n100_n73535# VSUBS 0.216482f
C2475 a_100_n72402# VSUBS 0.190616f
C2476 a_n158_n72402# VSUBS 0.190616f
C2477 a_n100_n72499# VSUBS 0.216482f
C2478 a_100_n71366# VSUBS 0.190616f
C2479 a_n158_n71366# VSUBS 0.190616f
C2480 a_n100_n71463# VSUBS 0.216482f
C2481 a_100_n70330# VSUBS 0.190616f
C2482 a_n158_n70330# VSUBS 0.190616f
C2483 a_n100_n70427# VSUBS 0.216482f
C2484 a_100_n69294# VSUBS 0.190616f
C2485 a_n158_n69294# VSUBS 0.190616f
C2486 a_n100_n69391# VSUBS 0.216482f
C2487 a_100_n68258# VSUBS 0.190616f
C2488 a_n158_n68258# VSUBS 0.190616f
C2489 a_n100_n68355# VSUBS 0.216482f
C2490 a_100_n67222# VSUBS 0.190616f
C2491 a_n158_n67222# VSUBS 0.190616f
C2492 a_n100_n67319# VSUBS 0.216482f
C2493 a_100_n66186# VSUBS 0.190616f
C2494 a_n158_n66186# VSUBS 0.190616f
C2495 a_n100_n66283# VSUBS 0.216482f
C2496 a_100_n65150# VSUBS 0.190616f
C2497 a_n158_n65150# VSUBS 0.190616f
C2498 a_n100_n65247# VSUBS 0.216482f
C2499 a_100_n64114# VSUBS 0.190616f
C2500 a_n158_n64114# VSUBS 0.190616f
C2501 a_n100_n64211# VSUBS 0.216482f
C2502 a_100_n63078# VSUBS 0.190616f
C2503 a_n158_n63078# VSUBS 0.190616f
C2504 a_n100_n63175# VSUBS 0.216482f
C2505 a_100_n62042# VSUBS 0.190616f
C2506 a_n158_n62042# VSUBS 0.190616f
C2507 a_n100_n62139# VSUBS 0.216482f
C2508 a_100_n61006# VSUBS 0.190616f
C2509 a_n158_n61006# VSUBS 0.190616f
C2510 a_n100_n61103# VSUBS 0.216482f
C2511 a_100_n59970# VSUBS 0.190616f
C2512 a_n158_n59970# VSUBS 0.190616f
C2513 a_n100_n60067# VSUBS 0.216482f
C2514 a_100_n58934# VSUBS 0.190616f
C2515 a_n158_n58934# VSUBS 0.190616f
C2516 a_n100_n59031# VSUBS 0.216482f
C2517 a_100_n57898# VSUBS 0.190616f
C2518 a_n158_n57898# VSUBS 0.190616f
C2519 a_n100_n57995# VSUBS 0.216482f
C2520 a_100_n56862# VSUBS 0.190616f
C2521 a_n158_n56862# VSUBS 0.190616f
C2522 a_n100_n56959# VSUBS 0.216482f
C2523 a_100_n55826# VSUBS 0.190616f
C2524 a_n158_n55826# VSUBS 0.190616f
C2525 a_n100_n55923# VSUBS 0.216482f
C2526 a_100_n54790# VSUBS 0.190616f
C2527 a_n158_n54790# VSUBS 0.190616f
C2528 a_n100_n54887# VSUBS 0.216482f
C2529 a_100_n53754# VSUBS 0.190616f
C2530 a_n158_n53754# VSUBS 0.190616f
C2531 a_n100_n53851# VSUBS 0.216482f
C2532 a_100_n52718# VSUBS 0.190616f
C2533 a_n158_n52718# VSUBS 0.190616f
C2534 a_n100_n52815# VSUBS 0.216482f
C2535 a_100_n51682# VSUBS 0.190616f
C2536 a_n158_n51682# VSUBS 0.190616f
C2537 a_n100_n51779# VSUBS 0.216482f
C2538 a_100_n50646# VSUBS 0.190616f
C2539 a_n158_n50646# VSUBS 0.190616f
C2540 a_n100_n50743# VSUBS 0.216482f
C2541 a_100_n49610# VSUBS 0.190616f
C2542 a_n158_n49610# VSUBS 0.190616f
C2543 a_n100_n49707# VSUBS 0.216482f
C2544 a_100_n48574# VSUBS 0.190616f
C2545 a_n158_n48574# VSUBS 0.190616f
C2546 a_n100_n48671# VSUBS 0.216482f
C2547 a_100_n47538# VSUBS 0.190616f
C2548 a_n158_n47538# VSUBS 0.190616f
C2549 a_n100_n47635# VSUBS 0.216482f
C2550 a_100_n46502# VSUBS 0.190616f
C2551 a_n158_n46502# VSUBS 0.190616f
C2552 a_n100_n46599# VSUBS 0.216482f
C2553 a_100_n45466# VSUBS 0.190616f
C2554 a_n158_n45466# VSUBS 0.190616f
C2555 a_n100_n45563# VSUBS 0.216482f
C2556 a_100_n44430# VSUBS 0.190616f
C2557 a_n158_n44430# VSUBS 0.190616f
C2558 a_n100_n44527# VSUBS 0.216482f
C2559 a_100_n43394# VSUBS 0.190616f
C2560 a_n158_n43394# VSUBS 0.190616f
C2561 a_n100_n43491# VSUBS 0.216482f
C2562 a_100_n42358# VSUBS 0.190616f
C2563 a_n158_n42358# VSUBS 0.190616f
C2564 a_n100_n42455# VSUBS 0.216482f
C2565 a_100_n41322# VSUBS 0.190616f
C2566 a_n158_n41322# VSUBS 0.190616f
C2567 a_n100_n41419# VSUBS 0.216482f
C2568 a_100_n40286# VSUBS 0.190616f
C2569 a_n158_n40286# VSUBS 0.190616f
C2570 a_n100_n40383# VSUBS 0.216482f
C2571 a_100_n39250# VSUBS 0.190616f
C2572 a_n158_n39250# VSUBS 0.190616f
C2573 a_n100_n39347# VSUBS 0.216482f
C2574 a_100_n38214# VSUBS 0.190616f
C2575 a_n158_n38214# VSUBS 0.190616f
C2576 a_n100_n38311# VSUBS 0.216482f
C2577 a_100_n37178# VSUBS 0.190616f
C2578 a_n158_n37178# VSUBS 0.190616f
C2579 a_n100_n37275# VSUBS 0.216482f
C2580 a_100_n36142# VSUBS 0.190616f
C2581 a_n158_n36142# VSUBS 0.190616f
C2582 a_n100_n36239# VSUBS 0.216482f
C2583 a_100_n35106# VSUBS 0.190616f
C2584 a_n158_n35106# VSUBS 0.190616f
C2585 a_n100_n35203# VSUBS 0.216482f
C2586 a_100_n34070# VSUBS 0.190616f
C2587 a_n158_n34070# VSUBS 0.190616f
C2588 a_n100_n34167# VSUBS 0.216482f
C2589 a_100_n33034# VSUBS 0.190616f
C2590 a_n158_n33034# VSUBS 0.190616f
C2591 a_n100_n33131# VSUBS 0.216482f
C2592 a_100_n31998# VSUBS 0.190616f
C2593 a_n158_n31998# VSUBS 0.190616f
C2594 a_n100_n32095# VSUBS 0.216482f
C2595 a_100_n30962# VSUBS 0.190616f
C2596 a_n158_n30962# VSUBS 0.190616f
C2597 a_n100_n31059# VSUBS 0.216482f
C2598 a_100_n29926# VSUBS 0.190616f
C2599 a_n158_n29926# VSUBS 0.190616f
C2600 a_n100_n30023# VSUBS 0.216482f
C2601 a_100_n28890# VSUBS 0.190616f
C2602 a_n158_n28890# VSUBS 0.190616f
C2603 a_n100_n28987# VSUBS 0.216482f
C2604 a_100_n27854# VSUBS 0.190616f
C2605 a_n158_n27854# VSUBS 0.190616f
C2606 a_n100_n27951# VSUBS 0.216482f
C2607 a_100_n26818# VSUBS 0.190616f
C2608 a_n158_n26818# VSUBS 0.190616f
C2609 a_n100_n26915# VSUBS 0.216482f
C2610 a_100_n25782# VSUBS 0.190616f
C2611 a_n158_n25782# VSUBS 0.190616f
C2612 a_n100_n25879# VSUBS 0.216482f
C2613 a_100_n24746# VSUBS 0.190616f
C2614 a_n158_n24746# VSUBS 0.190616f
C2615 a_n100_n24843# VSUBS 0.216482f
C2616 a_100_n23710# VSUBS 0.190616f
C2617 a_n158_n23710# VSUBS 0.190616f
C2618 a_n100_n23807# VSUBS 0.216482f
C2619 a_100_n22674# VSUBS 0.190616f
C2620 a_n158_n22674# VSUBS 0.190616f
C2621 a_n100_n22771# VSUBS 0.216482f
C2622 a_100_n21638# VSUBS 0.190616f
C2623 a_n158_n21638# VSUBS 0.190616f
C2624 a_n100_n21735# VSUBS 0.216482f
C2625 a_100_n20602# VSUBS 0.190616f
C2626 a_n158_n20602# VSUBS 0.190616f
C2627 a_n100_n20699# VSUBS 0.216482f
C2628 a_100_n19566# VSUBS 0.190616f
C2629 a_n158_n19566# VSUBS 0.190616f
C2630 a_n100_n19663# VSUBS 0.216482f
C2631 a_100_n18530# VSUBS 0.190616f
C2632 a_n158_n18530# VSUBS 0.190616f
C2633 a_n100_n18627# VSUBS 0.216482f
C2634 a_100_n17494# VSUBS 0.190616f
C2635 a_n158_n17494# VSUBS 0.190616f
C2636 a_n100_n17591# VSUBS 0.216482f
C2637 a_100_n16458# VSUBS 0.190616f
C2638 a_n158_n16458# VSUBS 0.190616f
C2639 a_n100_n16555# VSUBS 0.216482f
C2640 a_100_n15422# VSUBS 0.190616f
C2641 a_n158_n15422# VSUBS 0.190616f
C2642 a_n100_n15519# VSUBS 0.216482f
C2643 a_100_n14386# VSUBS 0.190616f
C2644 a_n158_n14386# VSUBS 0.190616f
C2645 a_n100_n14483# VSUBS 0.216482f
C2646 a_100_n13350# VSUBS 0.190616f
C2647 a_n158_n13350# VSUBS 0.190616f
C2648 a_n100_n13447# VSUBS 0.216482f
C2649 a_100_n12314# VSUBS 0.190616f
C2650 a_n158_n12314# VSUBS 0.190616f
C2651 a_n100_n12411# VSUBS 0.216482f
C2652 a_100_n11278# VSUBS 0.190616f
C2653 a_n158_n11278# VSUBS 0.190616f
C2654 a_n100_n11375# VSUBS 0.216482f
C2655 a_100_n10242# VSUBS 0.190616f
C2656 a_n158_n10242# VSUBS 0.190616f
C2657 a_n100_n10339# VSUBS 0.216482f
C2658 a_100_n9206# VSUBS 0.190616f
C2659 a_n158_n9206# VSUBS 0.190616f
C2660 a_n100_n9303# VSUBS 0.216482f
C2661 a_100_n8170# VSUBS 0.190616f
C2662 a_n158_n8170# VSUBS 0.190616f
C2663 a_n100_n8267# VSUBS 0.216482f
C2664 a_100_n7134# VSUBS 0.190616f
C2665 a_n158_n7134# VSUBS 0.190616f
C2666 a_n100_n7231# VSUBS 0.216482f
C2667 a_100_n6098# VSUBS 0.190616f
C2668 a_n158_n6098# VSUBS 0.190616f
C2669 a_n100_n6195# VSUBS 0.216482f
C2670 a_100_n5062# VSUBS 0.190616f
C2671 a_n158_n5062# VSUBS 0.190616f
C2672 a_n100_n5159# VSUBS 0.216482f
C2673 a_100_n4026# VSUBS 0.190616f
C2674 a_n158_n4026# VSUBS 0.190616f
C2675 a_n100_n4123# VSUBS 0.216482f
C2676 a_100_n2990# VSUBS 0.190616f
C2677 a_n158_n2990# VSUBS 0.190616f
C2678 a_n100_n3087# VSUBS 0.216482f
C2679 a_100_n1954# VSUBS 0.190616f
C2680 a_n158_n1954# VSUBS 0.190616f
C2681 a_n100_n2051# VSUBS 0.216482f
C2682 a_100_n918# VSUBS 0.190616f
C2683 a_n158_n918# VSUBS 0.190616f
C2684 a_n100_n1015# VSUBS 0.216482f
C2685 a_100_118# VSUBS 0.190616f
C2686 a_n158_118# VSUBS 0.190616f
C2687 a_n100_21# VSUBS 0.216482f
C2688 a_100_1154# VSUBS 0.190616f
C2689 a_n158_1154# VSUBS 0.190616f
C2690 a_n100_1057# VSUBS 0.216482f
C2691 a_100_2190# VSUBS 0.190616f
C2692 a_n158_2190# VSUBS 0.190616f
C2693 a_n100_2093# VSUBS 0.216482f
C2694 a_100_3226# VSUBS 0.190616f
C2695 a_n158_3226# VSUBS 0.190616f
C2696 a_n100_3129# VSUBS 0.216482f
C2697 a_100_4262# VSUBS 0.190616f
C2698 a_n158_4262# VSUBS 0.190616f
C2699 a_n100_4165# VSUBS 0.216482f
C2700 a_100_5298# VSUBS 0.190616f
C2701 a_n158_5298# VSUBS 0.190616f
C2702 a_n100_5201# VSUBS 0.216482f
C2703 a_100_6334# VSUBS 0.190616f
C2704 a_n158_6334# VSUBS 0.190616f
C2705 a_n100_6237# VSUBS 0.216482f
C2706 a_100_7370# VSUBS 0.190616f
C2707 a_n158_7370# VSUBS 0.190616f
C2708 a_n100_7273# VSUBS 0.216482f
C2709 a_100_8406# VSUBS 0.190616f
C2710 a_n158_8406# VSUBS 0.190616f
C2711 a_n100_8309# VSUBS 0.216482f
C2712 a_100_9442# VSUBS 0.190616f
C2713 a_n158_9442# VSUBS 0.190616f
C2714 a_n100_9345# VSUBS 0.216482f
C2715 a_100_10478# VSUBS 0.190616f
C2716 a_n158_10478# VSUBS 0.190616f
C2717 a_n100_10381# VSUBS 0.216482f
C2718 a_100_11514# VSUBS 0.190616f
C2719 a_n158_11514# VSUBS 0.190616f
C2720 a_n100_11417# VSUBS 0.216482f
C2721 a_100_12550# VSUBS 0.190616f
C2722 a_n158_12550# VSUBS 0.190616f
C2723 a_n100_12453# VSUBS 0.216482f
C2724 a_100_13586# VSUBS 0.190616f
C2725 a_n158_13586# VSUBS 0.190616f
C2726 a_n100_13489# VSUBS 0.216482f
C2727 a_100_14622# VSUBS 0.190616f
C2728 a_n158_14622# VSUBS 0.190616f
C2729 a_n100_14525# VSUBS 0.216482f
C2730 a_100_15658# VSUBS 0.190616f
C2731 a_n158_15658# VSUBS 0.190616f
C2732 a_n100_15561# VSUBS 0.216482f
C2733 a_100_16694# VSUBS 0.190616f
C2734 a_n158_16694# VSUBS 0.190616f
C2735 a_n100_16597# VSUBS 0.216482f
C2736 a_100_17730# VSUBS 0.190616f
C2737 a_n158_17730# VSUBS 0.190616f
C2738 a_n100_17633# VSUBS 0.216482f
C2739 a_100_18766# VSUBS 0.190616f
C2740 a_n158_18766# VSUBS 0.190616f
C2741 a_n100_18669# VSUBS 0.216482f
C2742 a_100_19802# VSUBS 0.190616f
C2743 a_n158_19802# VSUBS 0.190616f
C2744 a_n100_19705# VSUBS 0.216482f
C2745 a_100_20838# VSUBS 0.190616f
C2746 a_n158_20838# VSUBS 0.190616f
C2747 a_n100_20741# VSUBS 0.216482f
C2748 a_100_21874# VSUBS 0.190616f
C2749 a_n158_21874# VSUBS 0.190616f
C2750 a_n100_21777# VSUBS 0.216482f
C2751 a_100_22910# VSUBS 0.190616f
C2752 a_n158_22910# VSUBS 0.190616f
C2753 a_n100_22813# VSUBS 0.216482f
C2754 a_100_23946# VSUBS 0.190616f
C2755 a_n158_23946# VSUBS 0.190616f
C2756 a_n100_23849# VSUBS 0.216482f
C2757 a_100_24982# VSUBS 0.190616f
C2758 a_n158_24982# VSUBS 0.190616f
C2759 a_n100_24885# VSUBS 0.216482f
C2760 a_100_26018# VSUBS 0.190616f
C2761 a_n158_26018# VSUBS 0.190616f
C2762 a_n100_25921# VSUBS 0.216482f
C2763 a_100_27054# VSUBS 0.190616f
C2764 a_n158_27054# VSUBS 0.190616f
C2765 a_n100_26957# VSUBS 0.216482f
C2766 a_100_28090# VSUBS 0.190616f
C2767 a_n158_28090# VSUBS 0.190616f
C2768 a_n100_27993# VSUBS 0.216482f
C2769 a_100_29126# VSUBS 0.190616f
C2770 a_n158_29126# VSUBS 0.190616f
C2771 a_n100_29029# VSUBS 0.216482f
C2772 a_100_30162# VSUBS 0.190616f
C2773 a_n158_30162# VSUBS 0.190616f
C2774 a_n100_30065# VSUBS 0.216482f
C2775 a_100_31198# VSUBS 0.190616f
C2776 a_n158_31198# VSUBS 0.190616f
C2777 a_n100_31101# VSUBS 0.216482f
C2778 a_100_32234# VSUBS 0.190616f
C2779 a_n158_32234# VSUBS 0.190616f
C2780 a_n100_32137# VSUBS 0.216482f
C2781 a_100_33270# VSUBS 0.190616f
C2782 a_n158_33270# VSUBS 0.190616f
C2783 a_n100_33173# VSUBS 0.216482f
C2784 a_100_34306# VSUBS 0.190616f
C2785 a_n158_34306# VSUBS 0.190616f
C2786 a_n100_34209# VSUBS 0.216482f
C2787 a_100_35342# VSUBS 0.190616f
C2788 a_n158_35342# VSUBS 0.190616f
C2789 a_n100_35245# VSUBS 0.216482f
C2790 a_100_36378# VSUBS 0.190616f
C2791 a_n158_36378# VSUBS 0.190616f
C2792 a_n100_36281# VSUBS 0.216482f
C2793 a_100_37414# VSUBS 0.190616f
C2794 a_n158_37414# VSUBS 0.190616f
C2795 a_n100_37317# VSUBS 0.216482f
C2796 a_100_38450# VSUBS 0.190616f
C2797 a_n158_38450# VSUBS 0.190616f
C2798 a_n100_38353# VSUBS 0.216482f
C2799 a_100_39486# VSUBS 0.190616f
C2800 a_n158_39486# VSUBS 0.190616f
C2801 a_n100_39389# VSUBS 0.216482f
C2802 a_100_40522# VSUBS 0.190616f
C2803 a_n158_40522# VSUBS 0.190616f
C2804 a_n100_40425# VSUBS 0.216482f
C2805 a_100_41558# VSUBS 0.190616f
C2806 a_n158_41558# VSUBS 0.190616f
C2807 a_n100_41461# VSUBS 0.216482f
C2808 a_100_42594# VSUBS 0.190616f
C2809 a_n158_42594# VSUBS 0.190616f
C2810 a_n100_42497# VSUBS 0.216482f
C2811 a_100_43630# VSUBS 0.190616f
C2812 a_n158_43630# VSUBS 0.190616f
C2813 a_n100_43533# VSUBS 0.216482f
C2814 a_100_44666# VSUBS 0.190616f
C2815 a_n158_44666# VSUBS 0.190616f
C2816 a_n100_44569# VSUBS 0.216482f
C2817 a_100_45702# VSUBS 0.190616f
C2818 a_n158_45702# VSUBS 0.190616f
C2819 a_n100_45605# VSUBS 0.216482f
C2820 a_100_46738# VSUBS 0.190616f
C2821 a_n158_46738# VSUBS 0.190616f
C2822 a_n100_46641# VSUBS 0.216482f
C2823 a_100_47774# VSUBS 0.190616f
C2824 a_n158_47774# VSUBS 0.190616f
C2825 a_n100_47677# VSUBS 0.216482f
C2826 a_100_48810# VSUBS 0.190616f
C2827 a_n158_48810# VSUBS 0.190616f
C2828 a_n100_48713# VSUBS 0.216482f
C2829 a_100_49846# VSUBS 0.190616f
C2830 a_n158_49846# VSUBS 0.190616f
C2831 a_n100_49749# VSUBS 0.216482f
C2832 a_100_50882# VSUBS 0.190616f
C2833 a_n158_50882# VSUBS 0.190616f
C2834 a_n100_50785# VSUBS 0.216482f
C2835 a_100_51918# VSUBS 0.190616f
C2836 a_n158_51918# VSUBS 0.190616f
C2837 a_n100_51821# VSUBS 0.216482f
C2838 a_100_52954# VSUBS 0.190616f
C2839 a_n158_52954# VSUBS 0.190616f
C2840 a_n100_52857# VSUBS 0.216482f
C2841 a_100_53990# VSUBS 0.190616f
C2842 a_n158_53990# VSUBS 0.190616f
C2843 a_n100_53893# VSUBS 0.216482f
C2844 a_100_55026# VSUBS 0.190616f
C2845 a_n158_55026# VSUBS 0.190616f
C2846 a_n100_54929# VSUBS 0.216482f
C2847 a_100_56062# VSUBS 0.190616f
C2848 a_n158_56062# VSUBS 0.190616f
C2849 a_n100_55965# VSUBS 0.216482f
C2850 a_100_57098# VSUBS 0.190616f
C2851 a_n158_57098# VSUBS 0.190616f
C2852 a_n100_57001# VSUBS 0.216482f
C2853 a_100_58134# VSUBS 0.190616f
C2854 a_n158_58134# VSUBS 0.190616f
C2855 a_n100_58037# VSUBS 0.216482f
C2856 a_100_59170# VSUBS 0.190616f
C2857 a_n158_59170# VSUBS 0.190616f
C2858 a_n100_59073# VSUBS 0.216482f
C2859 a_100_60206# VSUBS 0.190616f
C2860 a_n158_60206# VSUBS 0.190616f
C2861 a_n100_60109# VSUBS 0.216482f
C2862 a_100_61242# VSUBS 0.190616f
C2863 a_n158_61242# VSUBS 0.190616f
C2864 a_n100_61145# VSUBS 0.216482f
C2865 a_100_62278# VSUBS 0.190616f
C2866 a_n158_62278# VSUBS 0.190616f
C2867 a_n100_62181# VSUBS 0.216482f
C2868 a_100_63314# VSUBS 0.190616f
C2869 a_n158_63314# VSUBS 0.190616f
C2870 a_n100_63217# VSUBS 0.216482f
C2871 a_100_64350# VSUBS 0.190616f
C2872 a_n158_64350# VSUBS 0.190616f
C2873 a_n100_64253# VSUBS 0.216482f
C2874 a_100_65386# VSUBS 0.190616f
C2875 a_n158_65386# VSUBS 0.190616f
C2876 a_n100_65289# VSUBS 0.216482f
C2877 a_100_66422# VSUBS 0.190616f
C2878 a_n158_66422# VSUBS 0.190616f
C2879 a_n100_66325# VSUBS 0.216482f
C2880 a_100_67458# VSUBS 0.190616f
C2881 a_n158_67458# VSUBS 0.190616f
C2882 a_n100_67361# VSUBS 0.216482f
C2883 a_100_68494# VSUBS 0.190616f
C2884 a_n158_68494# VSUBS 0.190616f
C2885 a_n100_68397# VSUBS 0.216482f
C2886 a_100_69530# VSUBS 0.190616f
C2887 a_n158_69530# VSUBS 0.190616f
C2888 a_n100_69433# VSUBS 0.216482f
C2889 a_100_70566# VSUBS 0.190616f
C2890 a_n158_70566# VSUBS 0.190616f
C2891 a_n100_70469# VSUBS 0.216482f
C2892 a_100_71602# VSUBS 0.190616f
C2893 a_n158_71602# VSUBS 0.190616f
C2894 a_n100_71505# VSUBS 0.216482f
C2895 a_100_72638# VSUBS 0.190616f
C2896 a_n158_72638# VSUBS 0.190616f
C2897 a_n100_72541# VSUBS 0.216482f
C2898 a_100_73674# VSUBS 0.190616f
C2899 a_n158_73674# VSUBS 0.190616f
C2900 a_n100_73577# VSUBS 0.216482f
C2901 a_100_74710# VSUBS 0.190616f
C2902 a_n158_74710# VSUBS 0.190616f
C2903 a_n100_74613# VSUBS 0.216482f
C2904 a_100_75746# VSUBS 0.190616f
C2905 a_n158_75746# VSUBS 0.190616f
C2906 a_n100_75649# VSUBS 0.216482f
C2907 a_100_76782# VSUBS 0.190616f
C2908 a_n158_76782# VSUBS 0.190616f
C2909 a_n100_76685# VSUBS 0.216482f
C2910 a_100_77818# VSUBS 0.190616f
C2911 a_n158_77818# VSUBS 0.190616f
C2912 a_n100_77721# VSUBS 0.216482f
C2913 a_100_78854# VSUBS 0.190616f
C2914 a_n158_78854# VSUBS 0.190616f
C2915 a_n100_78757# VSUBS 0.216482f
C2916 a_100_79890# VSUBS 0.190616f
C2917 a_n158_79890# VSUBS 0.190616f
C2918 a_n100_79793# VSUBS 0.216482f
C2919 a_100_80926# VSUBS 0.190616f
C2920 a_n158_80926# VSUBS 0.190616f
C2921 a_n100_80829# VSUBS 0.216482f
C2922 a_100_81962# VSUBS 0.190616f
C2923 a_n158_81962# VSUBS 0.190616f
C2924 a_n100_81865# VSUBS 0.216482f
C2925 a_100_82998# VSUBS 0.190616f
C2926 a_n158_82998# VSUBS 0.190616f
C2927 a_n100_82901# VSUBS 0.216482f
C2928 a_100_84034# VSUBS 0.190616f
C2929 a_n158_84034# VSUBS 0.190616f
C2930 a_n100_83937# VSUBS 0.216482f
C2931 a_100_85070# VSUBS 0.190616f
C2932 a_n158_85070# VSUBS 0.190616f
C2933 a_n100_84973# VSUBS 0.216482f
C2934 a_100_86106# VSUBS 0.190616f
C2935 a_n158_86106# VSUBS 0.190616f
C2936 a_n100_86009# VSUBS 0.216482f
C2937 a_100_87142# VSUBS 0.190616f
C2938 a_n158_87142# VSUBS 0.190616f
C2939 a_n100_87045# VSUBS 0.216482f
C2940 a_100_88178# VSUBS 0.190616f
C2941 a_n158_88178# VSUBS 0.190616f
C2942 a_n100_88081# VSUBS 0.216482f
C2943 a_100_89214# VSUBS 0.190616f
C2944 a_n158_89214# VSUBS 0.190616f
C2945 a_n100_89117# VSUBS 0.216482f
C2946 a_100_90250# VSUBS 0.190616f
C2947 a_n158_90250# VSUBS 0.190616f
C2948 a_n100_90153# VSUBS 0.216482f
C2949 a_100_91286# VSUBS 0.190616f
C2950 a_n158_91286# VSUBS 0.190616f
C2951 a_n100_91189# VSUBS 0.216482f
C2952 a_100_92322# VSUBS 0.190616f
C2953 a_n158_92322# VSUBS 0.190616f
C2954 a_n100_92225# VSUBS 0.216482f
C2955 a_100_93358# VSUBS 0.190616f
C2956 a_n158_93358# VSUBS 0.190616f
C2957 a_n100_93261# VSUBS 0.216482f
C2958 a_100_94394# VSUBS 0.190616f
C2959 a_n158_94394# VSUBS 0.190616f
C2960 a_n100_94297# VSUBS 0.216482f
C2961 a_100_95430# VSUBS 0.190616f
C2962 a_n158_95430# VSUBS 0.190616f
C2963 a_n100_95333# VSUBS 0.216482f
C2964 a_100_96466# VSUBS 0.190616f
C2965 a_n158_96466# VSUBS 0.190616f
C2966 a_n100_96369# VSUBS 0.216482f
C2967 a_100_97502# VSUBS 0.190616f
C2968 a_n158_97502# VSUBS 0.190616f
C2969 a_n100_97405# VSUBS 0.216482f
C2970 a_100_98538# VSUBS 0.190616f
C2971 a_n158_98538# VSUBS 0.190616f
C2972 a_n100_98441# VSUBS 0.216482f
C2973 a_100_99574# VSUBS 0.190616f
C2974 a_n158_99574# VSUBS 0.190616f
C2975 a_n100_99477# VSUBS 0.216482f
C2976 a_100_100610# VSUBS 0.190616f
C2977 a_n158_100610# VSUBS 0.190616f
C2978 a_n100_100513# VSUBS 0.216482f
C2979 a_100_101646# VSUBS 0.190616f
C2980 a_n158_101646# VSUBS 0.190616f
C2981 a_n100_101549# VSUBS 0.216482f
C2982 a_100_102682# VSUBS 0.190616f
C2983 a_n158_102682# VSUBS 0.190616f
C2984 a_n100_102585# VSUBS 0.216482f
C2985 a_100_103718# VSUBS 0.190616f
C2986 a_n158_103718# VSUBS 0.190616f
C2987 a_n100_103621# VSUBS 0.216482f
C2988 a_100_104754# VSUBS 0.190616f
C2989 a_n158_104754# VSUBS 0.190616f
C2990 a_n100_104657# VSUBS 0.216482f
C2991 a_100_105790# VSUBS 0.190616f
C2992 a_n158_105790# VSUBS 0.190616f
C2993 a_n100_105693# VSUBS 0.216482f
C2994 a_100_106826# VSUBS 0.190616f
C2995 a_n158_106826# VSUBS 0.190616f
C2996 a_n100_106729# VSUBS 0.216482f
C2997 a_100_107862# VSUBS 0.190616f
C2998 a_n158_107862# VSUBS 0.190616f
C2999 a_n100_107765# VSUBS 0.216482f
C3000 a_100_108898# VSUBS 0.190616f
C3001 a_n158_108898# VSUBS 0.190616f
C3002 a_n100_108801# VSUBS 0.216482f
C3003 a_100_109934# VSUBS 0.190616f
C3004 a_n158_109934# VSUBS 0.190616f
C3005 a_n100_109837# VSUBS 0.216482f
C3006 a_100_110970# VSUBS 0.190616f
C3007 a_n158_110970# VSUBS 0.190616f
C3008 a_n100_110873# VSUBS 0.216482f
C3009 a_100_112006# VSUBS 0.190616f
C3010 a_n158_112006# VSUBS 0.190616f
C3011 a_n100_111909# VSUBS 0.216482f
C3012 a_100_113042# VSUBS 0.190616f
C3013 a_n158_113042# VSUBS 0.190616f
C3014 a_n100_112945# VSUBS 0.216482f
C3015 a_100_114078# VSUBS 0.190616f
C3016 a_n158_114078# VSUBS 0.190616f
C3017 a_n100_113981# VSUBS 0.216482f
C3018 a_100_115114# VSUBS 0.190616f
C3019 a_n158_115114# VSUBS 0.190616f
C3020 a_n100_115017# VSUBS 0.216482f
C3021 a_100_116150# VSUBS 0.190616f
C3022 a_n158_116150# VSUBS 0.190616f
C3023 a_n100_116053# VSUBS 0.216482f
C3024 a_100_117186# VSUBS 0.190616f
C3025 a_n158_117186# VSUBS 0.190616f
C3026 a_n100_117089# VSUBS 0.216482f
C3027 a_100_118222# VSUBS 0.190616f
C3028 a_n158_118222# VSUBS 0.190616f
C3029 a_n100_118125# VSUBS 0.216482f
C3030 a_100_119258# VSUBS 0.190616f
C3031 a_n158_119258# VSUBS 0.190616f
C3032 a_n100_119161# VSUBS 0.216482f
C3033 a_100_120294# VSUBS 0.190616f
C3034 a_n158_120294# VSUBS 0.190616f
C3035 a_n100_120197# VSUBS 0.216482f
C3036 a_100_121330# VSUBS 0.190616f
C3037 a_n158_121330# VSUBS 0.190616f
C3038 a_n100_121233# VSUBS 0.216482f
C3039 a_100_122366# VSUBS 0.190616f
C3040 a_n158_122366# VSUBS 0.190616f
C3041 a_n100_122269# VSUBS 0.216482f
C3042 a_100_123402# VSUBS 0.190616f
C3043 a_n158_123402# VSUBS 0.190616f
C3044 a_n100_123305# VSUBS 0.216482f
C3045 a_100_124438# VSUBS 0.190616f
C3046 a_n158_124438# VSUBS 0.190616f
C3047 a_n100_124341# VSUBS 0.216482f
C3048 a_100_125474# VSUBS 0.190616f
C3049 a_n158_125474# VSUBS 0.190616f
C3050 a_n100_125377# VSUBS 0.216482f
C3051 a_100_126510# VSUBS 0.190616f
C3052 a_n158_126510# VSUBS 0.190616f
C3053 a_n100_126413# VSUBS 0.216482f
C3054 a_100_127546# VSUBS 0.190616f
C3055 a_n158_127546# VSUBS 0.190616f
C3056 a_n100_127449# VSUBS 0.216482f
C3057 a_100_128582# VSUBS 0.190616f
C3058 a_n158_128582# VSUBS 0.190616f
C3059 a_n100_128485# VSUBS 0.216482f
C3060 a_100_129618# VSUBS 0.190616f
C3061 a_n158_129618# VSUBS 0.190616f
C3062 a_n100_129521# VSUBS 0.216482f
C3063 a_100_130654# VSUBS 0.190616f
C3064 a_n158_130654# VSUBS 0.190616f
C3065 a_n100_130557# VSUBS 0.216482f
C3066 a_100_131690# VSUBS 0.196066f
C3067 a_n158_131690# VSUBS 0.196066f
C3068 a_n100_131593# VSUBS 0.260213f
C3069 w_n358_n132787# VSUBS 0.711293p
.ends

.subckt pcell256scs avdd pbias pcbias sw_b sw_bn iout_n iout
XXM1 XM1/a_n158_n84606# XM1/a_n158_60430# XM1/a_n100_n31571# XM1/a_n100_n45931# XM1/a_n158_n111890#
+ XM1/a_n100_38793# XM1/a_n158_n15678# XM1/a_n158_n71682# XM1/a_n158_n136302# XM1/a_100_4426#
+ XM1/a_n100_76129# XM1/a_n100_n106243# XM1/a_n100_n14339# XM1/a_n158_n27166# XM1/a_n100_n70343#
+ XM1/a_n158_n83170# XM1/a_n158_158078# XM1/a_n100_n84703# XM1/a_n158_n97530# XM1/a_n100_n133527#
+ XM1/a_n158_17350# XM1/a_100_5862# XM1/a_100_123614# XM1/a_n158_n150662# XM1/a_n100_77565#
+ XM1/a_n100_123517# XM1/a_n158_30274# XM1/a_n158_44634# XM1/a_n100_n15775# XM1/a_n100_90489#
+ XM1/a_100_86278# XM1/a_n100_n134963# XM1/a_100_110690# XM1/a_n158_71918# XM1/a_n100_110593#
+ XM1/a_n158_n55886# XM1/a_n100_124953# XM1/a_n100_n145015# XM1/a_100_135102# XM1/a_n158_n106146#
+ XM1/a_n100_89053# XM1/a_n100_135005# XM1/a_n158_n176510# XM1/a_n158_n162150# XM1/a_n158_n1318#
+ XM1/a_n158_56122# XM1/a_n100_n27263# XM1/a_n100_n132091# XM1/a_n100_n146451# XM1/a_n158_n107582#
+ XM1/a_n100_122081# XM1/a_n100_n40187# XM1/a_n158_83406# XM1/a_n100_136441# XM1/a_n158_n2754#
+ XM1/a_n100_n54547# XM1/a_n158_n67374# XM1/a_n100_n68907# XM1/a_100_107818# XM1/a_100_n32910#
+ XM1/a_n100_n173735# XM1/a_100_163822# XM1/a_n158_n134866# XM1/a_n100_163725# XM1/a_n158_n80298#
+ XM1/a_n158_n94658# XM1/a_n158_14478# XM1/a_n158_28838# XM1/a_n158_70482# XM1/a_n158_84842#
+ XM1/a_n100_n55983# XM1/a_n158_n119070# XM1/a_n100_n66035# XM1/a_n100_n129219# XM1/a_100_119306#
+ XM1/a_n158_n146354# XM1/a_n100_119209# XM1/a_100_175310# XM1/a_100_n120506# XM1/a_n100_175213#
+ XM1/a_n100_n93319# XM1/a_n100_n67471# XM1/a_n158_96330# XM1/a_n100_n116295# XM1/a_n158_n173638#
+ XM1/a_100_106382# XM1/a_n100_106285# XM1/a_n158_n147790# XM1/a_n100_n80395# XM1/a_n100_n94755#
+ XM1/a_100_n121942# XM1/a_n100_n157939# XM1/a_n100_n143579# XM1/a_100_133666# XM1/a_n100_133569#
+ XM1/a_n100_147929# XM1/a_n158_54686# XM1/a_100_11606# XM1/a_100_n133430# XM1/a_100_n14242#
+ XM1/a_n100_n155067# XM1/a_100_n28602# XM1/a_n158_n116198# XM1/a_n100_n169427# XM1/a_100_145154#
+ XM1/a_100_159514# XM1/a_n100_145057# XM1/a_n100_159417# XM1/a_100_n160714# XM1/a_100_n41526#
+ XM1/a_n158_66174# XM1/a_100_172438# XM1/a_100_146590# XM1/a_n158_93458# XM1/a_n100_146493#
+ XM1/a_n100_n64599# XM1/a_n158_123614# XM1/a_n100_n78959# XM1/a_n100_n183787# XM1/a_100_n42962#
+ XM1/a_100_10170# XM1/a_100_24530# XM1/a_100_173874# XM1/a_100_n172202# XM1/a_n100_173777#
+ XM1/a_100_n53014# XM1/a_n158_94894# XM1/a_n158_110690# XM1/a_100_51814# XM1/a_n100_n76087#
+ XM1/a_100_n103274# XM1/a_n158_135102# XM1/a_100_n117634# XM1/a_100_n40090# XM1/a_100_129358#
+ XM1/a_100_n54450# XM1/a_100_n68810# XM1/a_100_n130558# XM1/a_100_n144918# XM1/a_n100_11509#
+ XM1/a_100_n81734# XM1/a_100_63302# XM1/a_100_n129122# XM1/a_n158_107818# XM1/a_n158_n32910#
+ XM1/a_100_n131994# XM1/a_n158_163822# XM1/a_n100_12945# XM1/a_100_n142046# XM1/a_100_n156406#
+ XM1/a_100_n37218# XM1/a_100_n93222# XM1/a_100_21658# XM1/a_n100_7201# XM1/a_n158_119306#
+ XM1/a_n158_n8498# XM1/a_n158_175310# XM1/a_100_n157842# XM1/a_100_n143482# XM1/a_100_n24294#
+ XM1/a_100_n38654# XM1/a_n100_n179479# XM1/a_n100_10073# XM1/a_n100_24433# XM1/a_100_169566#
+ XM1/a_n100_169469# XM1/a_100_n170766# XM1/a_100_n51578# XM1/a_n158_106382# XM1/a_100_n65938#
+ XM1/a_100_33146# XM1/a_n100_51717# XM1/a_100_47506# XM1/a_n158_4426# XM1/a_100_n169330#
+ XM1/a_n158_133666# XM1/a_n100_n4287# XM1/a_100_34582# XM1/a_100_48942# XM1/a_100_n182254#
+ XM1/a_n158_5862# XM1/a_100_n63066# XM1/a_100_n77426# XM1/a_n100_63205# XM1/a_100_61866#
+ XM1/a_n158_n14242# XM1/a_n158_145154# XM1/a_n158_n28602# XM1/a_100_n127686# XM1/a_n158_159514#
+ XM1/a_n100_n120603# XM1/a_100_n183690# XM1/a_100_n5626# XM1/a_n100_4329# XM1/a_n100_50281#
+ XM1/a_100_n78862# XM1/a_100_46070# XM1/a_n100_64641# XM1/a_n158_n41526# XM1/a_n158_172438#
+ XM1/a_n158_31710# XM1/a_100_n91786# XM1/a_n100_91925# XM1/a_n158_146590# XM1/a_100_73354#
+ XM1/a_100_87714# XM1/a_100_n139174# XM1/a_n100_5765# XM1/a_n158_n42962# XM1/a_n158_173874#
+ XM1/a_n100_22997# XM1/a_n158_n53014# XM1/a_100_18786# XM1/a_100_n166458# XM1/a_100_n152098#
+ XM1/a_100_74790# XM1/a_n100_33049# XM1/a_n158_n120506# XM1/a_n100_47409# XM1/a_100_n4190#
+ XM1/a_100_99202# XM1/a_n158_n40090# XM1/a_n100_n41623# XM1/a_n158_129358# XM1/a_n158_n54450#
+ XM1/a_n158_n68810# XM1/a_n100_n104807# XM1/a_100_n167894# XM1/a_n100_n160811# XM1/a_n100_34485#
+ XM1/a_n100_48845# XM1/a_n158_n121942# XM1/a_n100_150801# XM1/a_n158_n81734# XM1/a_n158_118#
+ XM1/a_n158_15914# XM1/a_n100_61769# XM1/a_100_43198# XM1/a_100_57558# XM1/a_n100_21#
+ XM1/a_n100_n53111# XM1/a_100_n179382# XM1/a_n158_n133430# XM1/a_n158_n37218# XM1/a_n158_n93222#
+ XM1/a_n158_13042# XM1/a_100_58994# XM1/a_100_1554# XM1/a_n158_27402# XM1/a_100_n87478#
+ XM1/a_n100_73257# XM1/a_n100_87617# XM1/a_n100_n103371# XM1/a_n158_n160714# XM1/a_100_69046#
+ XM1/a_n100_n117731# XM1/a_n100_n11467# XM1/a_n158_40326# XM1/a_n100_107721# XM1/a_n158_n24294#
+ XM1/a_n100_n25827# XM1/a_n158_n38654# XM1/a_n158_169566# XM1/a_n100_n81831# XM1/a_n100_n130655#
+ XM1/a_100_2990# XM1/a_n100_18689# XM1/a_100_120742# XM1/a_n100_74693# XM1/a_n100_120645#
+ XM1/a_n158_n51578# XM1/a_n158_n65938# XM1/a_n158_41762# XM1/a_n158_n172202# XM1/a_n100_99105#
+ XM1/a_100_97766# XM1/a_n100_n37315# XM1/a_n100_n142143# XM1/a_n158_n103274# XM1/a_n100_n156503#
+ XM1/a_100_132230# XM1/a_n100_n50239# XM1/a_n158_n117634# XM1/a_n100_86181# XM1/a_n100_132133#
+ XM1/a_n158_n63066# XM1/a_n158_n77426# XM1/a_n100_n24391# XM1/a_n158_53250# XM1/a_n158_67610#
+ XM1/a_n100_n38751# XM1/a_n158_n130558# XM1/a_n158_n144918# XM1/a_n158_80534# XM1/a_n100_n51675#
+ XM1/a_n158_n78862# XM1/a_n100_n100499# XM1/a_n100_n114859# XM1/a_n158_n129122# XM1/a_n100_n170863#
+ XM1/a_100_104946# XM1/a_n158_n131994# XM1/a_n100_58897# XM1/a_n100_104849# XM1/a_100_160950#
+ XM1/a_n100_160853# XM1/a_n158_n91786# XM1/a_n158_n142046# XM1/a_n158_25966# XM1/a_100_171002#
+ XM1/a_n158_n156406# XM1/a_n158_81970# XM4/w_n358_n132787# XM1/a_n158_36018# XM1/a_n100_n63163#
+ XM1/a_100_n104710# XM1/a_n158_92022# XM1/a_n100_n77523# XM1/a_n100_n126347# XM1/a_100_102074#
+ XM1/a_100_116434# XM1/a_n100_n182351# XM1/a_n100_116337# XM1/a_n158_n157842# XM1/a_n158_n143482#
+ XM1/a_n100_172341# XM1/a_n100_n90447# XM1/a_100_n12806# XM1/a_n158_23094# XM1/a_n158_37454#
+ XM1/a_100_143718# XM1/a_n158_n170766# XM1/a_100_79098# XM1/a_n100_97669# XM1/a_n100_n127783#
+ XM1/a_n158_50378# XM1/a_100_117870# XM1/a_n100_n35879# XM1/a_n100_n89011# XM1/a_n158_64738#
+ XM1/a_n100_117773# XM1/a_n100_n91883# XM1/a_n158_38890# XM1/a_100_130794# XM1/a_n158_n169330#
+ XM1/a_n100_130697# XM1/a_n100_n165119# XM1/a_100_155206# XM1/a_n100_155109# XM1/a_n158_n182254#
+ XM1/a_n100_n139271# XM1/a_n158_76226# XM1/a_n100_129261# XM1/a_n100_n47367# XM1/a_n158_n9934#
+ XM1/a_100_n11370# XM1/a_100_n25730# XM1/a_n100_n166555# XM1/a_n100_n152195# XM1/a_100_142282#
+ XM1/a_n158_n127686# XM1/a_n100_142185# XM1/a_100_156642# XM1/a_100_n101838# XM1/a_n158_n183690#
+ XM1/a_n100_156545# XM1/a_n158_n87478# XM1/a_100_20222# XM1/a_n158_77662# XM1/a_n100_n167991#
+ XM1/a_n158_n7062# XM1/a_n158_90586# XM1/a_n158_120742# XM1/a_n100_157981# XM1/a_n100_n178043#
+ XM1/a_100_114998# XM1/a_100_168130# XM1/a_100_n113326# XM1/a_n158_n139174# XM1/a_n100_168033#
+ XM1/a_n100_n5723# XM1/a_n100_n86139# XM1/a_100_7298# XM1/a_100_n50142# XM1/a_100_n64502#
+ XM1/a_n158_89150# XM1/a_100_181054# XM1/a_n158_n166458# XM1/a_n158_n152098# XM1/a_n158_132230#
+ XM1/a_n100_n87575# XM1/a_100_n114762# XM1/a_n100_n136399# XM1/a_100_126486# XM1/a_n100_126389#
+ XM1/a_100_182490# XM1/a_n158_n167894# XM1/a_n100_182393# XM1/a_100_n22858# XM1/a_100_60430#
+ XM1/a_100_n126250# XM1/a_n158_104946# XM1/a_n100_n99063# XM1/a_n158_160950# XM1/a_n158_n179382#
+ XM1/a_n158_171002# XM1/a_100_n153534# XM1/a_100_n34346# XM1/a_n100_20125# XM1/a_100_n48706#
+ XM1/a_100_n90350# XM1/a_100_165258# XM1/a_100_179618# XM1/a_100_n180818# XM1/a_n158_102074#
+ XM1/a_n158_86278# XM1/a_n158_116434# XM1/a_100_n154970# XM1/a_100_n35782# XM1/a_100_n109018#
+ XM1/a_n100_21561# XM1/a_n100_35921# XM1/a_100_166694# XM1/a_n158_n12806# XM1/a_100_n165022#
+ XM1/a_100_17350# XM1/a_n158_143718# XM1/a_n100_166597# XM1/a_n158_117870# XM1/a_100_30274#
+ XM1/a_100_44634# XM1/a_n158_1554# XM1/a_100_n73118# XM1/a_n158_130794# XM1/a_100_n47270#
+ XM1/a_100_71918# XM1/a_100_178182# XM1/a_100_n123378# XM1/a_100_n137738# XM1/a_n158_155206#
+ XM1/a_n100_178085# XM1/a_100_n1318# XM1/a_100_n60194# XM1/a_n158_2990# XM1/a_100_n74554#
+ XM1/a_100_n88914# XM1/a_n100_60333# XM1/a_100_56122# XM1/a_n158_n11370# XM1/a_n100_n12903#
+ XM1/a_n158_n25730# XM1/a_n158_142282# XM1/a_n158_156642# XM1/a_100_83406# XM1/a_100_n2754#
+ XM1/a_100_n19986# XM1/a_100_n75990# XM1/a_n100_1457# XM1/a_100_n149226# XM1/a_100_n86042#
+ XM1/a_100_14478# XM1/a_100_28838# XM1/a_100_70482# XM1/a_100_84842# XM1/a_n100_n10031#
+ XM1/a_n100_2893# XM1/a_n158_114998# XM1/a_n158_168130# XM1/a_n100_17253# XM1/a_n158_n104710#
+ XM1/a_n158_n50142# XM1/a_n158_n64502# XM1/a_100_n163586# XM1/a_n158_181054# XM1/a_100_n177946#
+ XM1/a_100_n44398# XM1/a_100_n58758# XM1/a_n100_30177# XM1/a_n100_44537# XM1/a_100_96330#
+ XM1/a_n158_11606# XM1/a_n158_126486# XM1/a_n158_182490# XM1/a_n100_n101935# XM1/a_n100_45973#
+ XM1/a_n158_n22858# XM1/a_100_n175074# XM1/a_n100_56025# XM1/a_100_54686# XM1/a_n100_83309#
+ XM1/a_n100_n113423# XM1/a_100_103510# XM1/a_n100_57461# XM1/a_n100_103413# XM1/a_n100_n21519#
+ XM1/a_n158_n34346# XM1/a_n158_n48706# XM1/a_n158_165258# XM1/a_n158_n90350# XM1/a_n158_179618#
+ XM1/a_n100_n140707# XM1/a_n158_10170# XM1/a_n158_24530# XM1/a_n158_n101838# XM1/a_n100_70385#
+ XM1/a_100_n98966# XM1/a_100_66174# XM1/a_n100_84745# XM1/a_n100_n22955# XM1/a_n158_51814#
+ XM1/a_n158_n35782# XM1/a_n158_166694# XM1/a_100_93458# XM1/a_n100_n33007# XM1/a_100_n159278#
+ XM1/a_100_n96094# XM1/a_n158_n113326# XM1/a_n100_96233# XM1/a_n158_n73118# XM1/a_100_94894#
+ XM1/a_n100_n20083# XM1/a_n158_63302# XM1/a_n100_n34443# XM1/a_n158_n47270# XM1/a_n100_n48803#
+ XM1/a_n158_178182# XM1/a_n100_n153631# XM1/a_n158_n114762# XM1/a_n158_n60194# XM1/a_n100_n61727#
+ XM1/a_n158_n74554# XM1/a_n100_143621# XM1/a_n158_n88914# XM1/a_100_100638# XM1/a_n100_n180915#
+ XM1/a_n100_54589# XM1/a_n100_68949# XM1/a_n100_170905# XM1/a_n158_7298# XM1/a_n158_21658#
+ XM1/a_n158_n19986# XM1/a_n100_n109115# XM1/a_n158_n75990# XM1/a_n100_n111987# XM1/a_n158_n126250#
+ XM1/a_100_n100402# XM1/a_n100_101977# XM1/a_n100_n73215# XM1/a_n158_n86042# XM1/a_n100_n122039#
+ XM1/a_100_8734# XM1/a_100_112126# XM1/a_n100_66077# XM1/a_n100_112029# XM1/a_n158_n153534#
+ XM1/a_n158_33146# XM1/a_n100_n18647# XM1/a_n158_47506# XM1/a_n100_n60291# XM1/a_n100_n74651#
+ XM1/a_n100_n123475# XM1/a_n158_n180818# XM1/a_100_113562# XM1/a_100_n8498# XM1/a_n100_n137835#
+ XM1/a_100_127922# XM1/a_n158_n44398# XM1/a_n100_113465# XM1/a_n100_127825# XM1/a_n158_n58758#
+ XM1/a_n158_n154970# XM1/a_n158_n109018# XM1/a_n158_n165022# XM1/a_n100_n150759#
+ XM1/a_n158_34582# XM1/a_n158_48942# XM1/a_100_140846# XM1/a_n100_94797# XM1/a_n100_140749#
+ XM1/a_n158_61866# XM1/a_n100_n149323# XM1/a_100_125050# XM1/a_100_139410# XM1/a_n100_n43059#
+ XM1/a_n100_n57419# XM1/a_n100_139313# XM1/a_n158_n5626# XM1/a_100_n140610# XM1/a_100_n21422#
+ XM1/a_n100_n162247# XM1/a_n158_46070# XM1/a_100_152334# XM1/a_n158_n123378# XM1/a_n158_n137738#
+ XM1/a_n100_n176607# XM1/a_n100_152237# XM1/a_n100_n44495# XM1/a_n158_73354# XM1/a_n158_87714#
+ XM1/a_n158_103510# XM1/a_n100_n58855# XM1/a_n100_n107679# XM1/a_n100_n163683# XM1/a_100_153770#
+ XM1/a_n100_153673# XM1/a_n100_n71779# XM1/a_n158_n98966# XM1/a_n158_18786# XM1/a_n158_n149226#
+ XM1/a_n158_74790# XM1/a_n100_n1415# XM1/a_100_31710# XM1/a_n100_180957# XM1/a_n158_99202#
+ XM1/a_n158_n4190# XM1/a_n100_n119167# XM1/a_100_109254# XM1/a_n100_n175171# XM1/a_n100_109157#
+ XM1/a_n100_n2851# XM1/a_n100_n83267# XM1/a_n158_n96094# XM1/a_100_n110454# XM1/a_100_n124814#
+ XM1/a_n100_165161# XM1/a_n100_179521# XM1/a_n100_n97627# XM1/a_100_122178# XM1/a_100_136538#
+ XM1/a_100_n61630# XM1/a_n158_n163586# XM1/a_n158_n177946# XM1/a_n158_43198# XM1/a_n158_57558#
+ XM1/a_n100_n28699# XM1/a_100_n111890# XM1/a_n100_n147887# XM1/a_100_137974# XM1/a_n158_100638#
+ XM1/a_100_n136302# XM1/a_n100_137877# XM1/a_100_n17114# XM1/a_100_148026# XM1/a_100_150898#
+ XM1/a_n158_n175074# XM1/a_100_15914# XM1/a_n158_58994# XM1/a_100_n30038# XM1/a_n158_69046#
+ XM1/a_n100_n96191# XM1/a_n100_n159375# XM1/a_100_n18550# XM1/a_100_149462# XM1/a_n158_112126#
+ XM1/a_n100_149365# XM1/a_100_n150662# XM1/a_n100_n172299# XM1/a_100_n31474# XM1/a_100_n45834#
+ XM1/a_100_13042# XM1/a_n100_31613# XM1/a_100_162386# XM1/a_100_176746# XM1/a_100_27402#
+ XM1/a_n100_162289# XM1/a_n100_176649# XM1/a_n158_113562# XM1/a_100_40326# XM1/a_n158_97766#
+ XM1/a_n158_127922# XM1/a_100_n106146# XM1/a_100_118# XM1/a_100_n176510# XM1/a_100_n162150#
+ XM1/a_n158_140846# XM1/a_n100_43101# XM1/a_100_n57322# XM1/a_n158_n159278# XM1/a_100_41762#
+ XM1/a_100_n70246# XM1/a_100_n84606# XM1/a_100_n107582# XM1/a_n158_125050# XM1/a_n158_139410#
+ XM1/a_n158_n21422# XM1/a_n158_152334# XM1/a_100_n134866# XM1/a_100_n15678# XM1/a_n100_15817#
+ XM1/a_100_n71682# XM1/a_n100_71821# XM1/a_100_53250# XM1/a_100_67610# XM1/a_100_n119070#
+ XM1/a_100_80534# XM1/a_n158_153770# XM1/a_100_n146354# XM1/a_100_n27166# XM1/a_n158_n100402#
+ XM1/a_n100_27305# XM1/a_100_158078# XM1/a_100_n83170# XM1/a_100_n97530# XM1/a_100_25966#
+ XM1/a_100_n173638# XM1/a_100_81970# XM1/a_n100_40229# XM1/a_n158_79098# XM1/a_n158_109254#
+ XM1/a_100_36018# XM1/a_100_n147790# XM1/a_100_92022# XM1/a_n100_14381# XM1/a_n100_28741#
+ XM1/a_n158_122178# XM1/a_n158_n61630# XM1/a_n158_136538# XM1/a_n100_41665# XM1/a_n100_n7159#
+ XM1/a_100_n55886# XM1/a_100_23094# XM1/a_100_37454# XM1/a_n158_8734# XM1/a_100_50378#
+ XM1/a_n158_137974# XM1/a_100_64738# XM1/a_n158_n17114# XM1/a_100_n116198# XM1/a_n158_148026#
+ XM1/a_n100_n8595# XM1/a_100_38890# XM1/a_n158_150898# XM1/a_100_n67374# XM1/a_n100_53153#
+ XM1/a_n100_67513# XM1/a_n158_n30038# XM1/a_n158_n140610# XM1/a_n158_20222# XM1/a_n158_n18550#
+ XM1/a_100_n80298# XM1/a_n100_80437# XM1/a_100_n94658# XM1/a_100_76226# XM1/a_n158_149462#
+ XM1/a_n100_n110551# XM1/a_n100_n124911# XM1/a_100_n9934# XM1/a_n100_8637# XM1/a_n158_n31474#
+ XM1/a_n100_100541# XM1/a_n100_114901# XM1/a_n158_n45834# XM1/a_n158_162386# XM1/a_n158_176746#
+ XM1/a_n100_25869# XM1/a_n100_79001# XM1/a_n100_81873# XM1/a_100_77662# XM1/a_n100_n17211#
+ XM1/a_100_n7062# XM1/a_100_90586# VSUBS XM1/a_n100_n30135# XM1/a_n158_n57322# XM1/a_n100_37357#
+ XM1/a_n158_n110454# XM1/a_n158_n124814# XM1/a_n100_93361# XM1/a_n158_n70246# XM1/a_100_89150#
+ sky130_fd_pr__pfet_g5v0d10v5_BK8KVU
XXM2 XM2/a_n100_n42155# XM2/a_100_n252938# XM2/a_n158_26478# XM2/a_n100_n226675# XM2/a_n158_n268754#
+ XM2/a_n100_n181863# XM2/a_n100_n21067# XM2/a_n100_n205587# XM2/a_n158_n247666# XM2/a_n100_n160775#
+ XM2/a_n158_n5154# XM2/a_n100_n324207# XM2/a_100_n334654# XM2/a_n100_n308391# XM2/a_n100_10565#
+ XM2/a_n158_n226578# XM2/a_n158_n181766# XM2/a_100_n47330# XM2/a_n100_n303119# XM2/a_100_n107958#
+ XM2/a_100_n313566# XM2/a_n158_n78962# XM2/a_n158_n329382# XM2/a_n100_n242491# XM2/a_n158_n284570#
+ XM2/a_100_13298# XM2/a_n158_n160678# XM2/a_100_n26242# XM2/a_n100_n155503# XM2/a_100_n165950#
+ XM2/a_n158_n308294# XM2/a_n158_n57874# XM2/a_n158_n263482# XM2/a_n100_n134415# XM2/a_100_29114#
+ XM2/a_n158_n36786# XM2/a_100_n144862# XM2/a_n158_n242394# XM2/a_n100_n184499# XM2/a_n100_n113327#
+ XM2/a_n158_n15698# XM2/a_100_n123774# XM2/a_n158_n155406# XM2/a_n158_n139590# XM2/a_n100_n57971#
+ XM2/a_n100_n216131# XM2/a_n158_n258210# XM2/a_n158_n134318# XM2/a_n158_n73690# XM2/a_100_n102686#
+ XM2/a_100_n292478# XM2/a_n100_n36883# XM2/a_100_n221306# XM2/a_100_n205490# XM2/a_n158_n237122#
+ XM2/a_n100_n150231# XM2/a_n100_n179227# XM2/a_100_n189674# XM2/a_n158_n192310# XM2/a_n100_n7887#
+ XM2/a_n100_n15795# XM2/a_100_n118502# XM2/a_100_n324110# XM2/a_100_n200218# XM2/a_n158_n216034#
+ XM2/a_n100_29017# XM2/a_n100_n158139# XM2/a_n158_n171222# XM2/a_100_n168586# XM2/a_n100_7929#
+ XM2/a_n100_n318935# XM2/a_100_n303022# XM2/a_100_n287206# XM2/a_n158_n150134# XM2/a_100_n147498#
+ XM2/a_n158_n310930# XM2/a_n158_n47330# XM2/a_100_n266118# XM2/a_n100_n195043# XM2/a_n158_n26242#
+ XM2/a_n158_n318838# XM2/a_n158_2754# XM2/a_100_n7790# XM2/a_n100_n231947# XM2/a_100_n2518#
+ XM2/a_100_n113230# XM2/a_n100_n334751# XM2/a_n100_n210859# XM2/a_n158_n252938# XM2/a_n100_2657#
+ XM2/a_n100_n313663# XM2/a_n100_n297847# XM2/a_100_n52602# XM2/a_n100_n92239# XM2/a_100_n179130#
+ XM2/a_n158_n334654# XM2/a_n100_n276759# XM2/a_100_n31514# XM2/a_n158_n107958# XM2/a_100_n158042#
+ XM2/a_n158_n313566# XM2/a_100_n81598# XM2/a_100_n10426# XM2/a_100_18570# XM2/a_n100_n123871#
+ XM2/a_n158_n165950# XM2/a_100_n97414# XM2/a_n100_n102783# XM2/a_n158_n144862# XM2/a_n100_n337387#
+ XM2/a_n100_n292575# XM2/a_100_n76326# XM2/a_n100_n221403# XM2/a_n158_21206# XM2/a_100_n231850#
+ XM2/a_n100_n316299# XM2/a_n158_n123774# XM2/a_n100_n189771# XM2/a_n100_n271487#
+ XM2/a_100_n55238# XM2/a_n100_n200315# XM2/a_100_n210762# XM2/a_100_n239758# XM2/a_n158_n102686#
+ XM2/a_n100_n168683# XM2/a_100_n194946# XM2/a_n100_n250399# XM2/a_n158_n292478# XM2/a_100_5390#
+ XM2/a_n158_118# XM2/a_n158_n221306# XM2/a_n158_n205490# XM2/a_100_n297750# XM2/a_n100_n287303#
+ XM2/a_n100_18473# XM2/a_100_n173858# XM2/a_n100_n147595# XM2/a_n158_n189674# XM2/a_n100_21#
+ XM2/a_n158_n118502# XM2/a_n158_n324110# XM2/a_100_n92142# XM2/a_n158_n200218# XM2/a_n100_n266215#
+ XM2/a_100_n276662# XM2/a_n158_n168586# XM2/a_n100_n86967# XM2/a_n158_n52602# XM2/a_n158_n303022#
+ XM2/a_100_n71054# XM2/a_n100_n245127# XM2/a_n158_n287206# XM2/a_100_n255574# XM2/a_n158_n147498#
+ XM2/a_n100_n65879# XM2/a_n158_n31514# XM2/a_n100_n224039# XM2/a_n158_n266118# XM2/a_100_n234486#
+ XM2/a_n158_n81598# XM2/a_n158_n10426# XM2/a_100_n337290# XM2/a_100_n213398# XM2/a_n100_n282031#
+ XM2/a_100_n332018# XM2/a_n158_n97414# XM2/a_n158_n113230# XM2/a_n100_n31611# XM2/a_100_n271390#
+ XM2/a_n100_n81695# XM2/a_100_n229214# XM2/a_n158_15934# XM2/a_n158_n76326# XM2/a_100_n184402#
+ XM2/a_n100_n2615# XM2/a_n100_n10523# XM2/a_n100_n39519# XM2/a_100_n279298# XM2/a_100_n20970#
+ XM2/a_100_n49966# XM2/a_100_n208126# XM2/a_100_n163314# XM2/a_n158_n55238# XM2/a_n100_n137051#
+ XM2/a_n158_n179130# XM2/a_n100_n97511# XM2/a_100_n28878# XM2/a_100_n142226# XM2/a_100_23842#
+ XM2/a_n158_n158042# XM2/a_n100_n76423# XM2/a_100_n86870# XM2/a_100_n245030# XM2/a_100_n121138#
+ XM2/a_n158_n92142# XM2/a_n100_n55335# XM2/a_n158_10662# XM2/a_100_n65782# XM2/a_n100_n239855#
+ XM2/a_n158_n71054# XM2/a_n100_n34247# XM2/a_100_n44694# XM2/a_n100_n218767# XM2/a_n158_n231850#
+ XM2/a_n100_n173955# XM2/a_100_n187038# XM2/a_n100_n13159# XM2/a_n158_n210762# XM2/a_n158_n239758#
+ XM2/a_n100_23745# XM2/a_n100_n152867# XM2/a_n158_n194946# XM2/a_n100_n71151# XM2/a_100_n326746#
+ XM2/a_100_n281934# XM2/a_n158_n297750# XM2/a_n100_n255671# XM2/a_100_26478# XM2/a_n100_n131779#
+ XM2/a_n158_n173858# XM4/w_n358_n132787# XM2/a_n100_n50063# XM2/a_n100_n79059# XM2/a_100_n39422#
+ XM2/a_100_n305658# XM2/a_n158_5390# XM2/a_100_n260846# XM2/a_n100_n234583# XM2/a_n158_n276662#
+ XM2/a_100_n18334# XM2/a_100_n5154# XM2/a_n158_n20970# XM2/a_n158_n49966# XM2/a_n158_13298#
+ XM2/a_n100_n213495# XM2/a_n158_n255574# XM2/a_n100_n197679# XM2/a_n100_n126507#
+ XM2/a_n100_n332115# XM2/a_n158_n28878# XM2/a_100_n136954# XM2/a_n100_5293# XM2/a_n158_n234486#
+ XM2/a_n158_29114# XM2/a_n100_n229311# XM2/a_n100_n105419# XM2/a_n100_n311027# XM2/a_100_n115866#
+ XM2/a_100_n321474# XM2/a_n158_n86870# XM2/a_n158_n213398# XM2/a_n158_n337290# XM2/a_n100_n279395#
+ XM2/a_100_n34150# XM2/a_n100_n208223# XM2/a_n100_n163411# XM2/a_100_n218670# XM2/a_n158_n332018#
+ XM2/a_100_n300386# XM2/a_n158_n65782# XM2/a_n100_n28975# XM2/a_n158_n271390# XM2/a_100_n13062#
+ XM2/a_n158_n229214# XM2/a_n100_13201# XM2/a_n100_n142323# XM2/a_n158_n44694# XM2/a_100_n152770#
+ XM2/a_n158_n184402# XM2/a_100_8026# XM2/a_n158_n279298# XM2/a_100_n316202# XM2/a_n158_n208126#
+ XM2/a_n100_n121235# XM2/a_n158_n163314# XM2/a_100_n131682# XM2/a_100_n250302# XM2/a_n100_n100147#
+ XM2/a_100_n110594# XM2/a_n158_n142226# XM2/a_n100_n60607# XM2/a_n100_n44791# XM2/a_n158_n39422#
+ XM2/a_n158_n245030# XM2/a_n158_n121138# XM2/a_n100_n187135# XM2/a_100_n197582# XM2/a_n158_n18334#
+ XM2/a_100_n126410# XM2/a_n100_n166047# XM2/a_100_n176494# XM2/a_n158_n7790# XM2/a_100_n105322#
+ XM2/a_n100_n326843# XM2/a_100_n295114# XM2/a_n158_n187038# XM2/a_n158_n2518# XM2/a_n100_n305755#
+ XM2/a_100_n274026# XM2/a_n100_n260943# XM2/a_n100_n18431# XM2/a_n100_n289939# XM2/a_n158_n34150#
+ XM2/a_n158_n326746# XM2/a_100_n94778# XM2/a_n158_n281934# XM2/a_100_n23606# XM2/a_n158_n13062#
+ XM2/a_n158_n305658# XM2/a_n158_n260846# XM2/a_100_n100050# XM2/a_n100_n115963# XM2/a_100_n129046#
+ XM2/a_n100_n321571# XM2/a_100_n60510# XM2/a_100_n89506# XM2/a_n158_18570# XM2/a_n100_n300483#
+ XM2/a_n158_n136954# XM2/a_n100_n329479# XM2/a_n100_n284667# XM2/a_n100_n5251# XM2/a_100_n68418#
+ XM2/a_100_n223942# XM2/a_n158_n115866# XM2/a_n158_n321474# XM2/a_n100_n263579# XM2/a_100_n202854#
+ XM2/a_n158_n218670# XM2/a_n158_n300386# XM2/a_100_n289842# XM2/a_100_21206# XM2/a_n100_n110691#
+ XM2/a_n100_n139687# XM2/a_n158_n152770# XM2/a_n158_n316202# XM2/a_100_n84234# XM2/a_100_n268754#
+ XM2/a_n100_n258307# XM2/a_n100_n118599# XM2/a_n158_n131682# XM2/a_n158_8026# XM2/a_100_n63146#
+ XM2/a_n100_n237219# XM2/a_n158_n250302# XM2/a_100_n247666# XM2/a_n100_n192407# XM2/a_n158_n94778#
+ XM2/a_n158_n110594# XM2/a_n100_n176591# XM2/a_n158_n23606# XM2/a_100_n42058# XM2/a_100_n226578#
+ XM2/a_n100_n295211# XM2/a_n100_26381# XM2/a_n100_n171319# XM2/a_100_n181766# XM2/a_n158_n197582#
+ XM2/a_n158_n126410# XM2/a_100_n329382# XM2/a_n100_n274123# XM2/a_n100_21109# XM2/a_100_n284570#
+ XM2/a_100_n160678# XM2/a_100_118# XM2/a_n158_n176494# XM2/a_n100_n94875# XM2/a_n158_n60510#
+ XM2/a_n158_n89506# XM2/a_n158_n105322# XM2/a_100_n308294# XM2/a_n100_n253035# XM2/a_n158_n295114#
+ XM2/a_n100_n23703# XM2/a_100_n263482# XM2/a_n100_n73787# XM2/a_n158_n68418# XM2/a_n158_n274026#
+ XM2/a_100_n242394# XM2/a_n100_n52699# XM2/a_100_n155406# XM2/a_n100_n129143# XM2/a_100_n139590#
+ XM2/a_n100_n89603# XM2/a_100_n258210# XM2/a_100_n134318# XM2/a_100_15934# XM2/a_n100_n108055#
+ XM2/a_n100_n68515# XM2/a_n158_23842# XM2/a_100_n78962# XM2/a_100_n237122# XM2/a_100_n192310#
+ XM2/a_n158_n84234# XM2/a_n158_n100050# XM2/a_n158_n129046# XM2/a_n100_n47427# XM2/a_100_n57874#
+ XM2/a_n100_n202951# XM2/a_100_n216034# XM2/a_100_n171222# XM2/a_n158_n63146# XM2/a_n100_n26339#
+ XM2/a_100_n36786# XM2/a_n158_n223942# XM2/a_n158_n42058# XM2/a_100_n150134# XM2/a_100_2754#
+ XM2/a_n100_n84331# XM2/a_100_n310930# XM2/a_100_n15698# XM2/a_n158_n202854# XM2/a_n100_n268851#
+ XM2/a_100_10662# XM2/a_n100_15837# XM2/a_n100_n144959# XM2/a_n100_n63243# VSUBS
+ XM2/a_100_n318838# XM2/a_100_n73690# XM2/a_n100_n247763# XM2/a_n158_n289842# sky130_fd_pr__pfet_g5v0d10v5_AJ8KYZ
XXM3 m1_1634_n2388# m1_1634_n2388# XM3/a_n100_74613# m1_1634_n2388# XM3/a_n158_21874#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n63175# XM3/a_n100_n19663# XM3/a_n158_86106#
+ m1_1634_n2388# XM3/a_n158_n45466# XM3/a_n100_4165# XM3/a_n100_113981# m1_1634_n2388#
+ XM3/a_n100_n24843# XM3/a_n100_11417# XM3/a_n158_n50646# XM3/a_n158_82998# XM3/a_n100_n109795#
+ XM3/a_n158_n116950# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n114975# XM3/a_n100_95333#
+ XM3/a_n158_42594# XM3/a_n158_n10242# XM3/a_n100_n85967# m1_1634_n2388# m1_1634_n2388#
+ XM3/a_n100_115017# XM3/a_n158_n66186# m1_1634_n2388# XM3/a_n100_n45563# XM3/a_n100_32137#
+ XM3/a_n158_n27854# XM3/a_n158_n71366# XM3/a_n158_7370# m1_1634_n2388# XM3/a_n158_n109698#
+ XM3/a_n100_n50743# m1_1634_n2388# XM3/a_n158_105790# m1_1634_n2388# XM3/a_n158_n114878#
+ m1_1634_n2388# XM3/a_n158_110970# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_49749#
+ m1_1634_n2388# XM3/a_n158_n88978# XM3/a_n100_77721# XM3/a_n158_24982# XM3/a_n100_54929#
+ m1_1634_n2388# XM3/a_n100_82901# m1_1634_n2388# XM3/a_n100_n66283# XM3/a_n100_n100471#
+ XM3/a_n100_7273# XM3/a_n158_89214# XM3/a_n158_n48574# XM3/a_n158_n92086# XM3/a_n158_n1954#
+ m1_1634_n2388# XM3/a_n100_n27951# XM3/a_n100_n71463# XM3/a_n100_14525# XM3/a_n158_5298#
+ m1_1634_n2388# XM3/a_n158_112006# XM3/a_n158_n53754# m1_1634_n2388# m1_1634_n2388#
+ XM3/a_n158_131690# m1_1634_n2388# XM3/a_n158_26018# XM3/a_n100_98441# XM3/a_n158_n13350#
+ m1_1634_n2388# XM3/a_n100_75649# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_118125#
+ XM3/a_n158_129618# XM3/a_n158_50882# XM3/a_n100_n121191# XM3/a_n158_n100374# XM3/a_n100_80829#
+ m1_1634_n2388# XM3/a_n158_n69294# m1_1634_n2388# XM3/a_n100_n92183# XM3/a_n100_123305#
+ XM3/a_n100_n48671# XM3/a_n100_35245# XM3/a_n100_n25879# XM3/a_n158_n74474# m1_1634_n2388#
+ XM3/a_n100_n53851# XM3/a_n100_n119119# XM3/a_n100_40425# m1_1634_n2388# XM3/a_n158_n117986#
+ m1_1634_n2388# XM3/a_n158_n34070# m1_1634_n2388# XM3/a_n100_96369# XM3/a_n158_n11278#
+ m1_1634_n2388# XM3/a_n100_n1015# m1_1634_n2388# XM3/a_n158_n121094# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n100_n69391# XM3/a_n158_n95194# XM3/a_n100_n46599# XM3/a_n100_n74571#
+ XM3/a_n100_61145# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_17633# XM3/a_n158_97502#
+ XM3/a_n158_n56862# m1_1634_n2388# XM3/a_n158_115114# XM3/a_n100_n51779# m1_1634_n2388#
+ XM3/a_n100_22813# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_29126# m1_1634_n2388#
+ XM3/a_n100_n11375# XM3/a_n158_34306# XM3/a_n100_78757# XM3/a_n158_53990# m1_1634_n2388#
+ XM3/a_n158_n103482# XM3/a_n100_83937# m1_1634_n2388# XM3/a_n100_126413# XM3/a_n100_n95291#
+ XM3/a_n100_38353# m1_1634_n2388# XM3/a_n158_n77582# XM3/a_n100_n28987# XM3/a_n100_n72499#
+ m1_1634_n2388# XM3/a_n100_43533# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_n82762#
+ XM3/a_n100_n127407# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n32095# m1_1634_n2388#
+ XM3/a_n158_55026# XM3/a_n100_99477# XM3/a_n158_n14386# m1_1634_n2388# XM3/a_n100_n4123#
+ XM3/a_n158_60206# m1_1634_n2388# XM3/a_n100_59073# m1_1634_n2388# XM3/a_n100_108801#
+ XM3/a_n100_64253# XM3/a_n158_n59970# m1_1634_n2388# XM3/a_n158_118222# XM3/a_n100_n54887#
+ XM3/a_n158_77818# XM4/w_n358_n132787# m1_1634_n2388# XM3/a_n100_25921# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n158_123402# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n14483#
+ XM3/a_n158_37414# XM3/a_n158_n40286# XM3/a_n158_n106590# XM3/a_n158_n9206# XM3/a_n100_129521#
+ m1_1634_n2388# XM3/a_n158_n111770# XM3/a_n100_106729# XM3/a_n100_18669# XM3/a_n100_90153#
+ XM3/a_n158_98538# XM3/a_n100_46641# XM3/a_n158_n57898# XM3/a_n100_111909# XM3/a_n100_n80787#
+ XM3/a_n158_n85870# XM3/a_n100_23849# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_51821#
+ XM3/a_n158_58134# XM3/a_n158_n17494# m1_1634_n2388# XM3/a_n100_n7231# XM3/a_n100_n40383#
+ XM3/a_n158_63314# XM3/a_n158_19802# XM3/a_n158_n22674# XM3/a_n158_2190# m1_1634_n2388#
+ XM3/a_n158_n132490# XM3/a_n100_127449# m1_1634_n2388# XM3/a_n100_39389# XM3/a_n100_67361#
+ XM3/a_n100_n57995# XM3/a_n100_44569# XM3/a_n100_72541# m1_1634_n2388# XM3/a_n158_n83798#
+ m1_1634_n2388# XM3/a_n158_126510# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_103718#
+ m1_1634_n2388# XM3/a_n100_n17591# XM3/a_n158_84034# XM3/a_n158_118# XM3/a_n100_2093#
+ XM3/a_n100_n5159# XM3/a_n158_n43394# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n22771#
+ XM3/a_n158_45702# XM3/a_n100_n116011# XM3/a_n100_21# XM3/a_n100_88081# m1_1634_n2388#
+ XM3/a_n100_n87003# m1_1634_n2388# XM3/a_n100_109837# XM3/a_n100_65289# XM3/a_n100_93261#
+ XM3/a_n158_119258# m1_1634_n2388# XM3/a_n100_n83895# XM3/a_n100_26957# XM3/a_n100_70469#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_124438# m1_1634_n2388#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n43491# XM3/a_n100_30065# XM3/a_n158_66422#
+ m1_1634_n2388# XM3/a_n100_n20699# XM3/a_n158_n25782# XM3/a_n158_71602# m1_1634_n2388#
+ XM3/a_n158_n30962# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_47677# XM3/a_n100_91189#
+ m1_1634_n2388# XM3/a_n158_8406# m1_1634_n2388# XM3/a_n100_52857# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n158_106826# XM3/a_n158_87142# m1_1634_n2388# XM3/a_n100_n8267#
+ m1_1634_n2388# XM3/a_n100_100513# XM3/a_n100_12453# XM3/a_n158_92322# m1_1634_n2388#
+ XM3/a_n158_48810# XM3/a_n158_n51682# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_68397#
+ XM3/a_n100_n67319# m1_1634_n2388# XM3/a_n100_n101507# XM3/a_n100_8309# XM3/a_n100_73577#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n100_116053# XM3/a_n158_127546# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n100_121233# XM3/a_n100_33173# m1_1634_n2388# XM3/a_n158_69530#
+ XM3/a_n158_n28890# XM3/a_n158_n119022# m1_1634_n2388# XM3/a_n158_46738# XM3/a_n100_n117047#
+ XM3/a_n158_74710# XM3/a_n158_n124202# XM3/a_n100_n88039# m1_1634_n2388# XM3/a_n158_51918#
+ XM3/a_n100_n122227# m1_1634_n2388# XM3/a_n100_94297# XM3/a_n100_n93219# XM3/a_n158_n98302#
+ XM3/a_n100_n49707# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_11514# XM3/a_n100_55965#
+ XM3/a_n158_109934# XM3/a_n158_n35106# m1_1634_n2388# XM3/a_n158_67458# XM3/a_n100_103621#
+ XM3/a_n158_n2990# XM3/a_n100_15561# XM3/a_n158_95430# m1_1634_n2388# XM3/a_n158_113042#
+ XM3/a_n158_n54790# XM3/a_n158_72638# XM3/a_n158_n31998# XM3/a_n100_20741# m1_1634_n2388#
+ XM3/a_n158_27054# m1_1634_n2388# XM3/a_n100_n104615# XM3/a_n158_32234# XM3/a_n100_76685#
+ XM3/a_n100_n75607# m1_1634_n2388# XM3/a_n100_119161# m1_1634_n2388# XM3/a_n100_81865#
+ XM3/a_n158_n4026# m1_1634_n2388# XM3/a_n158_88178# XM3/a_n100_124341# XM3/a_n100_36281#
+ m1_1634_n2388# XM3/a_n100_n35203# XM3/a_n100_101549# XM3/a_n100_13489# XM3/a_n158_93358#
+ XM3/a_n158_n61006# XM3/a_n100_41461# XM3/a_n158_49846# XM3/a_n158_n80690# XM3/a_n158_n127310#
+ m1_1634_n2388# XM3/a_n100_n125335# XM3/a_n158_n104518# m1_1634_n2388# XM3/a_n158_100610#
+ XM3/a_n100_n96327# m1_1634_n2388# XM3/a_n100_n130515# m1_1634_n2388# XM3/a_n100_n2051#
+ XM3/a_n158_n78618# m1_1634_n2388# XM3/a_n158_14622# XM3/a_n100_117089# m1_1634_n2388#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n100_122269# XM3/a_n158_n38214# XM3/a_n100_62181#
+ XM3/a_n100_n61103# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_116150# XM3/a_n158_75746#
+ XM3/a_n158_n125238# XM3/a_n158_121330# m1_1634_n2388# XM3/a_n158_80926# XM3/a_n158_n130418#
+ XM3/a_n100_n107723# m1_1634_n2388# XM3/a_n158_n99338# XM3/a_n158_35342# XM3/a_n100_79793#
+ XM3/a_n100_n78715# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n112903# XM3/a_n158_40522#
+ XM3/a_n100_84973# XM3/a_n158_n7134# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n38311#
+ XM3/a_n100_104657# XM3/a_n158_n64114# XM3/a_n100_16597# XM3/a_n158_96466# XM3/a_n100_n15519#
+ XM3/a_n158_114078# XM3/a_n100_21777# XM3/a_n100_n128443# m1_1634_n2388# XM3/a_n158_n107626#
+ XM3/a_n158_56062# XM3/a_n100_n99435# m1_1634_n2388# XM3/a_n100_86009# XM3/a_n158_n112806#
+ XM3/a_n158_61242# XM3/a_n158_17730# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n158_n86906# XM3/a_n158_22910# m1_1634_n2388# XM3/a_n100_n59031#
+ XM3/a_n100_125377# m1_1634_n2388# XM3/a_n100_n36239# m1_1634_n2388# XM3/a_n100_n64211#
+ XM3/a_n100_130557# XM3/a_n100_42497# XM3/a_n158_n46502# XM3/a_n158_n90014# XM3/a_n100_5201#
+ XM3/a_n158_78854# XM3/a_n100_n41419# XM3/a_n158_n128346# m1_1634_n2388# m1_1634_n2388#
+ XM3/a_n158_3226# m1_1634_n2388# XM3/a_n158_101646# m1_1634_n2388# XM3/a_n158_38450#
+ XM3/a_n100_n3087# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_15658# XM3/a_n158_43630#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_20838# m1_1634_n2388# XM3/a_n100_107765#
+ XM3/a_n100_n62139# XM3/a_n158_n67222# XM3/a_n158_99574# XM3/a_n100_n18627# XM3/a_n100_n90111#
+ XM3/a_n158_117186# m1_1634_n2388# XM3/a_n100_3129# XM3/a_n100_112945# XM3/a_n100_24885#
+ XM3/a_n100_n23807# XM3/a_n158_n72402# XM3/a_n158_122366# m1_1634_n2388# XM3/a_n158_59170#
+ XM3/a_n100_n108759# XM3/a_n100_89117# XM3/a_n158_n115914# XM3/a_n158_36378# XM3/a_n158_64350#
+ m1_1634_n2388# XM3/a_n100_n113939# XM3/a_n158_41558# m1_1634_n2388# XM3/a_n100_128485#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n39347# XM3/a_n100_n44527# XM3/a_n158_n49610#
+ XM3/a_n158_n93122# m1_1634_n2388# XM3/a_n158_n26818# XM3/a_n158_6334# m1_1634_n2388#
+ XM3/a_n100_n129479# XM3/a_n100_50785# m1_1634_n2388# XM3/a_n158_104754# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n158_57098# XM3/a_n158_85070# XM3/a_n100_n6195# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n158_62278# XM3/a_n100_10381# XM3/a_n158_18766# XM3/a_n158_90250#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n158_23946# m1_1634_n2388# XM3/a_n158_n101410#
+ XM3/a_n100_n65247# m1_1634_n2388# XM3/a_n158_n47538# XM3/a_n100_6237# XM3/a_n158_n75510#
+ XM3/a_n100_27993# XM3/a_n100_n26915# XM3/a_n100_n70427# m1_1634_n2388# XM3/a_n158_125474#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n158_n52718# m1_1634_n2388# XM3/a_n158_130654#
+ XM3/a_n158_39486# m1_1634_n2388# XM3/a_n100_n30023# m1_1634_n2388# XM3/a_n100_97405#
+ XM3/a_n158_44666# XM3/a_n158_n12314# m1_1634_n2388# XM3/a_n158_n122130# m1_1634_n2388#
+ XM3/a_n100_n120155# XM3/a_n100_29029# XM3/a_n158_n68258# XM3/a_n100_57001# m1_1634_n2388#
+ XM3/a_n158_n96230# XM3/a_n100_n47635# XM3/a_n100_n91147# XM3/a_n100_34209# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n158_n29926# XM3/a_n158_n73438# XM3/a_n158_9442# XM3/a_n100_53893#
+ XM3/a_n100_n52815# m1_1634_n2388# XM3/a_n158_107862# m1_1634_n2388# m1_1634_n2388#
+ XM3/a_n158_n33034# m1_1634_n2388# XM3/a_n158_65386# m1_1634_n2388# XM3/a_n100_n12411#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n158_70566# XM3/a_n158_n120058# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n100_n68355# m1_1634_n2388# XM3/a_n100_n102543# XM3/a_n100_9345#
+ XM3/a_n158_n94158# XM3/a_n158_30162# XM3/a_n100_n73535# XM3/a_n100_60109# m1_1634_n2388#
+ m1_1634_n2388# XM3/a_n158_128582# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_n55826#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n33131# XM3/a_n158_91286#
+ XM3/a_n158_n15422# XM3/a_n158_47774# XM3/a_n100_n10339# XM3/a_n100_n118083# XM3/a_n158_52954#
+ XM3/a_n158_n20602# XM3/a_n100_n89075# XM3/a_n100_n123263# XM3/a_n158_n102446# m1_1634_n2388#
+ XM3/a_n100_n94255# XM3/a_n100_37317# m1_1634_n2388# XM3/a_n158_n76546# XM3/a_n158_12550#
+ m1_1634_n2388# XM3/a_n100_n55923# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_n81726#
+ m1_1634_n2388# XM3/a_n100_120197# m1_1634_n2388# XM3/a_n100_n31059# XM3/a_n158_n36142#
+ m1_1634_n2388# XM3/a_n158_68494# m1_1634_n2388# XM3/a_n158_73674# XM3/a_n158_n41322#
+ XM3/a_n158_n123166# m1_1634_n2388# XM3/a_n158_28090# XM3/a_n158_n918# XM3/a_n100_58037#
+ XM3/a_n158_n97266# XM3/a_n100_n105651# XM3/a_n158_33270# m1_1634_n2388# m1_1634_n2388#
+ XM3/a_n100_n76643# XM3/a_n100_63217# m1_1634_n2388# XM3/a_n100_n110831# XM3/a_n100_19705#
+ XM3/a_n158_n58934# XM3/a_n158_10478# m1_1634_n2388# XM3/a_n158_108898# XM3/a_n158_n5062#
+ m1_1634_n2388# XM3/a_n100_n81823# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388#
+ XM3/a_n100_102585# XM3/a_n158_94394# XM3/a_n100_n13447# XM3/a_n158_n18530# XM3/a_n158_n62042#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n158_n23710# XM3/a_n100_n126371# XM3/a_n158_n105554#
+ XM3/a_n100_n97363# XM3/a_n100_n103579# XM3/a_n100_n131551# XM3/a_n158_n110734# XM3/a_n158_31198#
+ XM3/a_n158_n79654# m1_1634_n2388# XM3/a_n100_45605# m1_1634_n2388# XM3/a_n158_n84834#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n34167# XM3/a_n158_n39250# m1_1634_n2388#
+ XM3/a_n158_n16458# XM3/a_n158_n44430# XM3/a_n158_76782# XM3/a_n158_n126274# m1_1634_n2388#
+ XM3/a_n158_n21638# XM3/a_n158_1154# XM3/a_n100_n124299# XM3/a_n158_81962# XM3/a_n158_n131454#
+ m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n79751# XM3/a_n100_66325# XM3/a_n158_13586#
+ XM3/a_n100_n56959# XM3/a_n158_n8170# m1_1634_n2388# XM3/a_n100_n84931# XM3/a_n100_71505#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM3/a_n158_n37178# m1_1634_n2388# m1_1634_n2388#
+ XM3/a_n100_105693# XM3/a_n158_n65150# m1_1634_n2388# XM3/a_n100_n16555# XM3/a_n100_n60067#
+ m1_1634_n2388# XM3/a_n100_1057# XM3/a_n100_31101# XM3/a_n100_110873# XM3/a_n158_n42358#
+ m1_1634_n2388# XM3/a_n158_n70330# XM3/a_n100_n21735# m1_1634_n2388# m1_1634_n2388#
+ XM3/a_n158_n108662# XM3/a_n158_120294# XM3/a_n100_n106687# XM3/a_n100_87045# XM3/a_n158_n113842#
+ m1_1634_n2388# XM3/a_n100_n77679# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n111867#
+ XM3/a_n100_92225# XM3/a_n100_48713# XM3/a_n158_n87942# XM3/a_n158_n6098# XM3/a_n100_n82859#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n37275#
+ m1_1634_n2388# XM3/a_n100_131593# XM3/a_n158_n19566# XM3/a_n158_n63078# m1_1634_n2388#
+ XM3/a_n100_n42455# XM3/a_n158_n91050# XM3/a_n158_79890# XM3/a_n100_n9303# XM3/a_n158_n129382#
+ m1_1634_n2388# XM3/a_n158_4262# m1_1634_n2388# XM3/a_n158_n24746# XM3/a_n158_102682#
+ m1_1634_n2388# VSUBS m1_1634_n2388# m1_1634_n2388# XM3/a_n100_n98399# m1_1634_n2388#
+ XM3/a_n100_n132587# XM3/a_n100_69433# XM3/a_n158_16694# sky130_fd_pr__pfet_g5v0d10v5_GK83LR
XXM4 XM4/a_100_n4026# XM4/a_100_n74474# XM4/a_n100_74613# XM4/a_100_88178# m1_1634_n2388#
+ XM4/a_100_93358# XM4/a_100_49846# XM4/a_n100_n63175# XM4/a_n100_n19663# m1_1634_n2388#
+ XM4/a_100_n34070# m1_1634_n2388# XM4/a_n100_4165# XM4/a_n100_113981# XM4/a_100_n11278#
+ XM4/a_n100_n24843# XM4/a_n100_11417# m1_1634_n2388# m1_1634_n2388# XM4/a_n100_n109795#
+ m1_1634_n2388# XM4/a_100_14622# XM4/a_100_n95194# XM4/a_n100_n114975# XM4/a_n100_95333#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_n100_n85967# XM4/a_100_115114# XM4/a_100_n56862#
+ XM4/a_n100_115017# m1_1634_n2388# XM4/a_100_75746# XM4/a_n100_n45563# XM4/a_n100_32137#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_80926# m1_1634_n2388# XM4/a_n100_n50743#
+ XM4/a_100_n106590# m1_1634_n2388# XM4/a_100_35342# m1_1634_n2388# XM4/a_100_n111770#
+ m1_1634_n2388# XM4/a_100_40522# XM4/a_100_n7134# XM4/a_100_2190# XM4/a_n100_49749#
+ XM4/a_100_n77582# m1_1634_n2388# XM4/a_n100_77721# m1_1634_n2388# XM4/a_n100_54929#
+ XM4/a_100_n82762# XM4/a_n100_82901# XM4/a_100_96466# XM4/a_n100_n66283# XM4/a_n100_n100471#
+ XM4/a_n100_7273# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n14386#
+ XM4/a_n100_n27951# XM4/a_n100_n71463# XM4/a_n100_14525# m1_1634_n2388# XM4/a_100_56062#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_100_n132490# XM4/a_100_61242# m1_1634_n2388#
+ XM4/a_100_17730# m1_1634_n2388# XM4/a_n100_98441# m1_1634_n2388# XM4/a_100_22910#
+ XM4/a_n100_75649# XM4/a_100_n59970# XM4/a_100_118222# XM4/a_n100_118125# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_n100_n121191# m1_1634_n2388# XM4/a_n100_80829# XM4/a_100_123402#
+ m1_1634_n2388# XM4/a_100_78854# XM4/a_n100_n92183# XM4/a_n100_123305# XM4/a_n100_n48671#
+ XM4/a_n100_35245# XM4/a_n100_n25879# m1_1634_n2388# XM4/a_100_n40286# XM4/a_n100_n53851#
+ XM4/a_n100_n119119# XM4/a_n100_40425# XM4/a_100_38450# m1_1634_n2388# XM4/a_100_15658#
+ m1_1634_n2388# XM4/a_100_43630# XM4/a_n100_96369# m1_1634_n2388# XM4/a_100_20838#
+ XM4/a_n100_n1015# XM4/a_100_n57898# m1_1634_n2388# XM4/a_100_n85870# XM4/a_100_99574#
+ XM4/a_n100_n69391# m1_1634_n2388# XM4/a_n100_n46599# XM4/a_n100_n74571# XM4/a_n100_61145#
+ XM4/a_100_n17494# XM4/a_100_8406# XM4/a_n100_17633# m1_1634_n2388# m1_1634_n2388#
+ XM4/a_100_59170# m1_1634_n2388# XM4/a_n100_n51779# XM4/a_100_n22674# XM4/a_n100_22813#
+ XM4/a_100_36378# XM4/a_100_64350# m1_1634_n2388# XM4/a_100_41558# XM4/a_n100_n11375#
+ m1_1634_n2388# XM4/a_n100_78757# m1_1634_n2388# XM4/a_100_n83798# m1_1634_n2388#
+ XM4/a_n100_83937# XM4/a_100_126510# XM4/a_n100_126413# XM4/a_n100_n95291# XM4/a_n100_38353#
+ XM4/a_100_103718# m1_1634_n2388# XM4/a_n100_n28987# XM4/a_n100_n72499# XM4/a_100_n43394#
+ XM4/a_n100_43533# XM4/a_100_57098# XM4/a_100_85070# m1_1634_n2388# XM4/a_n100_n127407#
+ XM4/a_100_18766# XM4/a_100_62278# XM4/a_n100_n32095# XM4/a_100_90250# m1_1634_n2388#
+ XM4/a_n100_99477# m1_1634_n2388# XM4/a_100_23946# XM4/a_n100_n4123# m1_1634_n2388#
+ XM4/a_100_119258# XM4/a_n100_59073# XM4/a_100_124438# XM4/a_n100_108801# XM4/a_n100_64253#
+ m1_1634_n2388# XM4/a_100_n119022# m1_1634_n2388# XM4/a_n100_n54887# m1_1634_n2388#
+ XM4/w_n358_n132787# XM4/a_100_n25782# XM4/a_n100_25921# XM4/a_100_39486# XM4/a_100_n124202#
+ m1_1634_n2388# XM4/a_100_n30962# XM4/a_100_44666# XM4/a_n100_n14483# m1_1634_n2388#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_n100_129521# XM4/a_100_106826#
+ m1_1634_n2388# XM4/a_n100_106729# XM4/a_n100_18669# XM4/a_n100_90153# m1_1634_n2388#
+ XM4/a_n100_46641# m1_1634_n2388# XM4/a_n100_111909# XM4/a_n100_n80787# m1_1634_n2388#
+ XM4/a_n100_23849# XM4/a_100_n51682# XM4/a_100_65386# XM4/a_n100_51821# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_100_70566# XM4/a_n100_n7231# XM4/a_n100_n40383# m1_1634_n2388#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_127546# m1_1634_n2388# XM4/a_n100_127449#
+ XM4/a_100_30162# XM4/a_n100_39389# XM4/a_n100_67361# XM4/a_n100_n57995# XM4/a_n100_44569#
+ XM4/a_n100_72541# XM4/a_100_n28890# m1_1634_n2388# XM4/a_100_n127310# m1_1634_n2388#
+ XM4/a_100_47774# XM4/a_100_91286# m1_1634_n2388# XM4/a_100_n104518# XM4/a_n100_n17591#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_n100_2093# XM4/a_n100_n5159# m1_1634_n2388#
+ XM4/a_100_n98302# XM4/a_100_52954# XM4/a_n100_n22771# m1_1634_n2388# XM4/a_n100_n116011#
+ XM4/a_n100_21# XM4/a_n100_88081# XM4/a_100_109934# XM4/a_n100_n87003# XM4/a_100_12550#
+ XM4/a_n100_109837# XM4/a_n100_65289# XM4/a_n100_93261# m1_1634_n2388# XM4/a_100_n35106#
+ XM4/a_n100_n83895# XM4/a_n100_26957# XM4/a_n100_70469# XM4/a_100_113042# XM4/a_100_n54790#
+ XM4/a_100_n125238# XM4/a_100_68494# m1_1634_n2388# XM4/a_100_n31998# XM4/a_100_73674#
+ XM4/a_100_n130418# XM4/a_n100_n43491# XM4/a_n100_30065# m1_1634_n2388# XM4/a_100_28090#
+ XM4/a_n100_n20699# m1_1634_n2388# m1_1634_n2388# XM4/a_100_33270# m1_1634_n2388#
+ XM4/a_100_10478# XM4/a_100_n5062# XM4/a_n100_47677# XM4/a_n100_91189# XM4/a_100_n61006#
+ m1_1634_n2388# XM4/a_100_n80690# XM4/a_n100_52857# XM4/a_100_94394# XM4/a_100_n107626#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_100_100610# XM4/a_n100_n8267# XM4/a_100_n112806#
+ XM4/a_n100_100513# XM4/a_n100_12453# m1_1634_n2388# XM4/a_100_3226# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_100_n78618# XM4/a_100_31198# XM4/a_n100_68397# XM4/a_n100_n67319#
+ XM4/a_100_n38214# XM4/a_n100_n101507# XM4/a_n100_8309# XM4/a_n100_73577# XM4/a_100_116150#
+ XM4/a_100_n128346# XM4/a_n100_116053# m1_1634_n2388# XM4/a_100_76782# XM4/a_100_121330#
+ XM4/a_n100_121233# XM4/a_n100_33173# XM4/a_100_n99338# m1_1634_n2388# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_100_81962# m1_1634_n2388# XM4/a_n100_n117047# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_n100_n88039# XM4/a_100_13586# m1_1634_n2388# XM4/a_n100_n122227#
+ XM4/a_100_n8170# XM4/a_n100_94297# XM4/a_n100_n93219# m1_1634_n2388# XM4/a_n100_n49707#
+ XM4/a_100_n64114# XM4/a_100_114078# m1_1634_n2388# XM4/a_n100_55965# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_100_n115914# m1_1634_n2388# XM4/a_n100_103621# m1_1634_n2388#
+ XM4/a_n100_15561# m1_1634_n2388# XM4/a_100_6334# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_n100_20741# XM4/a_100_n86906# m1_1634_n2388# XM4/a_100_n6098#
+ XM4/a_n100_n104615# m1_1634_n2388# XM4/a_n100_76685# XM4/a_n100_n75607# XM4/a_100_n90014#
+ XM4/a_n100_119161# XM4/a_100_n46502# XM4/a_n100_81865# m1_1634_n2388# XM4/a_100_79890#
+ m1_1634_n2388# XM4/a_n100_124341# XM4/a_n100_36281# XM4/a_100_101646# XM4/a_n100_n35203#
+ XM4/a_n100_101549# XM4/a_n100_13489# m1_1634_n2388# m1_1634_n2388# XM4/a_n100_41461#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_16694# XM4/a_n100_n125335#
+ m1_1634_n2388# XM4/a_100_n101410# m1_1634_n2388# XM4/a_n100_n96327# XM4/a_100_n67222#
+ XM4/a_n100_n130515# XM4/a_100_21874# XM4/a_n100_n2051# m1_1634_n2388# XM4/a_100_117186#
+ m1_1634_n2388# XM4/a_n100_117089# XM4/a_100_n72402# XM4/a_100_86106# XM4/a_100_122366#
+ XM4/a_n100_122269# m1_1634_n2388# XM4/a_n100_62181# XM4/a_n100_n61103# XM4/a_100_9442#
+ XM4/a_100_82998# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n122130#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_n100_n107723# XM4/a_100_42594# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_n100_79793# XM4/a_n100_n78715# XM4/a_100_n49610# XM4/a_100_n93122#
+ XM4/a_n100_n112903# m1_1634_n2388# XM4/a_n100_84973# m1_1634_n2388# XM4/a_100_n26818#
+ XM4/a_100_104754# XM4/a_n100_n38311# XM4/a_n100_104657# m1_1634_n2388# XM4/a_n100_16597#
+ m1_1634_n2388# XM4/a_n100_n15519# m1_1634_n2388# XM4/a_n100_21777# XM4/a_n100_n128443#
+ XM4/a_100_n120058# m1_1634_n2388# m1_1634_n2388# XM4/a_n100_n99435# XM4/a_100_24982#
+ XM4/a_n100_86009# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n47538#
+ XM4/a_100_n75510# XM4/a_100_89214# XM4/a_100_125474# m1_1634_n2388# m1_1634_n2388#
+ XM4/a_100_n52718# XM4/a_n100_n59031# XM4/a_n100_125377# XM4/a_100_n1954# XM4/a_n100_n36239#
+ XM4/a_100_130654# XM4/a_n100_n64211# XM4/a_n100_130557# XM4/a_n100_42497# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_n100_5201# m1_1634_n2388# XM4/a_n100_n41419# m1_1634_n2388#
+ XM4/a_100_n12314# XM4/a_100_26018# m1_1634_n2388# XM4/a_100_n102446# m1_1634_n2388#
+ XM4/a_100_n68258# m1_1634_n2388# XM4/a_n100_n3087# XM4/a_100_50882# XM4/a_100_n96230#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_100_n29926# XM4/a_100_n73438# XM4/a_100_n918#
+ m1_1634_n2388# XM4/a_100_107862# XM4/a_n100_107765# XM4/a_n100_n62139# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_n100_n18627# XM4/a_n100_n90111# m1_1634_n2388# XM4/a_100_n33034#
+ XM4/a_n100_3129# XM4/a_n100_112945# XM4/a_n100_24885# XM4/a_n100_n23807# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_100_n123166# m1_1634_n2388# XM4/a_n100_n108759# XM4/a_n100_89117#
+ m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n94158# XM4/a_n100_n113939#
+ m1_1634_n2388# XM4/a_100_128582# XM4/a_n100_128485# XM4/a_100_n55826# XM4/a_100_97502#
+ XM4/a_n100_n39347# XM4/a_n100_n44527# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n15422#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_100_29126# XM4/a_n100_n129479# XM4/a_n100_50785#
+ XM4/a_100_n105554# m1_1634_n2388# XM4/a_100_n20602# XM4/a_100_34306# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_n100_n6195# XM4/a_100_n110734# XM4/a_100_53990# m1_1634_n2388#
+ XM4/a_n100_10381# m1_1634_n2388# m1_1634_n2388# XM4/a_100_1154# XM4/a_100_n76546#
+ m1_1634_n2388# XM4/a_100_n81726# m1_1634_n2388# XM4/a_n100_n65247# XM4/a_100_n36142#
+ m1_1634_n2388# XM4/a_n100_6237# m1_1634_n2388# XM4/a_n100_27993# XM4/a_n100_n26915#
+ XM4/a_n100_n70427# XM4/a_100_n126274# m1_1634_n2388# XM4/a_100_n41322# XM4/a_100_55026#
+ m1_1634_n2388# XM4/a_100_n131454# m1_1634_n2388# m1_1634_n2388# XM4/a_100_60206#
+ XM4/a_n100_n30023# XM4/a_100_n97266# XM4/a_n100_97405# m1_1634_n2388# m1_1634_n2388#
+ XM4/a_100_n58934# m1_1634_n2388# XM4/a_100_108898# XM4/a_n100_n120155# XM4/a_n100_29029#
+ m1_1634_n2388# XM4/a_n100_57001# XM4/a_100_77818# m1_1634_n2388# XM4/a_n100_n47635#
+ XM4/a_n100_n91147# XM4/a_n100_34209# XM4/a_100_n18530# XM4/a_100_n62042# m1_1634_n2388#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_n100_53893# XM4/a_n100_n52815# XM4/a_100_n108662#
+ m1_1634_n2388# XM4/a_100_n23710# XM4/a_100_37414# m1_1634_n2388# XM4/a_100_n113842#
+ m1_1634_n2388# XM4/a_100_n9206# XM4/a_n100_n12411# XM4/a_100_n79654# XM4/a_100_4262#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_100_n84834# XM4/a_100_98538# XM4/a_n100_n68355#
+ XM4/a_100_n39250# XM4/a_n100_n102543# XM4/a_n100_9345# m1_1634_n2388# m1_1634_n2388#
+ XM4/a_n100_n73535# XM4/a_n100_60109# XM4/a_100_n16458# XM4/a_100_n129382# m1_1634_n2388#
+ XM4/a_100_n44430# XM4/a_100_58134# m1_1634_n2388# XM4/a_100_n21638# XM4/a_100_63314#
+ XM4/a_100_19802# XM4/a_n100_n33131# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388#
+ XM4/a_n100_n10339# XM4/a_n100_n118083# m1_1634_n2388# m1_1634_n2388# XM4/a_n100_n89075#
+ XM4/a_n100_n123263# m1_1634_n2388# XM4/a_100_n37178# XM4/a_n100_n94255# XM4/a_n100_37317#
+ XM4/a_100_n65150# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n42358# XM4/a_n100_n55923#
+ XM4/a_100_n70330# XM4/a_100_84034# m1_1634_n2388# XM4/a_100_120294# XM4/a_n100_120197#
+ XM4/a_100_n116950# XM4/a_n100_n31059# m1_1634_n2388# XM4/a_100_45702# m1_1634_n2388#
+ XM4/a_100_7370# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n87942# m1_1634_n2388#
+ m1_1634_n2388# XM4/a_n100_58037# m1_1634_n2388# XM4/a_n100_n105651# m1_1634_n2388#
+ XM4/a_100_n19566# XM4/a_100_n63078# XM4/a_n100_n76643# XM4/a_n100_63217# XM4/a_100_n91050#
+ XM4/a_n100_n110831# XM4/a_n100_19705# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n109698#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_100_n24746# XM4/a_n100_n81823# XM4/a_100_118#
+ XM4/a_100_66422# XM4/a_100_102682# XM4/a_100_n114878# XM4/a_n100_102585# m1_1634_n2388#
+ XM4/a_n100_n13447# m1_1634_n2388# m1_1634_n2388# XM4/a_100_5298# XM4/a_100_71602#
+ m1_1634_n2388# XM4/a_n100_n126371# m1_1634_n2388# XM4/a_n100_n97363# XM4/a_n100_n103579#
+ XM4/a_n100_n131551# m1_1634_n2388# m1_1634_n2388# m1_1634_n2388# XM4/a_100_n45466#
+ XM4/a_n100_45605# XM4/a_100_87142# m1_1634_n2388# XM4/a_100_n50646# XM4/a_100_92322#
+ XM4/a_n100_n34167# m1_1634_n2388# XM4/a_100_48810# m1_1634_n2388# m1_1634_n2388#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_100_n10242# m1_1634_n2388# m1_1634_n2388# XM4/a_n100_n124299#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_100_n100374# XM4/a_100_n66186# XM4/a_n100_n79751#
+ XM4/a_n100_66325# m1_1634_n2388# XM4/a_n100_n56959# m1_1634_n2388# XM4/a_100_n71366#
+ XM4/a_n100_n84931# XM4/a_n100_71505# XM4/a_100_n27854# XM4/a_100_69530# XM4/a_100_105790#
+ m1_1634_n2388# XM4/a_100_n117986# XM4/a_100_46738# XM4/a_n100_105693# m1_1634_n2388#
+ XM4/a_100_74710# XM4/a_n100_n16555# XM4/a_n100_n60067# XM4/a_100_110970# XM4/a_n100_1057#
+ XM4/a_n100_31101# XM4/a_n100_110873# m1_1634_n2388# XM4/a_100_51918# m1_1634_n2388#
+ XM4/a_n100_n21735# XM4/a_100_n88978# XM4/a_100_n121094# m1_1634_n2388# m1_1634_n2388#
+ XM4/a_n100_n106687# XM4/a_n100_87045# m1_1634_n2388# XM4/a_100_11514# XM4/a_n100_n77679#
+ XM4/a_100_n48574# XM4/a_100_n92086# XM4/a_n100_n111867# XM4/a_n100_92225# XM4/a_n100_48713#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_n100_n82859# XM4/a_100_n53754# XM4/a_100_67458#
+ XM4/a_100_112006# XM4/a_100_n2990# XM4/a_100_95430# XM4/a_n100_n37275# XM4/a_100_131690#
+ XM4/a_n100_131593# m1_1634_n2388# m1_1634_n2388# XM4/a_100_72638# XM4/a_n100_n42455#
+ m1_1634_n2388# m1_1634_n2388# XM4/a_n100_n9303# m1_1634_n2388# XM4/a_100_n13350#
+ m1_1634_n2388# XM4/a_100_27054# m1_1634_n2388# m1_1634_n2388# XM4/a_100_129618#
+ VSUBS XM4/a_100_n103482# XM4/a_100_32234# XM4/a_n100_n98399# XM4/a_100_n69294# XM4/a_n100_n132587#
+ XM4/a_n100_69433# m1_1634_n2388# sky130_fd_pr__pfet_g5v0d10v5_GK83LR
C0 XM1/a_n100_24433# XM3/a_n158_76782# 2.85e-20
C1 XM1/a_100_n166458# XM4/w_n358_n132787# 0.054058f
C2 XM4/w_n358_n132787# XM4/a_n100_5201# -0.004445f
C3 XM1/a_100_n173638# XM2/a_100_n326746# 4.64e-21
C4 XM1/a_n100_n63163# XM2/a_n158_n218670# 0.005074f
C5 XM1/a_n100_n44495# m1_1634_n2388# 1.3e-19
C6 XM1/a_n158_n9934# XM2/a_n158_n163314# 4.64e-21
C7 XM1/a_100_114998# XM2/a_n158_n39422# 0.116862f
C8 XM4/w_n358_n132787# XM4/a_n100_116053# -0.004445f
C9 XM2/a_n100_n129143# XM3/a_n158_75746# 1.66e-19
C10 XM2/a_100_n242394# XM3/a_n100_n35203# 1.93e-19
C11 XM4/w_n358_n132787# XM3/a_n158_n63078# 0.032295f
C12 XM4/a_n100_n49707# m1_1634_n2388# 0.072015f
C13 XM2/a_n100_n10523# XM1/a_100_142282# 0.005074f
C14 XM1/a_n100_103413# XM2/a_n158_n49966# 0.005074f
C15 XM2/a_n100_n171319# XM3/a_n158_33270# 0.005074f
C16 XM2/a_n100_26381# XM1/a_100_179618# 0.005074f
C17 XM2/a_n100_n282031# XM3/a_n100_n75607# 0.004501f
C18 XM1/a_n100_n109115# XM2/a_n158_n263482# 0.010147f
C19 XM2/a_n100_n102783# m1_1634_n2388# 9.96e-19
C20 XM3/a_n100_81865# XM4/a_n100_81865# 0.009521f
C21 XM1/a_100_18786# XM3/a_n100_70469# 1.72e-19
C22 XM1/a_n158_5862# XM3/a_n100_57001# 2.02e-20
C23 XM1/a_100_n84606# XM2/a_n100_n237219# 0.005074f
C24 XM1/a_100_n47270# XM2/a_100_n200218# 4.64e-21
C25 XM3/a_n100_47677# m1_1634_n2388# 0.072015f
C26 XM1/a_n158_4426# XM3/a_n100_54929# 1.94e-20
C27 XM2/a_n100_n92239# XM4/a_100_115114# 1.08e-20
C28 XM1/a_n100_n176607# m1_1634_n2388# 9.78e-20
C29 XM4/w_n358_n132787# XM2/a_100_n168586# 0.10588f
C30 XM2/a_100_n287206# m1_1634_n2388# 0.017213f
C31 XM1/a_n100_n94755# XM2/a_n158_n250302# 0.005074f
C32 XM1/a_100_n25730# XM4/w_n358_n132787# 0.053508f
C33 XM1/a_n100_n119167# XM4/w_n358_n132787# 0.012918f
C34 XM1/a_100_n97530# XM3/a_n158_n46502# 0.001362f
C35 XM4/w_n358_n132787# XM3/a_n158_89214# 0.032295f
C36 XM1/a_100_n163586# XM2/a_n100_n316299# 0.005074f
C37 XM2/a_100_n274026# XM3/a_n158_n69294# 0.071295f
C38 XM2/a_100_n316202# XM3/a_n100_n110831# 0.010147f
C39 XM1/a_n100_163725# XM2/a_n158_10662# 0.005074f
C40 XM1/a_n100_96233# XM2/a_100_n57874# 1.45e-19
C41 XM4/w_n358_n132787# XM4/a_n100_76685# -0.004445f
C42 XM1/a_100_n111890# XM2/a_n158_n266118# 0.116862f
C43 XM3/a_n100_n30023# m1_1634_n2388# 0.072015f
C44 XM4/w_n358_n132787# XM3/a_n158_34306# 0.032295f
C45 XM1/a_n100_79001# XM2/a_100_n76326# 7.26e-20
C46 XM1/a_100_100638# XM2/a_n158_n52602# 0.08181f
C47 XM2/a_n158_n89506# XM3/a_n100_117089# 7.26e-20
C48 XM2/a_n100_n89603# XM3/a_n158_117186# 0.005074f
C49 XM4/w_n358_n132787# XM3/a_n158_n102446# 0.032295f
C50 XM4/a_n100_n89075# m1_1634_n2388# 0.072015f
C51 XM1/a_100_n91786# XM2/a_n158_n245030# 0.0822f
C52 XM2/a_n158_n226578# XM3/a_n100_n22771# 7.48e-22
C53 XM1/a_n158_n50142# XM3/a_n100_2093# 1.94e-20
C54 XM1/a_n100_170905# XM2/a_100_18570# 7.26e-20
C55 XM1/a_n158_n74554# XM3/a_n100_n22771# 1.94e-20
C56 XM2/a_n158_n310930# XM3/a_n158_n104518# 4.64e-21
C57 XM3/a_n158_5298# m1_1634_n2388# 6.1e-20
C58 XM1/a_100_n179382# m1_1634_n2388# 0.002487f
C59 XM2/a_100_n223942# XM3/a_n100_n17591# 0.005074f
C60 XM1/a_n158_n180818# XM2/a_n158_n334654# 9.28e-21
C61 XM2/a_100_n200218# XM3/a_n100_5201# 0.010147f
C62 XM1/a_100_n44398# XM2/a_100_n197582# 4.64e-21
C63 XM4/w_n358_n132787# XM2/a_n100_n108055# 0.025717f
C64 XM1/a_n100_n106243# XM4/w_n358_n132787# 0.013376f
C65 XM2/a_n100_n226675# m1_1634_n2388# 0.002312f
C66 XM4/a_100_110970# m1_1634_n2388# 6.1e-20
C67 XM1/a_100_n55886# XM2/a_100_n210762# 4.64e-21
C68 XM1/a_n100_2893# m1_1634_n2388# 1.3e-19
C69 XM2/a_100_n105322# XM3/a_n100_99477# 0.010128f
C70 XM4/w_n358_n132787# XM2/a_100_n292478# 0.103341f
C71 XM1/a_100_n28602# XM3/a_n100_21777# 2.85e-20
C72 XM4/w_n358_n132787# XM4/a_n100_37317# -0.004445f
C73 XM3/a_n158_72638# m1_1634_n2388# 6.1e-20
C74 XM1/a_100_n100402# XM3/a_n100_n48671# 2.85e-20
C75 XM1/a_n100_157981# XM2/a_n158_5390# 0.005074f
C76 XM3/a_n100_103621# m1_1634_n2388# 0.072015f
C77 XM3/a_n100_n69391# m1_1634_n2388# 0.072015f
C78 XM1/a_n100_n25827# m1_1634_n2388# 1.05e-19
C79 XM2/a_100_n147498# XM3/a_n100_57001# 0.005074f
C80 XM4/a_n100_n128443# m1_1634_n2388# 0.072015f
C81 XM1/a_n100_n111987# XM2/a_n158_n266118# 0.010147f
C82 XM3/a_n158_17730# m1_1634_n2388# 6.1e-20
C83 XM1/a_n100_11509# XM2/a_n158_n142226# 0.010147f
C84 XM3/a_n100_n16555# XM4/a_n100_n16555# 0.009521f
C85 XM1/a_n100_45973# XM3/a_n100_96369# 5.2e-20
C86 XM1/a_100_n84606# XM4/w_n358_n132787# 0.054609f
C87 XM1/a_n100_124953# XM2/a_n158_n28878# 0.010147f
C88 XM2/a_n100_n260943# XM4/a_100_n56862# 2.13e-20
C89 XM2/a_100_n189674# XM3/a_n100_14525# 0.005074f
C90 XM2/a_100_n297750# XM3/a_n100_n93219# 0.005074f
C91 XM1/a_100_120742# XM2/a_n158_n34150# 0.107904f
C92 XM1/a_n158_40326# XM3/a_n100_92225# 1.94e-20
C93 XM2/a_n100_n144959# XM3/a_n158_62278# 0.005074f
C94 XM1/a_100_n57322# XM3/a_n158_n6098# 0.003402f
C95 XM4/w_n358_n132787# XM4/a_n100_n34167# -0.004445f
C96 XM3/a_n158_n5062# m1_1634_n2388# 6.1e-20
C97 XM1/a_100_66174# XM2/a_n100_n89603# 0.005074f
C98 XM1/a_n100_n25827# XM2/a_n158_n179130# 0.005074f
C99 XM2/a_n100_n187135# XM3/a_n158_19802# 0.005074f
C100 XM4/w_n358_n132787# XM1/a_n100_140749# 0.012279f
C101 XM4/a_100_71602# m1_1634_n2388# 6.1e-20
C102 XM1/a_100_44634# XM2/a_n100_n110691# 0.005074f
C103 XM4/w_n358_n132787# XM1/a_n100_n155067# 0.013408f
C104 XM2/a_n100_n147595# XM4/a_100_57098# 2.56e-20
C105 XM1/a_n158_2990# XM2/a_n158_n150134# 4.64e-21
C106 XM1/a_100_n78862# XM3/a_n158_n27854# 0.005291f
C107 XM1/a_n158_n75990# XM3/a_n100_n24843# 2.83e-20
C108 XM2/a_n158_n334654# XM3/a_n100_n128443# 1.41e-19
C109 XM3/a_n100_n108759# m1_1634_n2388# 0.072015f
C110 XM1/a_n100_n113423# XM2/a_100_n268754# 7.26e-20
C111 XM4/w_n358_n132787# XM2/a_n100_n231947# 0.025653f
C112 XM1/a_n158_n25730# XM3/a_n158_24982# 1.14e-21
C113 XM3/a_n158_128582# m1_1634_n2388# 6.1e-20
C114 XM1/a_n100_n126347# m1_1634_n2388# 1.3e-19
C115 XM3/a_n100_n36239# XM4/a_n100_n36239# 0.009521f
C116 XM2/a_100_n134318# XM3/a_n100_71505# 0.010147f
C117 XM2/a_n100_n245127# XM3/a_n100_n40383# 0.001266f
C118 XM1/a_n158_n73118# XM2/a_n100_n226675# 7.26e-20
C119 XM1/a_100_n8498# XM4/w_n358_n132787# 0.048914f
C120 XM1/a_n158_117870# XM2/a_n158_n36786# 9.28e-21
C121 XM4/w_n358_n132787# XM3/a_n100_101549# 0.009093f
C122 XM1/a_n100_n143579# XM3/a_n158_n91050# 1.99e-20
C123 XM1/a_100_n98966# XM3/a_n100_n47635# 5.71e-20
C124 XM1/a_n100_153673# XM4/w_n358_n132787# 0.01231f
C125 XM4/w_n358_n132787# XM3/a_n100_n14483# 0.00903f
C126 XM1/a_n100_113465# XM2/a_n158_n42058# 0.005074f
C127 XM1/a_100_n173638# XM2/a_n158_n326746# 0.068958f
C128 XM2/a_100_n176494# XM3/a_n100_29029# 0.010147f
C129 XM3/a_n100_49749# XM4/a_n100_49749# 0.009521f
C130 XM2/a_n100_n329479# XM3/a_n158_n122130# 0.003292f
C131 XM1/a_n158_n9934# XM2/a_n100_n163411# 7.26e-20
C132 XM4/w_n358_n132787# XM4/a_n100_n73535# -0.004445f
C133 XM3/a_n158_n44430# m1_1634_n2388# 6.1e-20
C134 XM2/a_n158_n242394# XM3/a_n100_n35203# 9.72e-21
C135 XM1/a_100_51814# XM3/a_n100_103621# 2.85e-20
C136 XM4/a_100_32234# m1_1634_n2388# 6.1e-20
C137 XM1/a_100_20222# XM3/a_n100_71505# 5.71e-20
C138 XM1/a_100_n45834# XM4/w_n358_n132787# 0.048442f
C139 XM1/a_n100_n127783# XM3/a_n158_n75510# 2.85e-20
C140 XM1/a_100_n120506# XM3/a_n100_n68355# 2.85e-20
C141 XM2/a_100_n100050# m1_1634_n2388# 0.017459f
C142 XM4/w_n358_n132787# XM3/a_n100_82901# 0.009157f
C143 XM1/a_100_n47270# XM2/a_n158_n200218# 0.05338f
C144 XM1/a_n100_n110551# m1_1634_n2388# 9.96e-20
C145 XM4/w_n358_n132787# XM3/a_n100_n3087# 0.009186f
C146 XM4/w_n358_n132787# XM2/a_n158_n168586# 0.107093f
C147 XM3/a_n100_n55923# XM4/a_n100_n55923# 0.009521f
C148 XM4/w_n358_n132787# XM3/a_n100_27993# 0.008742f
C149 XM1/a_n100_n165119# XM3/a_n158_n113842# 6.68e-21
C150 XM2/a_n100_n21067# XM1/a_100_135102# 0.001535f
C151 XM4/a_n100_95333# m1_1634_n2388# 0.072015f
C152 XM2/a_100_n121138# XM3/a_n100_86009# 0.003994f
C153 XM2/a_n158_n274026# XM3/a_n158_n69294# 4.64e-21
C154 XM4/w_n358_n132787# XM3/a_n100_n53851# 0.009186f
C155 XM4/a_100_n39250# m1_1634_n2388# 6.1e-20
C156 XM1/a_n158_n68810# XM2/a_n158_n221306# 4.64e-21
C157 XM4/w_n358_n132787# XM3/a_n158_126510# 0.032295f
C158 XM2/a_n158_n316202# XM3/a_n100_n110831# 1.45e-19
C159 XM4/w_n358_n132787# XM4/a_n100_n112903# -0.004445f
C160 XM2/a_100_n163314# XM3/a_n100_43533# 0.005074f
C161 XM1/a_n100_79001# XM2/a_n158_n76326# 0.005074f
C162 XM3/a_n158_n83798# m1_1634_n2388# 6.1e-20
C163 XM3/a_n158_n918# m1_1634_n2388# 6.1e-20
C164 XM2/a_100_n86870# XM3/a_n158_117186# 0.005476f
C165 XM1/a_100_n91786# XM2/a_n100_n245127# 0.005074f
C166 XM2/a_n100_n226675# XM3/a_n100_n22771# 0.005067f
C167 XM2/a_100_n205490# XM3/a_n158_1154# 0.054158f
C168 XM2/a_n158_n52602# XM4/w_n358_n132787# 0.104815f
C169 XM1/a_n100_66077# XM4/w_n358_n132787# 0.01363f
C170 XM1/a_n100_n71779# XM3/a_n158_n19566# 6.07e-19
C171 XM2/a_n100_n311027# XM3/a_n158_n104518# 2.47e-19
C172 XM1/a_n100_n97627# m1_1634_n2388# 1.3e-19
C173 XM2/a_n158_n223942# XM3/a_n100_n17591# 7.26e-20
C174 XM3/a_n100_66325# m1_1634_n2388# 0.072015f
C175 XM1/a_n100_15817# XM2/a_100_n139590# 7.26e-20
C176 XM3/a_n100_n75607# XM4/a_n100_n75607# 0.009521f
C177 XM2/a_n158_n200218# XM3/a_n100_5201# 1.45e-19
C178 XM1/a_100_n44398# XM2/a_n158_n197582# 0.076358f
C179 XM1/a_100_125050# XM4/w_n358_n132787# 0.048442f
C180 XM4/w_n358_n132787# XM2/a_100_n105322# 0.104259f
C181 XM1/a_n100_n150759# XM2/a_100_n303022# 4.26e-20
C182 XM2/a_100_n223942# m1_1634_n2388# 0.017213f
C183 XM4/a_n100_55965# m1_1634_n2388# 0.072015f
C184 XM4/w_n358_n132787# XM3/a_n100_n93219# 0.008254f
C185 XM4/a_100_n78618# m1_1634_n2388# 6.1e-20
C186 XM1/a_100_n55886# XM2/a_n158_n210762# 0.109462f
C187 XM3/a_n100_11417# m1_1634_n2388# 0.072015f
C188 XM2/a_n158_n105322# XM3/a_n100_99477# 1.44e-19
C189 XM1/a_n100_n166555# XM4/w_n358_n132787# 0.013101f
C190 XM4/w_n358_n132787# XM2/a_n158_n292478# 0.103107f
C191 XM1/a_n100_90489# XM2/a_n158_n63146# 0.010147f
C192 XM1/a_n100_n61727# XM3/a_n100_n9303# 3.12e-19
C193 XM3/a_n158_n123166# m1_1634_n2388# 6.1e-20
C194 XM1/a_100_n183690# XM3/a_n100_n132587# 2.85e-20
C195 XM4/w_n358_n132787# XM3/a_n158_52954# 0.032295f
C196 XM2/a_n158_n147498# XM3/a_n100_57001# 7.26e-20
C197 XM1/a_100_n71682# XM2/a_100_n226578# 4.64e-21
C198 XM1/a_n100_53153# XM2/a_100_n102686# 7.26e-20
C199 XM1/a_100_n182254# XM3/a_n100_n130515# 2.85e-20
C200 XM1/a_100_n176510# XM3/a_n100_n124299# 2.85e-20
C201 XM2/a_n158_n189674# XM3/a_n100_14525# 7.26e-20
C202 XM1/a_n158_n21422# XM3/a_n100_30065# 2.26e-20
C203 XM1/a_n100_157981# XM4/w_n358_n132787# 0.012279f
C204 XM2/a_n158_n297750# XM3/a_n100_n93219# 7.26e-20
C205 XM4/w_n358_n132787# XM3/a_n158_n28890# 0.032295f
C206 XM4/a_n100_n15519# m1_1634_n2388# 0.072015f
C207 XM2/a_100_n142226# XM3/a_n158_62278# 0.049095f
C208 XM3/a_n100_n95291# XM4/a_n100_n95291# 0.009521f
C209 XM1/a_100_66174# XM2/a_100_n86870# 4.64e-21
C210 XM1/a_n100_35921# XM3/a_n100_87045# 1.49e-19
C211 XM2/a_100_n252938# XM3/a_n158_n46502# 0.07441f
C212 XM1/a_n100_38793# XM4/w_n358_n132787# 0.013346f
C213 XM2/a_n100_n258307# XM4/a_100_n51682# 2.56e-20
C214 XM4/a_n100_16597# m1_1634_n2388# 0.072015f
C215 XM2/a_100_n184402# XM3/a_n158_19802# 0.019886f
C216 XM1/a_n100_n8595# XM2/a_100_n163314# 7.26e-20
C217 XM1/a_100_2990# XM2/a_100_n152770# 4.64e-21
C218 XM1/a_100_58994# XM2/a_n158_n94778# 0.116862f
C219 XM4/w_n358_n132787# XM3/a_n100_n132587# 0.011431f
C220 XM4/a_100_n117986# m1_1634_n2388# 6.1e-20
C221 XM2/a_100_n295114# XM3/a_n100_n88039# 0.005074f
C222 XM1/a_100_44634# XM2/a_100_n107958# 4.64e-21
C223 XM2/a_n100_n163411# m1_1634_n2388# 0.002793f
C224 XM1/a_n158_2990# XM2/a_n100_n150231# 7.26e-20
C225 XM1/a_n100_n44495# XM3/a_n158_7370# 2.85e-20
C226 XM3/a_n100_17633# XM4/a_n100_17633# 0.009521f
C227 XM2/a_n100_n334751# XM3/a_n100_n128443# 7.77e-20
C228 XM1/a_n100_n113423# XM2/a_n158_n268754# 0.005074f
C229 XM4/w_n358_n132787# XM2/a_100_n229214# 0.103342f
C230 XM1/a_n100_120645# XM2/a_n158_n34150# 0.005074f
C231 XM3/a_n158_91286# m1_1634_n2388# 6.1e-20
C232 XM3/a_n100_128485# m1_1634_n2388# 0.072015f
C233 XM4/w_n358_n132787# XM4/a_n100_110873# -0.004445f
C234 XM1/a_n100_n40187# XM3/a_n100_11417# 0.002268f
C235 XM1/a_n100_116337# XM2/a_n158_n39422# 0.005074f
C236 XM1/a_n100_n157939# XM3/a_n158_n105554# 2.85e-20
C237 XM2/a_n158_n134318# XM3/a_n100_71505# 1.45e-19
C238 XM2/a_n100_n144959# XM4/a_100_62278# 2.56e-20
C239 XM3/a_n158_36378# m1_1634_n2388# 6.1e-20
C240 XM1/a_n158_n183690# XM4/w_n358_n132787# 9.95e-32
C241 XM1/a_n100_n150759# m1_1634_n2388# 6.58e-20
C242 XM4/w_n358_n132787# XM3/a_n158_n68258# 0.032295f
C243 XM4/a_n100_n54887# m1_1634_n2388# 0.072015f
C244 XM1/a_100_n34346# XM3/a_n100_17633# 0.00124f
C245 XM1/a_100_n173638# XM2/a_n100_n326843# 0.005074f
C246 XM2/a_n158_n176494# XM3/a_n100_29029# 1.45e-19
C247 XM1/a_n100_30177# XM3/a_n158_81962# 2.67e-20
C248 XM1/a_n158_20222# XM3/a_n100_72541# 1.62e-20
C249 XM2/a_100_n326746# XM3/a_n158_n122130# 0.06f
C250 XM1/a_n100_n63163# XM2/a_100_n216034# 7.26e-20
C251 XM2/a_100_n129046# XM3/a_n158_76782# 0.077916f
C252 XM2/a_n100_n332115# XM4/a_100_n127310# 2.42e-20
C253 XM1/a_n100_n120603# XM3/a_n100_n69391# 0.001725f
C254 XM3/a_n100_n114975# XM4/a_n100_n114975# 0.009521f
C255 XM2/a_n100_n242491# XM3/a_n100_n35203# 0.00445f
C256 XM1/a_n158_17350# XM3/a_n100_68397# 1.94e-20
C257 XM2/a_100_n171222# XM3/a_n158_34306# 0.077916f
C258 XM1/a_100_77662# XM4/w_n358_n132787# 0.048442f
C259 XM1/a_100_168130# XM4/w_n358_n132787# 0.049181f
C260 XM1/a_n100_160853# XM2/a_n158_8026# 0.005074f
C261 XM2/a_n158_n100050# m1_1634_n2388# 2.36e-21
C262 XM1/a_100_n47270# XM2/a_n100_n200315# 0.005074f
C263 XM1/a_n100_100541# XM2/a_100_n52602# 7.26e-20
C264 XM2/a_100_n234486# XM3/a_n158_n28890# 0.077916f
C265 XM4/w_n358_n132787# XM2/a_n100_n168683# 0.024478f
C266 XM1/a_n100_166597# XM2/a_n158_10662# 0.004433f
C267 XM4/w_n358_n132787# XM4/a_n100_71505# -0.004445f
C268 XM2/a_n100_n287303# m1_1634_n2388# 7.61e-19
C269 XM3/a_n100_n35203# m1_1634_n2388# 0.072015f
C270 XM1/a_n100_133569# XM4/w_n358_n132787# 0.012279f
C271 XM1/a_n158_n136302# XM3/a_n100_n85967# 1.38e-20
C272 XM2/a_100_n276662# XM3/a_n100_n70427# 0.008289f
C273 XM1/a_n100_n94755# XM2/a_100_n247666# 7.26e-20
C274 XM2/a_n158_n121138# XM3/a_n100_86009# 4.26e-20
C275 XM4/w_n358_n132787# XM3/a_n158_n107626# 0.032295f
C276 XM4/a_n100_n94255# m1_1634_n2388# 0.072015f
C277 XM2/a_n100_n274123# XM3/a_n158_n69294# 0.003215f
C278 XM1/a_n158_n68810# XM2/a_n100_n221403# 7.26e-20
C279 XM4/w_n358_n132787# XM3/a_n100_126413# 0.009026f
C280 XM2/a_n100_n68515# XM4/w_n358_n132787# 0.011915f
C281 XM1/a_n100_n68907# XM4/w_n358_n132787# 0.013471f
C282 XM1/a_n100_n90447# XM3/a_n158_n38214# 2.85e-20
C283 XM2/a_n158_n163314# XM3/a_n100_43533# 7.26e-20
C284 XM2/a_100_n115866# XM3/a_n158_91286# 0.004697f
C285 XM1/a_n100_n31571# XM3/a_n100_18669# 2.27e-19
C286 XM2/a_n158_n86870# XM3/a_n158_117186# 4.64e-21
C287 XM2/a_100_n86870# XM3/a_n100_117089# 0.005074f
C288 XM1/a_n100_25869# XM2/a_100_n129046# 7.26e-20
C289 XM2/a_n158_n205490# XM3/a_n158_1154# 4.64e-21
C290 XM1/a_100_93458# XM4/w_n358_n132787# 0.048442f
C291 XM2/a_100_n158042# XM3/a_n158_48810# 0.033906f
C292 XM4/a_100_105790# m1_1634_n2388# 6.1e-20
C293 XM1/a_n158_123614# XM2/a_n100_n31611# 7.26e-20
C294 XM1/a_n100_n183787# XM2/a_100_n337290# 7.26e-20
C295 XM2/a_100_23842# XM1/a_n100_176649# 7.26e-20
C296 XM1/a_n100_n139271# m1_1634_n2388# 8.36e-20
C297 XM1/a_n100_n74651# XM3/a_n158_n22674# 2.85e-20
C298 XM2/a_n100_n224039# XM3/a_n100_n17591# 0.002257f
C299 XM4/w_n358_n132787# XM4/a_n100_32137# -0.004445f
C300 XM1/a_n100_15817# XM2/a_n158_n139590# 0.005074f
C301 XM3/a_n100_n74571# m1_1634_n2388# 0.072015f
C302 XM1/a_100_n44398# XM2/a_n100_n197679# 0.005074f
C303 XM1/a_n100_68949# XM2/a_100_n86870# 7.26e-20
C304 XM4/w_n358_n132787# XM2/a_n158_n105322# 0.107093f
C305 XM1/a_n100_93361# XM2/a_n158_n60510# 0.010147f
C306 XM1/a_n100_n150759# XM2/a_n158_n303022# 0.004271f
C307 XM4/w_n358_n132787# XM3/a_n100_46641# 0.009085f
C308 XM1/a_100_n55886# XM2/a_n100_n210859# 0.003918f
C309 XM2/a_n100_n105419# XM3/a_n100_99477# 3.11e-20
C310 XM1/a_100_63302# XM4/w_n358_n132787# 0.054708f
C311 XM4/w_n358_n132787# XM2/a_n100_n292575# 0.026631f
C312 XM1/a_n100_123517# XM2/a_n158_n28878# 0.005074f
C313 XM1/a_n158_n86042# XM3/a_n100_n34167# 1.94e-20
C314 XM3/a_n158_104754# m1_1634_n2388# 6.1e-20
C315 avdd pcbias 0.002316f
C316 XM2/a_100_n216034# XM3/a_n158_n11278# 0.073632f
C317 XM1/a_n100_n14339# m1_1634_n2388# 1.02e-19
C318 XM4/a_100_n131454# m1_1634_n2388# 6.1e-20
C319 XM2/a_100_n258210# XM3/a_n100_n52815# 0.010147f
C320 XM1/a_n158_84842# XM2/a_n100_n71151# 7.26e-20
C321 XM4/w_n358_n132787# XM4/a_n100_n39347# -0.004445f
C322 XM3/a_n158_n10242# m1_1634_n2388# 6.1e-20
C323 XM1/a_n100_48845# XM3/a_n158_99574# 2.85e-20
C324 XM1/a_100_n71682# XM2/a_n158_n226578# 0.107515f
C325 XM1/a_n100_53153# XM2/a_n158_n102686# 0.005074f
C326 XM2/a_n100_n305755# XM4/a_n100_n99435# 1.15e-20
C327 XM1/a_n100_169469# XM2/a_100_15934# 9.65e-20
C328 XM2/a_n158_n5154# XM4/w_n358_n132787# 0.106043f
C329 XM4/a_100_66422# m1_1634_n2388# 6.1e-20
C330 XM3/a_n100_70469# XM4/a_n100_70469# 0.009521f
C331 XM1/a_n100_n137835# XM2/a_100_n292478# 1.21e-19
C332 XM2/a_n158_n142226# XM3/a_n158_62278# 4.64e-21
C333 XM1/a_n100_n67471# XM4/w_n358_n132787# 0.01363f
C334 XM1/a_n100_n64599# XM3/a_n158_n12314# 2.85e-20
C335 XM1/a_100_66174# XM2/a_n158_n86870# 0.062727f
C336 XM3/a_n100_n113939# m1_1634_n2388# 0.072015f
C337 XM2/a_n158_n252938# XM3/a_n158_n46502# 4.64e-21
C338 XM1/a_n158_86278# XM2/a_n158_n68418# 9.28e-21
C339 XM3/a_n100_84973# m1_1634_n2388# 0.072015f
C340 XM1/a_n158_n54450# XM3/a_n100_n3087# 3.89e-20
C341 XM1/a_n158_n47270# XM2/a_n158_n202854# 4.64e-21
C342 XM2/a_n158_n184402# XM3/a_n158_19802# 4.64e-21
C343 XM1/a_n100_n8595# XM2/a_n158_n163314# 0.005074f
C344 XM1/a_100_2990# XM2/a_n158_n152770# 0.023391f
C345 XM2/a_n158_n295114# XM3/a_n100_n88039# 7.26e-20
C346 XM1/a_100_44634# XM2/a_n158_n107958# 0.018717f
C347 XM2/a_100_n160678# m1_1634_n2388# 0.018414f
C348 XM3/a_n100_30065# m1_1634_n2388# 0.072014f
C349 XM1/a_n100_147929# XM4/w_n358_n132787# 0.012279f
C350 XM1/a_n100_n100499# XM3/a_n158_n48574# 2.85e-20
C351 XM1/a_100_n30038# XM4/w_n358_n132787# 0.048442f
C352 XM4/a_n100_129521# m1_1634_n2388# 0.072015f
C353 XM4/w_n358_n132787# XM2/a_n158_n229214# 0.105525f
C354 XM4/w_n358_n132787# XM3/a_n100_n19663# 0.009186f
C355 XM4/a_100_n5062# m1_1634_n2388# 6.1e-20
C356 XM1/a_100_79098# XM2/a_n100_n73787# 0.005074f
C357 XM1/a_100_64738# XM3/a_n100_115017# 2.23e-20
C358 XM4/w_n358_n132787# XM4/a_n100_n78715# -0.004445f
C359 XM3/a_n158_n49610# m1_1634_n2388# 6.1e-20
C360 XM4/w_n358_n132787# XM3/a_n158_71602# 0.032295f
C361 XM4/w_n358_n132787# XM3/a_n158_102682# 0.032295f
C362 XM4/a_100_27054# m1_1634_n2388# 6.1e-20
C363 XM2/a_100_n200218# XM3/a_n158_6334# 0.063116f
C364 XM4/w_n358_n132787# XM3/a_n158_16694# 0.032295f
C365 XM1/a_n100_56025# m1_1634_n2388# 9.68e-20
C366 XM2/a_n158_n326746# XM3/a_n158_n122130# 4.64e-21
C367 XM1/a_n158_n170766# XM3/a_n100_n120155# 1.94e-20
C368 XM1/a_n100_n63163# XM2/a_n158_n216034# 0.005074f
C369 XM1/a_n158_n78862# XM3/a_n100_n27951# 1.86e-20
C370 XM2/a_100_n105322# XM3/a_n158_100610# 0.077916f
C371 XM2/a_100_n239758# XM3/a_n100_n35203# 0.005074f
C372 XM3/a_n100_126413# XM4/a_n100_126413# 0.009521f
C373 XM2/a_100_n324110# XM3/a_n158_n116950# 0.003918f
C374 XM1/a_n100_n4287# XM4/w_n358_n132787# 0.01363f
C375 XM1/a_n100_53153# XM3/a_n158_103718# 2.85e-20
C376 XM2/a_n100_n329479# XM4/a_100_n122130# 1.19e-20
C377 XM1/a_n158_n2754# XM3/a_n100_47677# 1.94e-20
C378 XM2/a_n100_n100147# m1_1634_n2388# 0.00103f
C379 XM4/a_n100_90153# m1_1634_n2388# 0.072015f
C380 XM4/w_n358_n132787# XM3/a_n100_n59031# 0.009131f
C381 XM4/a_100_n44430# m1_1634_n2388# 6.1e-20
C382 XM4/w_n358_n132787# XM2/a_100_n165950# 0.103341f
C383 XM2/a_n100_n89603# XM4/a_100_115114# 2.56e-20
C384 XM1/a_100_107818# XM2/a_n100_n44791# 0.005074f
C385 XM4/w_n358_n132787# XM4/a_n100_n118083# -0.004445f
C386 XM3/a_n158_n88978# m1_1634_n2388# 6.1e-20
C387 XM2/a_100_n284570# m1_1634_n2388# 0.021401f
C388 XM2/a_n158_n276662# XM3/a_n100_n70427# 1.27e-19
C389 XM1/a_n100_n94755# XM2/a_n158_n247666# 0.005074f
C390 XM2/a_n100_n121235# XM3/a_n100_86009# 0.001461f
C391 XM1/a_n100_n1415# XM3/a_n158_50882# 2.85e-20
C392 XM3/a_n158_55026# m1_1634_n2388# 6.1e-20
C393 XM1/a_n158_27402# XM2/a_n158_n126410# 9.28e-21
C394 XM1/a_100_n109018# XM4/w_n358_n132787# 0.048442f
C395 XM1/a_n158_n101838# XM3/a_n100_n49707# 1.94e-20
C396 XM1/a_n100_142185# XM2/a_100_n13062# 7.26e-20
C397 XM2/a_n158_n115866# XM3/a_n158_91286# 4.64e-21
C398 XM2/a_n158_n86870# XM3/a_n100_117089# 7.26e-20
C399 XM2/a_n100_n86967# XM3/a_n158_117186# 0.005074f
C400 XM1/a_n100_25869# XM2/a_n158_n129046# 0.005074f
C401 XM2/a_n100_n271487# XM3/a_n158_n64114# 0.001183f
C402 XM2/a_n100_n205587# XM3/a_n158_1154# 0.005074f
C403 XM1/a_100_182490# XM4/w_n358_n132787# 0.053288f
C404 XM1/a_100_171002# XM2/a_n100_15837# 0.005074f
C405 XM1/a_100_n169330# XM2/a_n158_n324110# 0.116862f
C406 XM2/a_n158_n158042# XM3/a_n158_48810# 4.64e-21
C407 XM4/a_n100_50785# m1_1634_n2388# 0.072015f
C408 XM4/w_n358_n132787# XM3/a_n100_n98399# 0.009601f
C409 XM4/a_100_n83798# m1_1634_n2388# 6.1e-20
C410 XM1/a_100_n133430# XM2/a_n158_n287206# 0.116862f
C411 XM1/a_n100_n183787# XM2/a_n158_n337290# 0.005078f
C412 XM1/a_n158_n45834# XM3/a_n100_6237# 1.94e-20
C413 XM1/a_n158_n150662# XM3/a_n100_n98399# 1.18e-20
C414 XM1/a_n100_n142143# XM2/a_100_n297750# 7.26e-20
C415 XM1/a_100_n106146# XM3/a_n100_n54887# 5.71e-20
C416 XM1/a_n100_68949# XM2/a_n158_n86870# 0.005074f
C417 XM4/w_n358_n132787# XM2/a_n100_n105419# 0.025057f
C418 XM3/a_n158_n128346# m1_1634_n2388# 6.1e-20
C419 XM1/a_n100_n150759# XM2/a_n100_n303119# 0.001243f
C420 XM2/a_n100_n224039# m1_1634_n2388# 0.002744f
C421 XM2/a_100_n305658# XM3/a_n158_n99338# 0.077916f
C422 XM1/a_n158_132230# XM2/a_n100_n21067# 7.26e-20
C423 XM2/a_n100_n311027# XM4/a_100_n104518# 3.16e-21
C424 XM3/a_n100_109837# XM4/a_n100_109837# 0.009521f
C425 XM4/w_n358_n132787# XM2/a_100_n289842# 0.106289f
C426 XM2/a_n100_n21067# XM4/w_n358_n132787# 0.011815f
C427 XM1/a_100_n173638# XM3/a_n158_n122130# 0.003891f
C428 XM1/a_n100_n157939# m1_1634_n2388# 9.55e-20
C429 XM3/a_n100_38353# XM4/a_n100_38353# 0.009521f
C430 XM3/a_n100_104657# m1_1634_n2388# 0.072015f
C431 XM4/w_n358_n132787# XM3/a_n158_n34070# 0.032295f
C432 XM4/a_n100_n20699# m1_1634_n2388# 0.072015f
C433 XM2/a_n158_n216034# XM3/a_n158_n11278# 4.64e-21
C434 XM2/a_n100_n10523# XM1/a_n158_142282# 7.26e-20
C435 XM1/a_n100_n123475# XM3/a_n158_n71366# 2.85e-20
C436 XM1/a_n158_n106146# XM3/a_n100_n54887# 3.89e-20
C437 XM2/a_n158_n258210# XM3/a_n100_n52815# 1.45e-19
C438 XM1/a_n100_n78959# XM3/a_n158_n26818# 2.85e-20
C439 XM1/a_n100_n35879# XM3/a_n158_14622# 2.85e-20
C440 XM1/a_100_n71682# XM2/a_n100_n226675# 0.005055f
C441 XM1/a_n100_n123475# m1_1634_n2388# 1.3e-19
C442 XM2/a_n100_n197679# XM4/a_100_9442# 2.56e-20
C443 XM4/a_n100_11417# m1_1634_n2388# 0.072015f
C444 XM1/a_n158_11606# XM2/a_n158_n142226# 9.28e-21
C445 XM4/a_100_n123166# m1_1634_n2388# 6.1e-20
C446 XM1/a_n100_n137835# XM2/a_n158_n292478# 0.007586f
C447 XM2/a_n100_n142323# XM3/a_n158_62278# 0.005074f
C448 XM1/a_100_n63066# XM3/a_n158_n11278# 0.001549f
C449 XM1/a_100_66174# XM2/a_n100_n86967# 0.005074f
C450 XM2/a_n100_n253035# XM3/a_n158_n46502# 7.31e-19
C451 XM1/a_n100_n156503# XM3/a_n158_n104518# 2.85e-20
C452 XM1/a_n158_n47270# XM2/a_n100_n202951# 7.26e-20
C453 XM2/a_n100_n184499# XM3/a_n158_19802# 0.005074f
C454 XM1/a_n100_n8595# XM2/a_n100_n163411# 0.005243f
C455 XM1/a_100_2990# XM2/a_n100_n152867# 0.005074f
C456 XM4/w_n358_n132787# XM4/a_n100_105693# -0.004445f
C457 XM1/a_n158_116434# XM2/a_n158_n39422# 4.64e-21
C458 XM1/a_100_44634# XM2/a_n100_n108055# 0.005074f
C459 XM2/a_n158_n160678# m1_1634_n2388# 2.36e-21
C460 XM4/w_n358_n132787# XM3/a_n100_65289# 0.009186f
C461 XM4/w_n358_n132787# XM2/a_n100_n229311# 0.025061f
C462 XM4/w_n358_n132787# XM3/a_n158_n73438# 0.032295f
C463 XM1/a_n100_n113423# XM2/a_100_n266118# 7.26e-20
C464 XM4/a_n100_n60067# m1_1634_n2388# 0.072015f
C465 XM2/a_n100_26381# XM4/w_n358_n132787# 0.012096f
C466 XM4/w_n358_n132787# XM3/a_n100_10381# 0.009186f
C467 XM1/a_n100_n7159# XM2/a_100_n160678# 8.45e-20
C468 XM3/a_n158_129618# m1_1634_n2388# 6.1e-20
C469 XM1/a_100_n94658# XM4/w_n358_n132787# 0.054609f
C470 XM1/a_100_n22858# XM3/a_n100_29029# 2.85e-20
C471 XM1/a_n100_28741# XM3/a_n158_79890# 2.85e-20
C472 XM2/a_100_n287206# XM3/a_n158_n81726# 0.077916f
C473 XM4/w_n358_n132787# XM3/a_n100_102585# 0.009186f
C474 XM1/a_100_37454# XM2/a_100_n118502# 4.64e-21
C475 XM2/a_100_n329382# XM3/a_n100_n123263# 0.010147f
C476 XM2/a_n158_n200218# XM3/a_n158_6334# 4.64e-21
C477 XM2/a_100_n15698# XM1/a_n100_139313# 7.26e-20
C478 XM1/a_100_79098# XM4/w_n358_n132787# 0.054609f
C479 XM2/a_n100_n326843# XM3/a_n158_n122130# 0.005074f
C480 XM4/a_n100_n131551# XM4/w_n358_n132787# -0.004445f
C481 XM1/a_n100_n35879# XM4/w_n358_n132787# 0.013388f
C482 XM2/a_100_n105322# XM3/a_n100_100513# 0.010147f
C483 XM2/a_n158_n239758# XM3/a_n100_n35203# 7.26e-20
C484 XM4/w_n358_n132787# XM4/a_n100_66325# -0.004445f
C485 XM1/a_n100_n57419# XM3/a_n158_n5062# 2.85e-20
C486 XM3/a_n100_n40383# m1_1634_n2388# 0.072015f
C487 XM2/a_n158_n324110# XM3/a_n158_n116950# 4.64e-21
C488 XM2/a_100_n97414# m1_1634_n2388# 0.019728f
C489 XM1/a_n158_5862# XM3/a_n100_58037# 1.94e-20
C490 XM4/w_n358_n132787# XM3/a_n158_n112806# 0.032295f
C491 XM4/a_n100_n99435# m1_1634_n2388# 0.072015f
C492 XM2/a_100_n237122# XM3/a_n100_n30023# 0.005074f
C493 XM3/a_n100_48713# m1_1634_n2388# 0.072015f
C494 XM2/a_100_n10426# XM1/a_n100_145057# 7.26e-20
C495 XM4/w_n358_n132787# XM2/a_n158_n165950# 0.106739f
C496 XM1/a_n158_4426# XM3/a_n100_55965# 1.94e-20
C497 XM1/a_n100_47409# m1_1634_n2388# 1.3e-19
C498 XM2/a_n158_n284570# m1_1634_n2388# 2.36e-21
C499 XM1/a_n158_n77426# XM3/a_n100_n25879# 1.94e-20
C500 XM2/a_n100_n276759# XM3/a_n100_n70427# 8.38e-19
C501 XM2/a_100_n118502# XM3/a_n100_86009# 0.005074f
C502 XM4/w_n358_n132787# XM3/a_n158_90250# 0.032295f
C503 XM4/w_n358_n132787# XM3/a_n158_127546# 0.034847f
C504 XM1/a_n100_n160811# XM4/w_n358_n132787# 0.01363f
C505 XM4/w_n358_n132787# XM4/a_n100_n5159# -0.004445f
C506 XM1/a_100_103510# XM4/w_n358_n132787# 0.051269f
C507 XM2/a_n100_n86967# XM4/a_100_120294# 2.56e-20
C508 XM4/w_n358_n132787# XM3/a_n100_4165# 0.009093f
C509 XM2/a_100_n160678# XM3/a_n100_43533# 0.005074f
C510 XM4/w_n358_n132787# XM1/a_n100_n142143# 0.01363f
C511 XM4/w_n358_n132787# XM3/a_n158_35342# 0.036937f
C512 XM4/a_100_100610# m1_1634_n2388# 6.1e-20
C513 XM2/a_n100_n115963# XM3/a_n158_91286# 0.005074f
C514 XM1/a_n158_n53014# XM3/a_n100_n2051# 1.94e-20
C515 XM3/a_n100_3129# XM4/a_n100_3129# 0.009521f
C516 XM2/a_100_n86870# XM3/a_n158_118222# 0.077916f
C517 XM2/a_100_n268754# XM3/a_n158_n64114# 0.062337f
C518 XM1/a_n100_n99063# m1_1634_n2388# 8.14e-20
C519 XM4/w_n358_n132787# XM4/a_n100_26957# -0.004445f
C520 XM3/a_n100_n79751# m1_1634_n2388# 0.072015f
C521 XM2/a_n100_n274123# XM4/a_100_n69294# 1.79e-20
C522 XM2/a_100_n202854# XM3/a_n158_1154# 8.02e-19
C523 XM1/a_n100_20125# XM2/a_100_n134318# 1.45e-19
C524 XM2/a_100_n310930# XM3/a_n100_n105651# 0.010147f
C525 XM2/a_n100_n158139# XM3/a_n158_48810# 0.005074f
C526 XM1/a_n100_63205# XM2/a_100_n92142# 7.26e-20
C527 XM1/a_100_57558# XM4/w_n358_n132787# 0.053586f
C528 XM3/a_n100_91189# XM4/a_n100_91189# 0.009521f
C529 XM1/a_n100_n183787# XM2/a_n100_n337387# 0.006572f
C530 XM3/a_n100_n21735# XM4/a_n100_n21735# 0.009521f
C531 XM4/a_100_n918# m1_1634_n2388# 6.1e-20
C532 XM1/a_n100_15817# XM2/a_100_n136954# 7.26e-20
C533 XM1/a_n100_n142143# XM2/a_n158_n297750# 0.005074f
C534 XM1/a_100_n124814# XM3/a_n100_n73535# 5.71e-20
C535 XM1/a_n158_n113326# XM3/a_n100_n62139# 3.63e-20
C536 XM4/w_n358_n132787# XM2/a_100_n102686# 0.103341f
C537 XM1/a_n100_n170863# m1_1634_n2388# 1.3e-19
C538 XM2/a_100_n221306# m1_1634_n2388# 0.019664f
C539 XM1/a_100_n91786# m1_1634_n2388# 7.88e-19
C540 XM4/w_n358_n132787# XM4/a_n100_n44527# -0.004445f
C541 XM3/a_n158_n15422# m1_1634_n2388# 6.1e-20
C542 XM4/w_n358_n132787# XM2/a_n158_n289842# 0.101988f
C543 XM2/a_100_n218670# XM3/a_n100_n12411# 0.006179f
C544 XM1/a_100_n28602# XM3/a_n100_22813# 7.45e-19
C545 XM1/a_100_92022# XM2/a_100_n63146# 4.64e-21
C546 XM3/a_n158_73674# m1_1634_n2388# 6.1e-20
C547 XM4/a_100_61242# m1_1634_n2388# 6.1e-20
C548 XM1/a_100_n150662# XM2/a_100_n305658# 4.64e-21
C549 XM2/a_n100_n216131# XM3/a_n158_n11278# 0.001105f
C550 XM1/a_100_129358# XM2/a_100_n26242# 4.64e-21
C551 XM2/a_100_n147498# XM3/a_n100_58037# 0.010147f
C552 XM1/a_n100_n130655# m1_1634_n2388# 1.3e-19
C553 XM1/a_n158_48942# XM3/a_n100_99477# 1.94e-20
C554 XM3/a_n158_18766# m1_1634_n2388# 6.1e-20
C555 XM3/a_n100_n119119# m1_1634_n2388# 0.072015f
C556 XM1/a_n100_179521# XM2/a_n158_23842# 0.005074f
C557 XM1/a_n100_53153# XM2/a_100_n100050# 7.26e-20
C558 XM1/a_n100_n58855# XM2/a_100_n213398# 1.45e-19
C559 XM2/a_100_n189674# XM3/a_n100_15561# 0.010147f
C560 XM1/a_n100_n137835# XM2/a_n100_n292575# 0.001572f
C561 XM1/a_n158_n101838# XM2/a_n158_n255574# 9.28e-21
C562 XM3/a_n100_n41419# XM4/a_n100_n41419# 0.009521f
C563 XM1/a_100_162386# XM2/a_n158_8026# 0.116862f
C564 XM4/a_n100_124341# m1_1634_n2388# 0.072015f
C565 XM4/w_n358_n132787# XM3/a_n100_n24843# 0.009017f
C566 XM4/a_100_n10242# m1_1634_n2388# 6.1e-20
C567 XM1/a_100_2990# XM2/a_100_n150134# 4.64e-21
C568 XM2/a_100_n292478# XM3/a_n100_n88039# 0.005074f
C569 XM4/w_n358_n132787# XM1/a_n100_n149323# 0.01363f
C570 XM4/w_n358_n132787# XM4/a_n100_n83895# -0.004445f
C571 XM1/a_n100_n134963# XM3/a_n158_n82762# 7.81e-19
C572 XM3/a_n158_n54790# m1_1634_n2388# 6.1e-20
C573 XM2/a_n100_n160775# m1_1634_n2388# 0.001932f
C574 XM1/a_n100_n136399# XM2/a_n100_n292575# 7.47e-19
C575 XM4/w_n358_n132787# XM2/a_100_n226578# 0.105653f
C576 XM4/a_100_21874# m1_1634_n2388# 6.1e-20
C577 XM1/a_n100_n113423# XM2/a_n158_n266118# 0.005074f
C578 XM1/a_100_n83170# XM3/a_n100_n31059# 2.85e-20
C579 XM1/a_n100_n7159# XM2/a_n158_n160678# 0.005401f
C580 XM3/a_n100_129521# m1_1634_n2388# 0.072015f
C581 XM1/a_100_n153534# XM3/a_n100_n102543# 2.85e-20
C582 XM2/a_100_n134318# XM3/a_n100_72541# 0.005074f
C583 XM2/a_n100_n142323# XM4/a_100_62278# 2.56e-20
C584 XM1/a_100_37454# XM2/a_n158_n118502# 0.004307f
C585 XM2/a_n158_n329382# XM3/a_n100_n123263# 1.45e-19
C586 XM1/a_n158_n64502# XM2/a_n158_n218670# 9.28e-21
C587 XM2/a_n100_n200315# XM3/a_n158_6334# 0.005074f
C588 XM2/a_100_n176494# XM3/a_n100_30065# 0.005074f
C589 XM2/a_n158_n18334# XM1/a_n158_135102# 4.64e-21
C590 XM1/a_n100_113465# XM2/a_n158_n39422# 0.005074f
C591 XM3/a_n100_n61103# XM4/a_n100_n61103# 0.009521f
C592 XM1/a_100_21658# XM3/a_n158_72638# 0.00544f
C593 XM2/a_n100_n247763# XM4/a_n100_n41419# 4.28e-20
C594 XM1/a_n100_n1415# XM4/w_n358_n132787# 0.013436f
C595 XM1/a_100_n32910# XM4/w_n358_n132787# 0.048442f
C596 XM2/a_n158_n105322# XM3/a_n100_100513# 1.45e-19
C597 XM4/a_n100_84973# m1_1634_n2388# 0.072015f
C598 XM4/w_n358_n132787# XM3/a_n100_n64211# 0.008451f
C599 XM4/a_100_n49610# m1_1634_n2388# 6.1e-20
C600 XM4/a_n100_4165# m1_1634_n2388# 0.072015f
C601 XM1/a_100_143718# XM2/a_n158_n10426# 0.116862f
C602 XM1/a_n158_n167894# XM3/a_n100_n117047# 1.94e-20
C603 XM1/a_100_20222# XM3/a_n100_72541# 2.46e-20
C604 XM4/w_n358_n132787# XM4/a_n100_n123263# -0.004445f
C605 XM3/a_n158_n94158# m1_1634_n2388# 6.1e-20
C606 XM1/a_n100_n51675# XM3/a_n158_n918# 2.85e-20
C607 XM1/a_100_5862# XM3/a_n100_57001# 1.57e-19
C608 XM2/a_n100_n324207# XM3/a_n158_n116950# 0.005074f
C609 XM2/a_n158_n97414# m1_1634_n2388# 2.36e-21
C610 XM4/w_n358_n132787# XM3/a_n100_83937# 0.009186f
C611 XM2/a_n158_n237122# XM3/a_n100_n30023# 7.26e-20
C612 XM1/a_n100_n169427# XM3/a_n100_n119119# 0.001197f
C613 XM4/w_n358_n132787# XM2/a_n100_n166047# 0.025083f
C614 XM4/w_n358_n132787# XM3/a_n100_n2051# 0.00888f
C615 XM2/a_n100_n284667# m1_1634_n2388# 0.001365f
C616 XM1/a_100_n114762# XM3/a_n100_n64211# 2.85e-20
C617 XM4/w_n358_n132787# XM3/a_n100_29029# 0.009186f
C618 XM1/a_100_n5626# XM3/a_n158_46738# 7.57e-19
C619 XM1/a_100_n14242# XM3/a_n100_36281# 2.85e-20
C620 XM2/a_n158_n118502# XM3/a_n100_86009# 7.26e-20
C621 XM2/a_n100_n18431# XM1/a_100_135102# 0.005074f
C622 XM1/a_100_n116198# m1_1634_n2388# 1.82e-19
C623 XM1/a_n158_n68810# XM3/a_n100_n16555# 9.62e-21
C624 XM4/w_n358_n132787# XM3/a_n100_127449# 0.008419f
C625 XM3/a_n100_n80787# XM4/a_n100_n80787# 0.009521f
C626 XM2/a_n158_n160678# XM3/a_n100_43533# 7.26e-20
C627 XM3/a_n100_59073# XM4/a_n100_59073# 0.009521f
C628 XM4/a_n100_45605# m1_1634_n2388# 0.072015f
C629 XM4/w_n358_n132787# XM3/a_n100_n103579# 0.007888f
C630 XM4/a_100_n88978# m1_1634_n2388# 6.1e-20
C631 XM2/a_100_n113230# XM3/a_n158_91286# 0.050264f
C632 XM2/a_100_n86870# XM3/a_n100_118125# 0.010147f
C633 XM1/a_n100_25869# XM2/a_100_n126410# 5.46e-20
C634 XM2/a_n158_n268754# XM3/a_n158_n64114# 4.64e-21
C635 XM2/a_n158_n49966# XM4/w_n358_n132787# 0.101988f
C636 XM2/a_n158_n202854# XM3/a_n158_1154# 4.64e-21
C637 XM1/a_n100_63205# XM2/a_n158_n92142# 0.005074f
C638 XM1/a_n100_54589# XM2/a_100_n100050# 1.24e-19
C639 XM1/a_n100_20125# XM2/a_n158_n134318# 0.010147f
C640 XM2/a_n158_n310930# XM3/a_n100_n105651# 1.45e-19
C641 XM2/a_100_n155406# XM3/a_n158_48810# 0.021054f
C642 XM1/a_n100_n33007# m1_1634_n2388# 1.15e-19
C643 XM1/a_n100_15817# XM2/a_n158_n136954# 0.005074f
C644 pcbias XM4/w_n358_n132787# 0.003693f
C645 XM2/a_100_n266118# XM3/a_n158_n58934# 0.001581f
C646 XM1/a_n100_n38751# XM2/a_100_n192310# 1.18e-19
C647 XM3/a_n100_67361# m1_1634_n2388# 0.072014f
C648 XM2/a_n100_n271487# XM4/a_100_n64114# 5.53e-21
C649 XM1/a_n100_68949# XM2/a_100_n84234# 7.26e-20
C650 XM4/w_n358_n132787# XM2/a_n158_n102686# 0.107093f
C651 XM4/w_n358_n132787# XM3/a_n158_n39250# 0.032295f
C652 XM4/a_n100_n25879# m1_1634_n2388# 0.072015f
C653 XM1/a_n100_n153631# XM3/a_n158_n101410# 0.001453f
C654 XM1/a_n158_n70246# XM2/a_n158_n223942# 9.28e-21
C655 XM3/a_n100_12453# m1_1634_n2388# 0.072015f
C656 XM3/a_n100_n100471# XM4/a_n100_n100471# 0.009521f
C657 XM4/w_n358_n132787# XM2/a_n100_n289939# 0.025125f
C658 XM1/a_100_n28602# XM2/a_100_n184402# 4.64e-21
C659 XM2/a_n158_n218670# XM3/a_n100_n12411# 1.09e-19
C660 XM3/a_n158_105790# m1_1634_n2388# 6.1e-20
C661 XM4/a_100_n128346# m1_1634_n2388# 6.1e-20
C662 XM1/a_100_n150662# XM2/a_n158_n305658# 0.097778f
C663 XM2/a_n158_n147498# XM3/a_n100_58037# 1.45e-19
C664 XM1/a_100_n157842# XM3/a_n100_n106687# 4.46e-20
C665 XM4/w_n358_n132787# XM3/a_n158_53990# 0.038462f
C666 XM1/a_n158_125050# XM2/a_n158_n28878# 9.28e-21
C667 XM1/a_n100_53153# XM2/a_n158_n100050# 0.005074f
C668 XM2/a_n158_n189674# XM3/a_n100_15561# 1.45e-19
C669 XM4/w_n358_n132787# XM1/a_100_n160714# 0.055027f
C670 XM1/a_n100_n58855# XM2/a_n158_n213398# 0.010147f
C671 XM4/w_n358_n132787# XM4/a_n100_100513# -0.004445f
C672 XM2/a_n100_n213495# XM3/a_n158_n6098# 1.17e-21
C673 XM2/a_100_n142226# XM3/a_n158_63314# 0.077916f
C674 XM3/a_n100_n6195# m1_1634_n2388# 0.072015f
C675 XM1/a_100_143718# XM4/w_n358_n132787# 0.048442f
C676 XM4/w_n358_n132787# XM3/a_n158_n78618# 0.032295f
C677 XM4/a_n100_n65247# m1_1634_n2388# 0.072015f
C678 XM1/a_n158_n47270# XM2/a_n158_n200218# 4.64e-21
C679 XM2/a_100_n184402# XM3/a_n158_20838# 0.077916f
C680 XM1/a_100_2990# XM2/a_n158_n150134# 0.070516f
C681 XM2/a_n158_n292478# XM3/a_n100_n88039# 7.26e-20
C682 XM1/a_100_n117634# XM3/a_n100_n66283# 5.71e-20
C683 XM1/a_100_150898# XM4/w_n358_n132787# 0.052496f
C684 XM1/a_n100_81873# XM2/a_100_n73690# 7.26e-20
C685 XM3/a_n100_n120155# XM4/a_n100_n120155# 0.009521f
C686 XM2/a_100_n158042# m1_1634_n2388# 0.017213f
C687 XM1/a_100_33146# XM3/a_n100_83937# 2.85e-20
C688 XM1/a_n100_27305# XM3/a_n158_79890# 3.44e-21
C689 XM4/w_n358_n132787# XM4/a_n100_n1015# -0.004445f
C690 XM1/a_n100_n136399# XM2/a_100_n289842# 7.26e-20
C691 XM1/a_n100_n78959# m1_1634_n2388# 1.3e-19
C692 XM4/w_n358_n132787# XM2/a_n158_n226578# 0.101988f
C693 XM2/a_n100_n253035# XM4/a_100_n46502# 9.49e-21
C694 XM2/a_100_n247666# XM3/a_n158_n41322# 0.077916f
C695 XM1/a_n100_79001# XM2/a_n158_n73690# 0.005074f
C696 XM1/a_100_64738# XM3/a_n100_116053# 5.71e-20
C697 XM3/a_n158_92322# m1_1634_n2388# 6.1e-20
C698 XM1/a_n100_n7159# XM2/a_n100_n160775# 0.005243f
C699 XM1/a_100_24530# XM3/a_n158_75746# 3.04e-19
C700 XM2/a_100_n289842# XM3/a_n100_n82859# 0.005074f
C701 XM1/a_n100_116337# XM2/a_n158_n36786# 0.005074f
C702 XM2/a_n158_n134318# XM3/a_n100_72541# 7.26e-20
C703 XM1/a_100_n149226# XM3/a_n100_n98399# 2.85e-20
C704 XM1/a_n100_n124911# XM3/a_n158_n74474# 1.17e-20
C705 XM1/a_n158_n103274# XM3/a_n100_n51779# 2.1e-20
C706 XM1/a_n158_27402# XM3/a_n100_77721# 1.94e-20
C707 XM3/a_n158_37414# m1_1634_n2388# 6.1e-20
C708 XM4/w_n358_n132787# XM3/a_n158_103718# 0.032389f
C709 XM1/a_100_37454# XM2/a_n100_n118599# 0.005074f
C710 XM4/w_n358_n132787# XM4/a_n100_61145# -0.004445f
C711 XM1/a_100_n94658# XM3/a_n100_n43491# 4.82e-20
C712 XM2/a_n158_n176494# XM3/a_n100_30065# 7.26e-20
C713 XM3/a_n100_n45563# m1_1634_n2388# 0.072015f
C714 XM2/a_100_n129046# XM3/a_n158_77818# 0.032738f
C715 XM2/a_100_n105322# XM3/a_n158_101646# 0.022612f
C716 XM2/a_n100_n139687# XM4/a_100_67458# 2.56e-20
C717 XM4/w_n358_n132787# XM3/a_n158_n117986# 0.032295f
C718 XM4/a_n100_n104615# m1_1634_n2388# 0.072015f
C719 XM1/a_100_n169330# XM3/a_n100_n118083# 5.71e-20
C720 XM1/a_n100_n140707# XM3/a_n100_n89075# 8.46e-19
C721 XM1/a_n158_17350# XM3/a_n100_69433# 1.94e-20
C722 XM2/a_100_n171222# XM3/a_n158_35342# 0.061948f
C723 XM1/a_n100_n127783# XM3/a_n100_n76643# 2.68e-19
C724 XM1/a_100_n104710# XM3/a_n100_n52815# 2.85e-20
C725 XM1/a_n100_n91883# XM3/a_n158_n41322# 2.85e-20
C726 XM2/a_100_n321474# XM3/a_n158_n116950# 0.051043f
C727 XM2/a_n100_n326843# XM4/a_100_n122130# 2.56e-20
C728 XM1/a_n100_n96191# m1_1634_n2388# 1.07e-19
C729 XM1/a_n100_147929# XM2/a_n158_n7790# 0.005074f
C730 XM2/a_n100_n97511# m1_1634_n2388# 0.002024f
C731 XM1/a_n100_57461# XM4/w_n358_n132787# 0.012521f
C732 XM4/w_n358_n132787# XM4/a_n100_n10339# -0.004445f
C733 XM3/a_n100_26957# XM4/a_n100_26957# 0.009521f
C734 XM4/w_n358_n132787# XM2/a_100_n163314# 0.104031f
C735 XM1/a_n100_166597# XM2/a_n158_13298# 0.005074f
C736 XM2/a_100_n281934# m1_1634_n2388# 0.017213f
C737 XM4/a_100_95430# m1_1634_n2388# 6.1e-20
C738 XM4/w_n358_n132787# XM4/a_n100_21777# -0.004445f
C739 XM1/a_n100_n113423# XM3/a_n100_n63175# 2.42e-19
C740 XM1/a_n158_n94658# XM3/a_n100_n43491# 3.23e-20
C741 XM2/a_n100_n65879# XM4/w_n358_n132787# 0.012279f
C742 XM3/a_n100_n84931# m1_1634_n2388# 0.072015f
C743 XM2/a_100_n229214# XM3/a_n158_n23710# 0.077916f
C744 XM1/a_n158_69046# XM3/a_n100_120197# 2.91e-20
C745 XM2/a_100_n271390# XM3/a_n100_n65247# 0.010147f
C746 XM2/a_n158_n113230# XM3/a_n158_91286# 4.64e-21
C747 XM1/a_n100_n31571# XM3/a_n100_19705# 2.73e-19
C748 XM2/a_n158_n86870# XM3/a_n100_118125# 1.45e-19
C749 XM1/a_n100_25869# XM2/a_n158_n126410# 0.004594f
C750 XM2/a_n100_n268851# XM3/a_n158_n64114# 0.005074f
C751 XM2/a_n100_n202951# XM3/a_n158_1154# 0.005074f
C752 XM1/a_n100_n44495# XM4/w_n358_n132787# 0.01363f
C753 XM1/a_n100_54589# XM2/a_n158_n100050# 0.007937f
C754 XM2/a_n158_n155406# XM3/a_n158_48810# 4.64e-21
C755 XM1/a_n158_123614# XM2/a_n100_n28975# 7.26e-20
C756 XM4/w_n358_n132787# XM4/a_n100_n49707# -0.004445f
C757 XM3/a_n158_n20602# m1_1634_n2388# 6.1e-20
C758 XM1/a_n100_129261# XM4/w_n358_n132787# 0.012279f
C759 XM2/a_n158_n266118# XM3/a_n158_n58934# 4.64e-21
C760 XM1/a_n100_n38751# XM2/a_n158_n192310# 0.007234f
C761 XM1/a_n100_68949# XM2/a_n158_n84234# 0.005074f
C762 XM1/a_n100_n142143# XM2/a_100_n295114# 7.26e-20
C763 XM4/w_n358_n132787# XM2/a_n100_n102783# 0.024108f
C764 XM4/a_100_56062# m1_1634_n2388# 6.1e-20
C765 XM2/a_n100_n221403# m1_1634_n2388# 0.003195f
C766 XM4/w_n358_n132787# XM3/a_n100_47677# 0.009186f
C767 XM1/a_n100_n176607# XM4/w_n358_n132787# 0.0135f
C768 XM1/a_n100_n86139# XM3/a_n158_n34070# 2.85e-20
C769 XM1/a_100_n28602# XM2/a_n158_n184402# 0.019496f
C770 XM3/a_n100_n124299# m1_1634_n2388# 0.072015f
C771 XM4/w_n358_n132787# XM2/a_100_n287206# 0.103341f
C772 XM1/a_n100_n182351# XM2/a_100_n337290# 7.26e-20
C773 XM2/a_n100_n218767# XM3/a_n100_n12411# 0.002506f
C774 XM1/a_100_86278# XM2/a_n158_n68418# 0.116862f
C775 XM3/a_n100_105693# m1_1634_n2388# 0.072015f
C776 XM1/a_100_n150662# XM2/a_n100_n305755# 0.005074f
C777 XM1/a_100_81970# XM2/a_n158_n73690# 0.033127f
C778 XM1/a_n100_38793# XM3/a_n158_89214# 6.97e-21
C779 XM1/a_n100_119209# XM2/a_n158_n36786# 1.06e-19
C780 XM1/a_n158_84842# XM2/a_n100_n68515# 7.26e-20
C781 XM4/a_n100_119161# m1_1634_n2388# 0.072014f
C782 XM4/w_n358_n132787# XM3/a_n100_n30023# 0.009096f
C783 XM4/a_100_n15422# m1_1634_n2388# 6.1e-20
C784 XM2/a_n158_n2518# XM4/w_n358_n132787# 0.101988f
C785 XM1/a_100_123614# XM2/a_n100_n31611# 0.005074f
C786 XM1/a_n158_n163586# XM3/a_n100_n112903# 1.94e-20
C787 XM2/a_n100_n195043# XM4/a_100_9442# 2.56e-20
C788 XM2/a_n100_n216131# XM4/a_100_n11278# 1.16e-20
C789 XM2/a_100_n210762# XM3/a_n158_n6098# 0.064674f
C790 XM1/a_n158_119306# XM2/a_n100_n36883# 3.74e-21
C791 XM1/a_100_87714# XM2/a_100_n65782# 4.64e-21
C792 XM4/w_n358_n132787# XM4/a_n100_n89075# -0.004445f
C793 XM3/a_n158_n59970# m1_1634_n2388# 6.1e-20
C794 XM1/a_100_36018# XM3/a_n100_87045# 2.85e-20
C795 XM1/a_n158_n175074# XM2/a_n158_n329382# 9.28e-21
C796 XM2/a_100_n252938# XM3/a_n100_n47635# 0.010147f
C797 XM2/a_100_n208126# XM3/a_n158_n2990# 0.077916f
C798 XM4/a_100_16694# m1_1634_n2388# 6.1e-20
C799 XM1/a_n100_1457# XM2/a_100_n152770# 1.45e-19
C800 XM1/a_n158_n47270# XM2/a_n100_n200315# 7.26e-20
C801 XM3/a_n100_86009# m1_1634_n2388# 0.072015f
C802 XM1/a_n158_n54450# XM3/a_n100_n2051# 2e-22
C803 XM4/w_n358_n132787# XM3/a_n158_5298# 0.032295f
C804 XM1/a_100_2990# XM2/a_n100_n150231# 0.005074f
C805 XM1/a_n158_31710# XM3/a_n100_82901# 3.71e-20
C806 XM1/a_100_n179382# XM4/w_n358_n132787# 0.055057f
C807 XM1/a_n100_n119167# XM3/a_n158_n68258# 2.85e-20
C808 XM1/a_n158_n61630# XM3/a_n100_n10339# 3.89e-20
C809 XM1/a_n100_n58855# XM3/a_n158_n7134# 7.86e-21
C810 XM3/a_n100_31101# m1_1634_n2388# 0.072015f
C811 XM1/a_n100_n136399# XM2/a_n158_n289842# 0.005074f
C812 XM4/w_n358_n132787# XM2/a_n100_n226675# 0.024087f
C813 XM1/a_n100_n157939# XM3/a_n100_n106687# 5.85e-19
C814 XM1/a_n100_2893# XM4/w_n358_n132787# 0.01363f
C815 XM3/a_n158_130654# m1_1634_n2388# 6.1e-20
C816 XM2/a_n158_n289842# XM3/a_n100_n82859# 7.26e-20
C817 XM4/w_n358_n132787# XM3/a_n100_103621# 0.007547f
C818 XM4/a_n100_79793# m1_1634_n2388# 0.072015f
C819 XM4/w_n358_n132787# XM3/a_n158_72638# 0.038462f
C820 XM4/w_n358_n132787# XM3/a_n100_n69391# 0.009997f
C821 XM4/a_100_n54790# m1_1634_n2388# 6.1e-20
C822 XM1/a_100_176746# XM2/a_n158_21206# 0.044811f
C823 XM1/a_100_37454# XM2/a_100_n115866# 4.64e-21
C824 XM1/a_n100_n25827# XM4/w_n358_n132787# 0.012832f
C825 XM4/w_n358_n132787# XM4/a_n100_n128443# -0.004445f
C826 XM3/a_n158_n99338# m1_1634_n2388# 6.1e-20
C827 XM4/w_n358_n132787# XM3/a_n158_17730# 0.03327f
C828 XM1/a_100_104946# XM2/a_n100_n50063# 0.005074f
C829 XM3/a_n100_79793# XM4/a_n100_79793# 0.009521f
C830 XM2/a_n158_n129046# XM3/a_n158_77818# 4.64e-21
C831 XM2/a_100_n105322# XM3/a_n100_101549# 0.005074f
C832 XM2/a_n158_n105322# XM3/a_n158_101646# 4.64e-21
C833 XM1/a_100_13042# XM3/a_n158_64350# 0.003891f
C834 XM1/a_n100_n50239# m1_1634_n2388# 9.19e-20
C835 XM1/a_n158_15914# XM3/a_n100_66325# 1.94e-20
C836 XM1/a_n100_11509# XM3/a_n158_62278# 2.85e-20
C837 XM1/a_100_n18550# XM2/a_100_n173858# 4.64e-21
C838 XM2/a_n158_n171222# XM3/a_n158_35342# 4.64e-21
C839 XM1/a_100_34582# XM2/a_100_n121138# 4.64e-21
C840 XM2/a_n158_n321474# XM3/a_n158_n116950# 4.64e-21
C841 XM4/w_n358_n132787# XM3/a_n158_n5062# 0.032295f
C842 XM2/a_100_n94778# m1_1634_n2388# 0.017213f
C843 XM1/a_n100_53153# XM3/a_n100_104657# 6.5e-21
C844 XM1/a_n158_n2754# XM3/a_n100_48713# 2.67e-20
C845 XM1/a_n100_172341# XM2/a_100_18570# 1.45e-19
C846 XM1/a_n100_n87575# XM3/a_n100_n37275# 7.19e-19
C847 XM1/a_n100_n80395# XM3/a_n158_n27854# 1.64e-20
C848 XM2/a_100_n234486# XM3/a_n100_n30023# 0.005074f
C849 XM4/w_n358_n132787# XM2/a_n158_n163314# 0.101988f
C850 XM4/a_n100_40425# m1_1634_n2388# 0.072015f
C851 XM2/a_100_n318838# XM3/a_n158_n111770# 0.012875f
C852 XM4/w_n358_n132787# XM3/a_n100_n108759# 0.009186f
C853 XM4/a_100_n94158# m1_1634_n2388# 6.1e-20
C854 XM2/a_n100_n324207# XM4/a_100_n116950# 2.56e-20
C855 XM4/w_n358_n132787# XM3/a_n158_128582# 0.032295f
C856 XM1/a_n100_61769# XM3/a_n158_113042# 7.86e-21
C857 XM1/a_n100_45973# m1_1634_n2388# 8.14e-20
C858 XM1/a_n100_n126347# XM4/w_n358_n132787# 0.01363f
C859 XM3/a_n158_56062# m1_1634_n2388# 6.1e-20
C860 XM1/a_n158_n165022# XM3/a_n100_n113939# 1.94e-20
C861 XM2/a_n100_n84331# XM4/a_100_120294# 2.56e-20
C862 XM1/a_100_n126250# m1_1634_n2388# 0.002183f
C863 XM1/a_100_25966# XM2/a_100_n129046# 4.64e-21
C864 XM2/a_n158_n271390# XM3/a_n100_n65247# 1.45e-19
C865 XM1/a_n100_142185# XM2/a_100_n10426# 7.26e-20
C866 XM2/a_n100_n113327# XM3/a_n158_91286# 0.005074f
C867 XM1/a_n100_99105# XM4/w_n358_n132787# 0.012279f
C868 XM2/a_100_n86870# XM3/a_n158_119258# 0.077916f
C869 XM1/a_n158_58994# XM2/a_n158_n94778# 9.28e-21
C870 XM1/a_n100_25869# XM2/a_n100_n126507# 7.46e-19
C871 XM1/a_100_n175074# XM2/a_n158_n329382# 0.116862f
C872 XM1/a_100_n51578# XM4/w_n358_n132787# 0.048442f
C873 XM1/a_100_171002# XM2/a_n100_18473# 0.005074f
C874 XM1/a_n100_63205# XM2/a_100_n89506# 7.26e-20
C875 XM1/a_n100_54589# XM2/a_n100_n100147# 0.001385f
C876 XM4/w_n358_n132787# XM3/a_n158_n44430# 0.032295f
C877 XM4/a_n100_n31059# m1_1634_n2388# 0.072015f
C878 XM2/a_n100_n155503# XM3/a_n158_48810# 0.005074f
C879 XM1/a_n158_n152098# XM3/a_n158_n101410# 2.84e-22
C880 XM1/a_n100_n81831# XM3/a_n158_n29926# 2.85e-20
C881 XM2/a_n100_n266215# XM3/a_n158_n58934# 0.005074f
C882 XM1/a_n100_n38751# XM2/a_n100_n192407# 0.001266f
C883 XM1/a_n100_n142143# XM2/a_n158_n295114# 0.005074f
C884 XM4/w_n358_n132787# XM2/a_100_n100050# 0.10336f
C885 XM2/a_100_n218670# m1_1634_n2388# 0.019664f
C886 XM1/a_n100_18689# XM2/a_100_n136954# 7.26e-20
C887 XM1/a_n100_n110551# XM4/w_n358_n132787# 0.013509f
C888 XM1/a_100_n28602# XM2/a_n100_n184499# 0.005074f
C889 XM4/w_n358_n132787# XM2/a_n158_n287206# 0.105974f
C890 XM1/a_n100_n73215# XM3/a_n158_n22674# 0.001222f
C891 XM1/a_n100_n182351# XM2/a_n158_n337290# 0.005074f
C892 XM2/a_n100_n18431# XM4/w_n358_n132787# 0.01219f
C893 XM4/w_n358_n132787# XM4/a_n100_95333# -0.004445f
C894 XM1/a_100_15914# XM2/a_100_n139590# 4.64e-21
C895 XM3/a_n100_n11375# m1_1634_n2388# 0.072015f
C896 XM1/a_n158_53250# XM2/a_n158_n102686# 4.64e-21
C897 XM2/a_100_n300386# XM3/a_n158_n94158# 0.077916f
C898 XM4/w_n358_n132787# XM3/a_n158_n83798# 0.032295f
C899 XM4/a_n100_n70427# m1_1634_n2388# 0.072015f
C900 XM2/a_n158_n210762# XM3/a_n158_n6098# 4.64e-21
C901 XM4/w_n358_n132787# XM3/a_n158_n918# 0.038241f
C902 XM1/a_n100_n107679# XM3/a_n158_n56862# 2.85e-20
C903 XM1/a_n100_n64599# XM3/a_n100_n13447# 6.24e-19
C904 XM1/a_100_153770# XM4/w_n358_n132787# 0.048442f
C905 XM2/a_n158_n252938# XM3/a_n100_n47635# 1.45e-19
C906 XM1/a_n158_n8498# XM2/a_n158_n163314# 4.64e-21
C907 XM1/a_n100_1457# XM2/a_n158_n152770# 0.010147f
C908 XM3/a_n100_117089# XM4/a_n100_117089# 0.009521f
C909 XM2/a_n100_n192407# XM4/a_100_14622# 2.56e-20
C910 XM1/a_n100_n97627# XM4/w_n358_n132787# 0.01363f
C911 XM2/a_n100_n158139# m1_1634_n2388# 0.001749f
C912 XM1/a_n158_116434# XM2/a_n158_n36786# 4.64e-21
C913 XM4/a_100_129618# m1_1634_n2388# 6.1e-20
C914 XM1/a_n100_n132091# XM3/a_n158_n79654# 2.85e-20
C915 XM4/w_n358_n132787# XM3/a_n100_66325# 0.009186f
C916 XM1/a_n100_112029# XM2/a_n158_n42058# 0.010147f
C917 XM1/a_n100_n136399# XM2/a_n100_n289939# 0.001572f
C918 XM4/w_n358_n132787# XM2/a_100_n223942# 0.103341f
C919 XM2/a_n158_26478# XM1/a_n158_181054# 9.28e-21
C920 XM2/a_100_26478# XM1/a_n100_180957# 1.45e-19
C921 XM4/w_n358_n132787# XM4/a_n100_55965# -0.004445f
C922 XM3/a_n100_47677# XM4/a_n100_47677# 0.009521f
C923 XM2/a_n100_29017# XM4/w_n358_n132787# 0.006139f
C924 XM1/a_n100_n149323# XM3/a_n158_n97266# 2.85e-20
C925 XM3/a_n100_n50743# m1_1634_n2388# 0.072015f
C926 XM4/w_n358_n132787# XM3/a_n100_11417# 0.009973f
C927 XM3/a_n100_130557# m1_1634_n2388# 0.072015f
C928 XM1/a_n158_41762# XM2/a_n158_n113230# 4.64e-21
C929 XM1/a_n100_28741# XM3/a_n158_80926# 2.85e-20
C930 XM2/a_100_n131682# XM3/a_n100_72541# 0.005074f
C931 XM4/w_n358_n132787# XM3/a_n158_n123166# 0.032295f
C932 XM4/a_n100_n109795# m1_1634_n2388# 0.072015f
C933 XM3/a_n100_n7231# XM4/a_n100_n7231# 0.009521f
C934 XM2/a_n100_n197679# XM3/a_n158_6334# 4.8e-19
C935 XM2/a_100_n13062# XM1/a_n100_139313# 7.26e-20
C936 XM1/a_100_37454# XM2/a_n158_n115866# 0.0896f
C937 XM2/a_100_n173858# XM3/a_n100_30065# 0.005074f
C938 XM1/a_n100_n12903# XM3/a_n100_37317# 1.01e-20
C939 XM1/a_100_n74554# XM3/a_n100_n23807# 2.85e-20
C940 XM1/a_n100_110593# XM2/a_100_n44694# 7.26e-20
C941 XM1/a_n100_71821# m1_1634_n2388# 5.9e-20
C942 XM2/a_n100_n129143# XM3/a_n158_77818# 0.005074f
C943 XM2/a_n100_n105419# XM3/a_n158_101646# 0.005074f
C944 XM2/a_n158_n105322# XM3/a_n100_101549# 7.26e-20
C945 XM1/a_n100_n146451# XM3/a_n158_n94158# 2.85e-20
C946 XM2/a_100_n281934# XM3/a_n158_n76546# 0.077916f
C947 XM4/w_n358_n132787# XM4/a_n100_n15519# -0.004445f
C948 XM2/a_100_n324110# XM3/a_n100_n118083# 0.010147f
C949 XM1/a_100_n150662# m1_1634_n2388# 0.002062f
C950 XM1/a_100_n18550# XM2/a_n158_n173858# 0.0674f
C951 XM2/a_n100_n171319# XM3/a_n158_35342# 0.005074f
C952 XM4/a_100_90250# m1_1634_n2388# 6.1e-20
C953 XM1/a_n100_n139271# XM3/a_n158_n86906# 2.85e-20
C954 XM1/a_100_34582# XM2/a_n158_n121138# 0.027285f
C955 XM2/a_n100_n321571# XM3/a_n158_n116950# 0.005074f
C956 XM1/a_n158_n78862# XM2/a_n158_n234486# 4.64e-21
C957 XM1/a_n158_48942# XM3/a_n100_100513# 1.94e-20
C958 XM4/w_n358_n132787# XM4/a_n100_16597# -0.004445f
C959 XM1/a_n100_17253# m1_1634_n2388# 1.02e-19
C960 XM2/a_n158_n234486# XM3/a_n100_n30023# 7.26e-20
C961 XM3/a_n100_49749# m1_1634_n2388# 0.072015f
C962 XM2/a_100_n7790# XM1/a_n100_145057# 7.26e-20
C963 XM3/a_n100_n90111# m1_1634_n2388# 0.072015f
C964 XM4/w_n358_n132787# XM2/a_n100_n163411# 0.025107f
C965 XM1/a_n158_n58758# XM2/a_n158_n213398# 9.28e-21
C966 XM1/a_100_4426# XM3/a_n100_54929# 2.85e-20
C967 XM2/a_n100_n282031# m1_1634_n2388# 0.001951f
C968 XM2/a_n158_n318838# XM3/a_n158_n111770# 4.64e-21
C969 XM1/a_n100_n100499# XM2/a_100_n255574# 7.26e-20
C970 XM1/a_100_n42962# XM2/a_n158_n197582# 0.116862f
C971 XM4/w_n358_n132787# XM3/a_n158_91286# 0.038786f
C972 XM2/a_100_n118502# XM3/a_n100_87045# 0.010147f
C973 XM3/a_n100_n26915# XM4/a_n100_n26915# 0.009521f
C974 XM2/a_100_n231850# XM3/a_n100_n24843# 0.005074f
C975 XM4/w_n358_n132787# XM3/a_n100_128485# 0.009186f
C976 XM1/a_n100_71821# XM3/a_n158_122366# 0.001033f
C977 XM1/a_n100_61769# XM3/a_n100_112945# 7.98e-19
C978 XM3/a_n100_100513# XM4/a_n100_100513# 0.009521f
C979 XM1/a_100_n156406# XM3/a_n100_n105651# 2.85e-20
C980 XM1/a_100_n18550# XM4/w_n358_n132787# 0.054609f
C981 XM2/a_100_n160678# XM3/a_n100_44569# 0.010147f
C982 XM4/w_n358_n132787# XM3/a_n158_36378# 0.032295f
C983 XM1/a_100_25966# XM2/a_n158_n129046# 0.09622f
C984 XM4/w_n358_n132787# XM1/a_n100_n150759# 0.012584f
C985 XM4/w_n358_n132787# XM4/a_n100_n54887# -0.004445f
C986 XM3/a_n158_n25782# m1_1634_n2388# 6.1e-20
C987 XM2/a_100_n86870# XM3/a_n100_119161# 0.010147f
C988 XM1/a_n158_n183690# XM3/a_n100_n132587# 1.94e-20
C989 XM1/a_100_n170766# XM4/w_n358_n132787# 0.054609f
C990 XM4/a_100_50882# m1_1634_n2388# 6.1e-20
C991 XM2/a_n100_n81695# XM4/a_100_125474# 2.56e-20
C992 XM1/a_n100_63205# XM2/a_n158_n89506# 0.005074f
C993 XM1/a_n158_n55886# XM2/a_n158_n210762# 4.64e-21
C994 XM1/a_100_41762# m1_1634_n2388# 2.75e-22
C995 XM1/a_n100_n178043# XM3/a_n158_n127310# 2.85e-20
C996 XM3/a_n100_n129479# m1_1634_n2388# 0.072015f
C997 XM1/a_100_n48706# XM3/a_n100_3129# 2.85e-20
C998 XM2/a_n100_n268851# XM4/a_100_n64114# 2.56e-20
C999 XM2/a_100_n263482# XM3/a_n158_n58934# 0.053379f
C1000 XM1/a_n158_127922# XM2/a_n158_n26242# 9.28e-21
C1001 XM4/w_n358_n132787# XM2/a_n158_n100050# 0.103141f
C1002 XM1/a_n100_n162247# m1_1634_n2388# 8.14e-20
C1003 XM2/a_100_n305658# XM3/a_n100_n100471# 0.010147f
C1004 XM1/a_n158_n41526# XM2/a_n100_n197679# 3.46e-20
C1005 XM3/a_n100_n46599# XM4/a_n100_n46599# 0.009521f
C1006 XM1/a_n100_93361# XM4/w_n358_n132787# 0.012279f
C1007 XM1/a_n100_18689# XM2/a_n158_n136954# 0.005074f
C1008 XM1/a_100_n28602# XM2/a_100_n181766# 4.64e-21
C1009 XM4/a_n100_113981# m1_1634_n2388# 0.072015f
C1010 XM1/a_100_n173638# XM3/a_n100_n123263# 2.85e-20
C1011 XM4/w_n358_n132787# XM2/a_n100_n287303# 0.025201f
C1012 XM1/a_n100_173777# XM4/w_n358_n132787# 0.012279f
C1013 XM4/w_n358_n132787# XM3/a_n100_n35203# 0.008376f
C1014 XM4/a_100_n20602# m1_1634_n2388# 6.1e-20
C1015 XM1/a_100_92022# XM2/a_100_n60510# 4.64e-21
C1016 XM3/a_n158_74710# m1_1634_n2388# 6.1e-20
C1017 XM3/a_n158_106826# m1_1634_n2388# 6.1e-20
C1018 XM1/a_100_15914# XM2/a_n158_n139590# 0.048316f
C1019 XM1/a_100_129358# XM2/a_100_n23606# 4.64e-21
C1020 XM2/a_100_n147498# XM3/a_n100_59073# 0.005074f
C1021 XM4/w_n358_n132787# XM4/a_n100_n94255# -0.004445f
C1022 XM3/a_n158_n65150# m1_1634_n2388# 6.1e-20
C1023 XM1/a_n158_53250# XM2/a_n100_n102783# 7.26e-20
C1024 XM3/a_n158_19802# m1_1634_n2388# 6.1e-20
C1025 XM1/a_100_126486# XM2/a_100_n28878# 4.64e-21
C1026 XM1/a_n100_45973# XM3/a_n100_98441# 8.85e-19
C1027 XM2/a_100_n213398# XM3/a_n100_n7231# 0.010147f
C1028 XM4/a_100_11514# m1_1634_n2388# 6.1e-20
C1029 XM1/a_n100_179521# XM2/a_n158_26478# 0.005074f
C1030 XM1/a_100_11606# XM2/a_n158_n142226# 0.116862f
C1031 XM2/a_100_n189674# XM3/a_n100_16597# 0.005724f
C1032 XM1/a_100_46070# XM3/a_n100_96369# 2.82e-20
C1033 XM4/w_n358_n132787# XM1/a_100_n157842# 0.054609f
C1034 XM2/a_n100_n210859# XM3/a_n158_n6098# 0.005074f
C1035 XM1/a_100_n90350# XM3/a_n100_n39347# 2.85e-20
C1036 XM1/a_n158_n71682# XM3/a_n100_n19663# 1.94e-20
C1037 XM1/a_100_n63066# XM3/a_n100_n12411# 0.001486f
C1038 XM3/a_n100_15561# XM4/a_n100_15561# 0.009521f
C1039 XM1/a_n158_n8498# XM2/a_n100_n163411# 1.2e-20
C1040 XM1/a_n100_n55983# XM3/a_n158_n5062# 2.85e-20
C1041 XM3/a_n100_n66283# XM4/a_n100_n66283# 0.009521f
C1042 XM1/a_100_117870# XM4/w_n358_n132787# 0.048442f
C1043 XM2/a_100_n155406# m1_1634_n2388# 0.021162f
C1044 XM2/a_100_n73690# m1_1634_n2388# 0.008614f
C1045 XM4/a_n100_74613# m1_1634_n2388# 0.072015f
C1046 XM4/w_n358_n132787# XM1/a_n100_n139271# 0.013423f
C1047 XM4/w_n358_n132787# XM3/a_n100_n74571# 0.00821f
C1048 XM4/a_100_n59970# m1_1634_n2388# 6.1e-20
C1049 XM4/w_n358_n132787# XM2/a_n158_n223942# 0.103555f
C1050 XM1/a_100_64738# XM3/a_n100_117089# 1.52e-20
C1051 XM3/a_n158_n104518# m1_1634_n2388# 6.1e-20
C1052 XM1/a_n158_n34346# XM2/a_n158_n189674# 4.64e-21
C1053 XM1/a_n158_41762# XM2/a_n100_n113327# 7.26e-20
C1054 XM2/a_100_n287206# XM3/a_n100_n82859# 0.005074f
C1055 XM1/a_n158_n91786# XM2/a_n158_n247666# 4.64e-21
C1056 XM2/a_n158_n131682# XM3/a_n100_72541# 7.26e-20
C1057 XM4/w_n358_n132787# XM3/a_n158_104754# 0.032295f
C1058 XM1/a_n100_n14339# XM4/w_n358_n132787# 0.0135f
C1059 XM1/a_n100_83309# XM4/w_n358_n132787# 0.012279f
C1060 XM1/a_100_37454# XM2/a_n100_n115963# 0.005074f
C1061 XM2/a_n158_n173858# XM3/a_n100_30065# 7.26e-20
C1062 XM1/a_n158_n90350# XM3/a_n100_n39347# 1.94e-20
C1063 XM4/w_n358_n132787# XM3/a_n158_n10242# 0.032295f
C1064 XM2/a_100_n126410# XM3/a_n158_77818# 0.022222f
C1065 XM2/a_100_n102686# XM3/a_n158_101646# 0.032348f
C1066 XM2/a_n100_n137051# XM4/a_100_67458# 2.56e-20
C1067 pbias pcbias 0.060867f
C1068 XM1/a_n100_n63163# XM3/a_n158_n12314# 2.85e-20
C1069 XM1/a_n100_n57419# XM3/a_n100_n6195# 8.12e-19
C1070 XM3/a_n100_n85967# XM4/a_n100_n85967# 0.009521f
C1071 XM1/a_n100_n53111# XM3/a_n158_n1954# 2.85e-20
C1072 XM1/a_n158_53250# XM3/a_n100_103621# 8.02e-22
C1073 XM2/a_n158_n324110# XM3/a_n100_n118083# 1.45e-19
C1074 XM1/a_100_n18550# XM2/a_n100_n173955# 0.005074f
C1075 XM1/a_100_5862# XM3/a_n100_58037# 2.85e-20
C1076 XM1/a_n158_n142046# XM3/a_n100_n90111# 1.94e-20
C1077 XM4/a_n100_35245# m1_1634_n2388# 0.072015f
C1078 XM1/a_100_34582# XM2/a_n100_n121235# 0.005074f
C1079 XM4/w_n358_n132787# XM3/a_n100_n113939# 0.009036f
C1080 XM4/a_100_n99338# m1_1634_n2388# 6.1e-20
C1081 XM1/a_n158_n78862# XM2/a_n100_n234583# 7.26e-20
C1082 XM1/a_n158_n22858# XM2/a_n158_n176494# 9.28e-21
C1083 XM2/a_n100_n94875# m1_1634_n2388# 8.05e-19
C1084 XM4/w_n358_n132787# XM3/a_n100_84973# 0.009186f
C1085 XM1/a_n158_176746# XM2/a_n158_21206# 4.64e-21
C1086 XM1/a_n158_2990# XM3/a_n100_53893# 1.94e-20
C1087 XM4/w_n358_n132787# XM2/a_100_n160678# 0.103535f
C1088 XM2/a_100_n279298# m1_1634_n2388# 0.018653f
C1089 XM4/w_n358_n132787# XM3/a_n100_30065# 0.008928f
C1090 XM1/a_100_n18550# XM3/a_n158_33270# 0.00544f
C1091 XM1/a_100_n14242# XM3/a_n100_37317# 2.85e-20
C1092 XM4/w_n358_n132787# XM4/a_n100_129521# -0.004445f
C1093 XM2/a_n100_n318935# XM3/a_n158_n111770# 0.005074f
C1094 XM1/a_n100_n100499# XM2/a_n158_n255574# 0.005074f
C1095 XM2/a_n158_n118502# XM3/a_n100_87045# 1.45e-19
C1096 XM2/a_n158_n231850# XM3/a_n100_n24843# 7.26e-20
C1097 XM1/a_n100_168033# XM2/a_n158_13298# 0.005074f
C1098 XM1/a_n158_n127686# XM3/a_n100_n75607# 1.94e-20
C1099 XM1/a_n100_149365# XM4/w_n358_n132787# 0.012279f
C1100 XM4/w_n358_n132787# XM3/a_n158_n49610# 0.032295f
C1101 XM4/a_n100_n36239# m1_1634_n2388# 0.072014f
C1102 XM2/a_n158_n160678# XM3/a_n100_44569# 1.45e-19
C1103 XM1/a_n158_103510# XM2/a_n158_n49966# 4.64e-21
C1104 XM1/a_n158_69046# XM3/a_n100_121233# 1.94e-20
C1105 XM1/a_100_25966# XM2/a_n100_n129143# 0.005074f
C1106 XM1/a_n100_99105# XM2/a_n158_n55238# 0.010147f
C1107 XM2/a_100_n113230# XM3/a_n158_92322# 0.077916f
C1108 XM3/a_n100_n105651# XM4/a_n100_n105651# 0.009521f
C1109 XM2/a_n158_n86870# XM3/a_n100_119161# 1.45e-19
C1110 XM2/a_n158_n47330# XM4/w_n358_n132787# 0.104266f
C1111 XM1/a_n100_56025# XM4/w_n358_n132787# 0.014434f
C1112 XM1/a_n158_n55886# XM2/a_n100_n210859# 6.08e-20
C1113 XM2/a_100_n155406# XM3/a_n158_49846# 0.077916f
C1114 XM3/a_n100_7273# m1_1634_n2388# 0.072015f
C1115 XM2/a_n158_n263482# XM3/a_n158_n58934# 4.64e-21
C1116 XM1/a_100_155206# XM2/a_100_118# 4.64e-21
C1117 XM3/a_n100_68397# m1_1634_n2388# 0.072015f
C1118 XM4/w_n358_n132787# XM2/a_n100_n100147# 0.024957f
C1119 XM4/w_n358_n132787# XM4/a_n100_90153# -0.004445f
C1120 XM2/a_n158_n305658# XM3/a_n100_n100471# 1.45e-19
C1121 XM2/a_n100_n218767# m1_1634_n2388# 0.003067f
C1122 XM3/a_n100_n16555# m1_1634_n2388# 0.072015f
C1123 XM1/a_n100_n21519# XM3/a_n100_30065# 0.001054f
C1124 XM3/a_n100_13489# m1_1634_n2388# 0.072015f
C1125 XM1/a_100_n28602# XM2/a_n158_n181766# 0.074411f
C1126 XM1/a_n158_n172202# XM3/a_n100_n121191# 1.94e-20
C1127 XM4/w_n358_n132787# XM2/a_100_n284570# 0.104891f
C1128 XM1/a_n100_n182351# XM2/a_100_n334654# 7.26e-20
C1129 XM4/w_n358_n132787# XM3/a_n158_n88978# 0.032295f
C1130 XM4/a_n100_n75607# m1_1634_n2388# 0.072015f
C1131 XM2/a_n100_n266215# XM4/a_100_n58934# 2.56e-20
C1132 XM2/a_100_n260846# XM3/a_n158_n53754# 0.010539f
C1133 XM3/a_n100_106729# m1_1634_n2388# 0.072015f
C1134 XM1/a_100_15914# XM2/a_n100_n139687# 0.005074f
C1135 XM1/a_100_n150662# XM2/a_n100_n303119# 0.004271f
C1136 XM1/a_n158_n91786# XM3/a_n100_n41419# 1.12e-20
C1137 XM4/w_n358_n132787# XM3/a_n158_55026# 0.032295f
C1138 XM3/a_n100_68397# XM4/a_n100_68397# 0.009521f
C1139 XM2/a_n158_n147498# XM3/a_n100_59073# 7.26e-20
C1140 XM3/a_n100_n125335# XM4/a_n100_n125335# 0.009521f
C1141 XM1/a_n100_10073# XM2/a_100_n144862# 7.26e-20
C1142 XM1/a_100_40326# XM3/a_n158_91286# 0.001549f
C1143 XM1/a_n100_n116295# m1_1634_n2388# 1.3e-19
C1144 XM2/a_n158_n213398# XM3/a_n100_n7231# 1.45e-19
C1145 XM2/a_n158_n189674# XM3/a_n100_16597# 9.65e-20
C1146 XM1/a_100_n142046# XM3/a_n100_n91147# 2.85e-20
C1147 XM1/a_n100_87617# XM4/w_n358_n132787# 0.011915f
C1148 XM4/a_100_124438# m1_1634_n2388# 6.1e-20
C1149 XM2/a_100_n142226# XM3/a_n158_64350# 0.060779f
C1150 XM1/a_n158_43198# XM2/a_n158_n110594# 9.28e-21
C1151 XM1/a_n158_112126# XM2/a_n158_n42058# 9.28e-21
C1152 XM4/w_n358_n132787# XM4/a_n100_50785# -0.004445f
C1153 XM2/a_100_n184402# XM3/a_n158_21874# 0.077916f
C1154 XM3/a_n100_n55923# m1_1634_n2388# 0.072015f
C1155 XM1/a_n158_n12806# XM2/a_n158_n168586# 4.64e-21
C1156 XM1/a_n158_n2754# XM2/a_n158_n158042# 4.64e-21
C1157 XM1/a_n100_81873# XM2/a_100_n71054# 7.26e-20
C1158 XM2/a_100_n334654# XM3/a_n158_n129382# 0.077916f
C1159 XM2/a_n158_n155406# m1_1634_n2388# 2.36e-21
C1160 XM1/a_100_33146# XM3/a_n100_84973# 2.85e-20
C1161 XM1/a_n158_n143482# XM3/a_n100_n91147# 1.3e-20
C1162 XM1/a_n100_54589# XM3/a_n158_105790# 2.84e-20
C1163 XM4/w_n358_n132787# XM3/a_n158_n128346# 0.032295f
C1164 XM4/a_n100_n114975# m1_1634_n2388# 0.072015f
C1165 XM4/w_n358_n132787# XM2/a_n100_n224039# 0.024769f
C1166 XM2/a_100_n18334# XM1/a_n100_136441# 7.26e-20
C1167 XM2/a_100_n20970# XM1/a_n100_135005# 2.27e-20
C1168 XM3/a_n158_93358# m1_1634_n2388# 6.1e-20
C1169 XM1/a_n158_n34346# XM2/a_n100_n189771# 7.26e-20
C1170 XM3/a_n158_131690# m1_1634_n2388# 3.05e-20
C1171 XM2/a_n158_n287206# XM3/a_n100_n82859# 7.26e-20
C1172 XM1/a_n158_n91786# XM2/a_n100_n247763# 7.26e-20
C1173 XM1/a_n100_74693# m1_1634_n2388# 1.3e-19
C1174 XM1/a_n158_27402# XM3/a_n100_78757# 3.89e-20
C1175 XM4/w_n358_n132787# XM3/a_n100_104657# 0.007543f
C1176 XM1/a_n158_36018# XM2/a_n158_n118502# 9.28e-21
C1177 XM4/w_n358_n132787# XM1/a_n100_n157939# 0.013487f
C1178 XM4/w_n358_n132787# XM4/a_n100_n20699# -0.004445f
C1179 XM3/a_n158_38450# m1_1634_n2388# 6.1e-20
C1180 XM1/a_100_25966# XM3/a_n100_76685# 2.85e-20
C1181 XM2/a_100_n242394# XM3/a_n158_n36142# 0.077916f
C1182 XM1/a_100_109254# XM2/a_n158_n44694# 0.116862f
C1183 XM4/a_100_85070# m1_1634_n2388# 6.1e-20
C1184 XM2/a_100_n284570# XM3/a_n100_n77679# 0.005074f
C1185 XM4/a_100_4262# m1_1634_n2388# 6.1e-20
C1186 XM1/a_n100_4329# XM3/a_n158_55026# 2.85e-20
C1187 XM2/a_n158_n126410# XM3/a_n158_77818# 4.64e-21
C1188 XM1/a_n100_17253# XM3/a_n158_68494# 1.73e-20
C1189 XM1/a_n158_n50142# XM2/a_n158_n205490# 4.64e-21
C1190 XM4/w_n358_n132787# XM4/a_n100_11417# -0.004445f
C1191 XM2/a_100_n102686# XM3/a_n100_101549# 0.005074f
C1192 XM2/a_n158_n102686# XM3/a_n158_101646# 4.64e-21
C1193 XM1/a_n100_n123475# XM4/w_n358_n132787# 0.01363f
C1194 XM3/a_n100_n95291# m1_1634_n2388# 0.072015f
C1195 XM1/a_100_n103274# XM2/a_100_n258210# 4.64e-21
C1196 XM1/a_100_n18550# XM2/a_100_n171222# 4.64e-21
C1197 XM1/a_n158_104946# XM2/a_n100_n50063# 7.26e-20
C1198 XM1/a_n158_173874# XM2/a_n158_18570# 4.64e-21
C1199 XM1/a_n100_53153# XM3/a_n100_105693# 7.02e-19
C1200 XM1/a_100_34582# XM2/a_100_n118502# 4.64e-21
C1201 XM2/a_100_n92142# m1_1634_n2388# 0.023368f
C1202 XM1/a_n100_147929# XM2/a_n158_n5154# 0.005074f
C1203 XM2/a_n100_n134415# XM4/a_100_72638# 2.56e-20
C1204 XM1/a_100_n182254# XM4/w_n358_n132787# 0.054609f
C1205 XM1/a_n100_n117731# XM3/a_n100_n65247# 0.001093f
C1206 XM1/a_n158_n111890# XM3/a_n100_n60067# 1.94e-20
C1207 XM4/w_n358_n132787# XM2/a_n158_n160678# 0.102342f
C1208 XM2/a_n158_n279298# m1_1634_n2388# 2.36e-21
C1209 XM2/a_n100_n321571# XM4/a_100_n116950# 2.56e-20
C1210 XM2/a_100_n316202# XM3/a_n158_n111770# 0.042085f
C1211 XM1/a_n158_n137738# XM3/a_n100_n85967# 1.94e-20
C1212 XM4/w_n358_n132787# XM4/a_n100_n60067# -0.004445f
C1213 XM1/a_n158_67610# XM3/a_n100_118125# 1.94e-20
C1214 XM1/a_n100_61769# XM3/a_n158_114078# 2.85e-20
C1215 XM3/a_n158_n30962# m1_1634_n2388# 6.1e-20
C1216 XM1/a_n100_n17211# XM3/a_n100_33173# 2.08e-19
C1217 XM4/w_n358_n132787# XM3/a_n158_129618# 0.032295f
C1218 XM1/a_n100_30177# XM2/a_100_n123774# 1.45e-19
C1219 XM4/a_100_45702# m1_1634_n2388# 6.1e-20
C1220 XM2/a_n100_n63243# XM4/w_n358_n132787# 0.011583f
C1221 XM2/a_100_n86870# XM3/a_n158_120294# 0.003528f
C1222 XM1/a_n158_20222# XM2/a_n158_n134318# 9.28e-21
C1223 XM1/a_n100_n94755# m1_1634_n2388# 9.31e-20
C1224 XM2/a_100_n223942# XM3/a_n158_n18530# 0.077916f
C1225 XM2/a_100_n266118# XM3/a_n100_n60067# 0.010147f
C1226 XM4/a_n100_108801# m1_1634_n2388# 0.072015f
C1227 XM2/a_n100_n263579# XM3/a_n158_n58934# 0.005074f
C1228 XM4/w_n358_n132787# XM3/a_n100_n40383# 0.010958f
C1229 XM4/a_100_n25782# m1_1634_n2388# 6.1e-20
C1230 XM3/a_n100_36281# XM4/a_n100_36281# 0.009521f
C1231 XM1/a_100_94894# XM2/a_100_n60510# 4.64e-21
C1232 XM1/a_n158_n41526# XM2/a_n158_n194946# 4.64e-21
C1233 XM4/w_n358_n132787# XM2/a_100_n97414# 0.104171f
C1234 XM2/a_100_n216034# m1_1634_n2388# 0.017213f
C1235 XM4/w_n358_n132787# XM3/a_n100_48713# 0.008991f
C1236 XM1/a_n100_132133# XM2/a_100_n23606# 7.26e-20
C1237 XM4/w_n358_n132787# XM4/a_n100_n99435# -0.004445f
C1238 XM3/a_n158_n70330# m1_1634_n2388# 6.1e-20
C1239 XM1/a_n100_47409# XM4/w_n358_n132787# 0.01363f
C1240 XM1/a_n100_18689# XM2/a_100_n134318# 7.26e-20
C1241 XM1/a_100_n28602# XM2/a_n100_n181863# 0.005074f
C1242 XM1/a_n158_47506# XM3/a_n100_98441# 9.22e-21
C1243 XM1/a_n100_n182351# XM2/a_n158_n334654# 0.005074f
C1244 XM4/w_n358_n132787# XM2/a_n158_n284570# 0.107093f
C1245 XM2/a_n158_n260846# XM3/a_n158_n53754# 4.64e-21
C1246 XM1/a_100_n57322# m1_1634_n2388# 3.95e-19
C1247 XM1/a_n158_155206# XM2/a_n158_118# 4.64e-21
C1248 XM1/a_100_81970# XM2/a_n158_n71054# 0.060779f
C1249 XM1/a_100_15914# XM2/a_100_n136954# 4.64e-21
C1250 XM1/a_n158_53250# XM2/a_n158_n100050# 4.64e-21
C1251 XM1/a_n100_10073# XM2/a_n158_n144862# 0.005074f
C1252 XM1/a_n100_119209# XM2/a_n158_n34150# 0.005074f
C1253 XM2/a_n100_n189771# XM3/a_n100_16597# 0.003522f
C1254 XM1/a_100_123614# XM2/a_n100_n28975# 0.005074f
C1255 XM1/a_100_116434# XM2/a_n158_n39422# 0.014044f
C1256 XM1/a_n158_119306# XM2/a_n100_n34247# 7.26e-20
C1257 XM1/a_100_36018# XM3/a_n100_88081# 2.85e-20
C1258 XM4/a_n100_69433# m1_1634_n2388# 0.072015f
C1259 XM2/a_n158_n142226# XM3/a_n158_64350# 4.64e-21
C1260 XM1/a_n100_n99063# XM4/w_n358_n132787# 0.013401f
C1261 XM4/w_n358_n132787# XM3/a_n100_n79751# 0.009186f
C1262 XM4/a_100_n65150# m1_1634_n2388# 6.1e-20
C1263 XM2/a_100_n208126# XM3/a_n158_n1954# 0.077916f
C1264 XM1/a_n158_n57322# XM3/a_n100_n5159# 1.94e-20
C1265 XM3/a_n100_87045# m1_1634_n2388# 0.072015f
C1266 XM1/a_n158_31710# XM3/a_n100_83937# 1.94e-20
C1267 XM3/a_n158_n109698# m1_1634_n2388# 6.1e-20
C1268 XM1/a_100_n75990# XM3/a_n100_n23807# 2.85e-20
C1269 XM1/a_n100_n50239# XM3/a_n100_1057# 1.3e-20
C1270 XM2/a_n100_n189771# XM4/a_100_14622# 2.56e-20
C1271 XM1/a_n158_n12806# XM2/a_n100_n168683# 7.26e-20
C1272 XM1/a_n158_n2754# XM2/a_n100_n158139# 7.26e-20
C1273 XM1/a_100_n159278# XM3/a_n100_n107723# 2.85e-20
C1274 XM2/a_n100_n210859# XM4/a_100_n6098# 2.56e-20
C1275 XM1/a_n158_n15678# XM3/a_n100_35245# 5.01e-21
C1276 XM2/a_n100_n155503# m1_1634_n2388# 0.001109f
C1277 XM2/a_100_n247666# XM3/a_n100_n42455# 0.010147f
C1278 XM1/a_n100_54589# XM3/a_n100_105693# 6.5e-21
C1279 XM1/a_n100_n170863# XM4/w_n358_n132787# 0.01363f
C1280 XM3/a_n100_32137# m1_1634_n2388# 0.072015f
C1281 XM4/w_n358_n132787# XM2/a_100_n221306# 0.103826f
C1282 XM1/a_100_84842# XM4/w_n358_n132787# 0.053546f
C1283 XM1/a_100_n91786# XM4/w_n358_n132787# 0.054831f
C1284 XM1/a_100_171002# XM4/w_n358_n132787# 0.053546f
C1285 XM3/a_n100_131593# m1_1634_n2388# 0.036019f
C1286 XM1/a_n158_n182254# XM3/a_n100_n130515# 1.94e-20
C1287 XM1/a_100_n152098# XM3/a_n100_n100471# 2.85e-20
C1288 XM4/w_n358_n132787# XM3/a_n158_n15422# 0.032295f
C1289 XM4/a_n100_n2051# m1_1634_n2388# 0.072015f
C1290 XM1/a_100_113562# XM2/a_n158_n42058# 0.037022f
C1291 XM4/w_n358_n132787# XM3/a_n158_73674# 0.032295f
C1292 XM1/a_100_n131994# XM2/a_100_n287206# 4.64e-21
C1293 XM1/a_100_176746# XM2/a_n158_23842# 0.049095f
C1294 XM1/a_n100_107721# XM2/a_n158_n47330# 0.005074f
C1295 XM1/a_n100_n139271# XM2/a_100_n295114# 7.26e-20
C1296 XM4/w_n358_n132787# XM1/a_n100_n130655# 0.01363f
C1297 XM4/w_n358_n132787# XM3/a_n158_18766# 0.032295f
C1298 XM4/a_n100_30065# m1_1634_n2388# 0.072014f
C1299 XM4/w_n358_n132787# XM3/a_n100_n119119# 0.008893f
C1300 XM4/a_100_n104518# m1_1634_n2388# 6.1e-20
C1301 XM2/a_n158_n284570# XM3/a_n100_n77679# 7.26e-20
C1302 XM2/a_n100_n126507# XM3/a_n158_77818# 0.005074f
C1303 XM1/a_n158_n50142# XM2/a_n100_n205587# 7.26e-20
C1304 XM1/a_100_173874# XM2/a_100_18570# 4.64e-21
C1305 XM2/a_n158_n102686# XM3/a_n100_101549# 7.26e-20
C1306 XM2/a_n100_n102783# XM3/a_n158_101646# 0.005074f
C1307 XM1/a_n100_n182351# XM3/a_n158_n130418# 2.85e-20
C1308 XM1/a_n158_n110454# XM3/a_n100_n59031# 3.55e-20
C1309 XM1/a_n158_15914# XM3/a_n100_67361# 3.07e-20
C1310 XM1/a_n100_11509# XM3/a_n158_63314# 2.85e-20
C1311 XM1/a_100_n137738# XM3/a_n100_n85967# 2.85e-20
C1312 XM1/a_100_n120506# XM3/a_n158_n69294# 0.001549f
C1313 XM1/a_100_n103274# XM2/a_n158_n258210# 0.10362f
C1314 XM1/a_100_n18550# XM2/a_n158_n171222# 0.026507f
C1315 XM2/a_n100_n168683# XM3/a_n158_35342# 0.001535f
C1316 XM1/a_n100_n2851# XM3/a_n158_47774# 2.85e-20
C1317 XM1/a_n100_1457# XM3/a_n100_51821# 4.68e-19
C1318 XM4/w_n358_n132787# XM4/a_n100_124341# -0.004445f
C1319 XM1/a_100_34582# XM2/a_n158_n118502# 0.066621f
C1320 XM1/a_100_n110454# XM2/a_100_n266118# 4.64e-21
C1321 XM1/a_n158_n78862# XM2/a_n158_n231850# 4.64e-21
C1322 XM1/a_n100_156545# XM2/a_n158_2754# 0.010147f
C1323 XM4/w_n358_n132787# XM2/a_n100_n160775# 0.024756f
C1324 XM2/a_n100_n279395# m1_1634_n2388# 0.002028f
C1325 XM4/w_n358_n132787# XM3/a_n158_n54790# 0.032295f
C1326 XM4/a_n100_n41419# m1_1634_n2388# 0.072015f
C1327 XM2/a_n158_n316202# XM3/a_n158_n111770# 4.64e-21
C1328 XM1/a_n100_n100499# XM2/a_100_n252938# 7.26e-20
C1329 XM2/a_100_n229214# XM3/a_n100_n24843# 0.005074f
C1330 XM4/w_n358_n132787# XM3/a_n100_129521# 0.009186f
C1331 XM1/a_n100_30177# XM2/a_n158_n123774# 0.010147f
C1332 XM3/a_n158_57098# m1_1634_n2388# 6.1e-20
C1333 XM1/a_100_n154970# XM3/a_n100_n104615# 5.9e-19
C1334 XM1/a_100_n179382# XM3/a_n100_n127407# 7.52e-19
C1335 XM2/a_n100_n318935# XM4/a_100_n111770# 2.56e-20
C1336 XM2/a_100_n313566# XM3/a_n158_n106590# 0.021833f
C1337 XM1/a_100_175310# XM4/w_n358_n132787# 0.048442f
C1338 XM3/a_n100_89117# XM4/a_n100_89117# 0.009521f
C1339 XM2/a_n158_n86870# XM3/a_n158_120294# 4.64e-21
C1340 XM2/a_100_n86870# XM3/a_n100_120197# 0.005074f
C1341 XM2/a_n100_n79059# XM4/a_100_125474# 2.56e-20
C1342 XM4/w_n358_n132787# XM4/a_n100_84973# -0.004445f
C1343 XM1/a_n100_n114859# m1_1634_n2388# 1.21e-19
C1344 XM4/w_n358_n132787# XM4/a_n100_4165# -0.004445f
C1345 XM1/a_100_n117634# XM2/a_n158_n271390# 0.116862f
C1346 XM2/a_n158_n266118# XM3/a_n100_n60067# 1.45e-19
C1347 XM3/a_n100_n21735# m1_1634_n2388# 0.072014f
C1348 XM1/a_100_23094# XM4/w_n358_n132787# 0.048442f
C1349 XM4/w_n358_n132787# XM3/a_n158_n94158# 0.032295f
C1350 XM4/a_n100_n80787# m1_1634_n2388# 0.072015f
C1351 XM1/a_n158_n41526# XM2/a_n100_n195043# 7.26e-20
C1352 XM4/w_n358_n132787# XM2/a_n158_n97414# 0.101988f
C1353 XM1/a_n100_146493# XM4/w_n358_n132787# 0.012279f
C1354 XM1/a_100_168130# XM2/a_100_13298# 4.64e-21
C1355 XM1/a_n100_18689# XM2/a_n158_n134318# 0.005074f
C1356 XM1/a_100_73354# XM2/a_100_n81598# 4.64e-21
C1357 XM4/w_n358_n132787# XM2/a_n100_n284667# 0.025032f
C1358 XM2/a_n100_n260943# XM3/a_n158_n53754# 0.005074f
C1359 XM2/a_n100_n15795# XM4/w_n358_n132787# 0.013155f
C1360 XM3/a_n158_107862# m1_1634_n2388# 6.1e-20
C1361 XM1/a_n158_n173638# XM2/a_n158_n329382# 4.64e-21
C1362 XM1/a_100_n139174# XM3/a_n100_n87003# 2.85e-20
C1363 XM1/a_n100_90489# XM4/w_n358_n132787# 0.012279f
C1364 XM1/a_100_15914# XM2/a_n158_n136954# 0.04559f
C1365 XM1/a_100_n116198# XM4/w_n358_n132787# 0.054694f
C1366 XM1/a_100_166694# XM2/a_n100_10565# 0.004433f
C1367 XM4/a_100_119258# m1_1634_n2388# 6.1e-20
C1368 XM2/a_100_n144862# XM3/a_n100_59073# 0.005074f
C1369 XM1/a_100_n176510# XM3/a_n158_n125238# 0.00544f
C1370 XM1/a_n100_n35879# XM3/a_n158_16694# 6.97e-21
C1371 XM1/a_n158_n19986# XM3/a_n100_31101# 1.94e-20
C1372 XM1/a_n158_53250# XM2/a_n100_n100147# 7.26e-20
C1373 XM1/a_n158_n44398# XM3/a_n100_6237# 2.6e-21
C1374 XM4/w_n358_n132787# XM4/a_n100_45605# -0.004445f
C1375 XM1/a_n100_5765# XM2/a_100_n150134# 7.26e-20
C1376 XM1/a_100_n63066# m1_1634_n2388# 5.46e-19
C1377 XM1/a_100_69046# XM2/a_100_n86870# 4.64e-21
C1378 XM3/a_n100_n61103# m1_1634_n2388# 0.072015f
C1379 XM1/a_n158_n71682# XM2/a_n158_n226578# 4.64e-21
C1380 XM2/a_n100_n142323# XM3/a_n158_64350# 0.005074f
C1381 XM1/a_100_n8498# XM2/a_100_n163314# 4.64e-21
C1382 XM4/a_n100_n120155# m1_1634_n2388# 0.072015f
C1383 XM2/a_100_n295114# XM3/a_n158_n88978# 0.077916f
C1384 XM3/a_n100_n12411# XM4/a_n100_n12411# 0.009521f
C1385 XM2/a_100_n337290# XM3/a_n100_n130515# 0.005074f
C1386 XM1/a_100_n136302# XM3/a_n100_n85967# 1.31e-19
C1387 XM1/a_n100_n33007# XM4/w_n358_n132787# 0.013564f
C1388 XM2/a_100_n152770# m1_1634_n2388# 0.017213f
C1389 XM4/w_n358_n132787# XM3/a_n100_67361# 0.009055f
C1390 XM2/a_n158_n247666# XM3/a_n100_n42455# 1.45e-19
C1391 XM4/w_n358_n132787# XM4/a_n100_n25879# -0.004445f
C1392 XM1/a_n158_n73118# XM3/a_n100_n21735# 3.89e-20
C1393 XM1/a_100_34582# XM3/a_n158_86106# 0.003892f
C1394 XM4/w_n358_n132787# XM2/a_n158_n221306# 0.107093f
C1395 XM2/a_n100_26381# XM1/a_100_182490# 0.004836f
C1396 XM2/a_100_26478# XM1/a_n100_182393# 6.36e-20
C1397 XM1/a_100_41762# XM2/a_100_n113230# 4.64e-21
C1398 XM4/w_n358_n132787# XM3/a_n100_12453# 0.008963f
C1399 XM4/a_100_79890# m1_1634_n2388# 6.1e-20
C1400 XM1/a_n158_n91786# XM2/a_n158_n245030# 4.64e-21
C1401 XM1/a_n158_n34346# XM2/a_n158_n187038# 4.64e-21
C1402 XM2/a_n100_n187135# XM4/a_100_19802# 2.56e-20
C1403 XM1/a_n158_41762# XM2/a_n100_n110691# 4.26e-20
C1404 sw_b XM4/w_n358_n132787# 0.006002f
C1405 XM1/a_n158_n163586# XM2/a_n158_n318838# 4.64e-21
C1406 XM2/a_100_n131682# XM3/a_n100_73577# 0.010147f
C1407 XM3/a_n158_8406# m1_1634_n2388# 6.1e-20
C1408 XM4/w_n358_n132787# XM3/a_n158_105790# 0.032295f
C1409 XM1/a_100_n131994# XM2/a_n158_n287206# 0.076747f
C1410 XM3/a_n100_n100471# m1_1634_n2388# 0.072015f
C1411 XM3/a_n100_124341# XM4/a_n100_124341# 0.009521f
C1412 XM1/a_n100_n139271# XM2/a_n158_n295114# 0.005074f
C1413 XM2/a_100_n173858# XM3/a_n100_31101# 0.010147f
C1414 XM1/a_n100_n12903# XM3/a_n100_38353# 5.33e-19
C1415 XM1/a_n100_110593# XM2/a_100_n42058# 7.26e-20
C1416 XM1/a_n158_100638# XM2/a_n100_n55335# 7.26e-20
C1417 XM3/a_n100_n32095# XM4/a_n100_n32095# 0.009521f
C1418 XM2/a_100_n102686# XM3/a_n158_102682# 0.077916f
C1419 XM1/a_100_n103274# XM2/a_n100_n258307# 0.005074f
C1420 XM4/w_n358_n132787# XM3/a_n100_n6195# 0.008086f
C1421 XM1/a_n158_53250# XM3/a_n100_104657# 2e-20
C1422 XM1/a_100_n18550# XM2/a_n100_n171319# 0.005074f
C1423 XM1/a_n100_5765# XM3/a_n158_58134# 2.85e-20
C1424 XM1/a_n100_n133527# XM3/a_n158_n82762# 2.85e-20
C1425 XM1/a_100_34582# XM2/a_n100_n118599# 0.005074f
C1426 XM1/a_n158_n121942# XM2/a_n158_n276662# 9.28e-21
C1427 XM4/w_n358_n132787# XM4/a_n100_n65247# -0.004445f
C1428 XM1/a_100_n110454# XM2/a_n158_n266118# 0.032738f
C1429 XM1/a_100_n87478# XM3/a_n100_n37275# 1.99e-22
C1430 XM1/a_n158_n78862# XM2/a_n100_n231947# 7.26e-20
C1431 XM2/a_n100_n73787# XM3/a_n158_130654# 0.005074f
C1432 XM2/a_n100_n92239# m1_1634_n2388# 0.001602f
C1433 XM2/a_100_n276662# XM3/a_n158_n71366# 0.077916f
C1434 XM3/a_n158_n36142# m1_1634_n2388# 6.1e-20
C1435 XM4/a_100_40522# m1_1634_n2388# 6.1e-20
C1436 XM3/a_n100_50785# m1_1634_n2388# 0.072015f
C1437 XM4/w_n358_n132787# XM2/a_100_n158042# 0.103342f
C1438 XM2/a_100_n318838# XM3/a_n100_n112903# 0.010147f
C1439 XM2/a_100_n276662# m1_1634_n2388# 0.019664f
C1440 XM1/a_n100_n10031# XM3/a_n100_42497# 8.59e-19
C1441 XM1/a_100_4426# XM3/a_n100_55965# 2.85e-20
C1442 XM3/a_n100_57001# XM4/a_n100_57001# 0.009521f
C1443 XM2/a_n100_n316299# XM3/a_n158_n111770# 0.005074f
C1444 XM1/a_n100_n100499# XM2/a_n158_n252938# 0.005074f
C1445 XM1/a_n100_n78959# XM4/w_n358_n132787# 0.01363f
C1446 XM1/a_100_58994# XM3/a_n100_109837# 2.85e-20
C1447 XM4/w_n358_n132787# XM3/a_n158_92322# 0.032295f
C1448 XM2/a_100_n118502# XM3/a_n100_88081# 0.005074f
C1449 XM2/a_n158_n229214# XM3/a_n100_n24843# 7.26e-20
C1450 XM1/a_100_n31474# XM3/a_n158_19802# 0.00544f
C1451 XM1/a_100_97766# XM2/a_n100_n57971# 0.005074f
C1452 XM4/w_n358_n132787# XM3/a_n158_37414# 0.032295f
C1453 XM2/a_100_n160678# XM3/a_n100_45605# 0.005482f
C1454 XM3/a_n100_n51779# XM4/a_n100_n51779# 0.009521f
C1455 XM1/a_100_25966# XM2/a_n100_n126507# 0.004594f
C1456 XM2/a_n158_n313566# XM3/a_n158_n106590# 4.64e-21
C1457 XM1/a_100_n38654# XM3/a_n100_12453# 3.05e-20
C1458 XM4/a_n100_103621# m1_1634_n2388# 0.072015f
C1459 XM1/a_n158_n123378# XM2/a_n158_n279298# 4.64e-21
C1460 XM2/a_100_n226578# XM3/a_n100_n19663# 0.005074f
C1461 XM2/a_n158_n86870# XM3/a_n100_120197# 7.26e-20
C1462 XM2/a_n100_n86967# XM3/a_n158_120294# 0.005074f
C1463 XM4/w_n358_n132787# XM3/a_n100_n45563# 0.008913f
C1464 XM4/a_100_n30962# m1_1634_n2388# 6.1e-20
C1465 XM4/w_n358_n132787# XM4/a_n100_n104615# -0.004445f
C1466 XM1/a_100_n28602# m1_1634_n2388# 0.001516f
C1467 XM3/a_n158_n75510# m1_1634_n2388# 6.1e-20
C1468 XM3/a_n100_107765# XM4/a_n100_107765# 0.009521f
C1469 XM2/a_n100_n76423# XM4/a_100_130654# 2.56e-20
C1470 XM4/w_n358_n132787# XM2/a_n100_n97511# 0.025292f
C1471 XM1/a_100_18786# XM2/a_100_n136954# 4.64e-21
C1472 XM1/a_n100_n96191# XM4/w_n358_n132787# 0.013525f
C1473 XM2/a_n100_n216131# m1_1634_n2388# 0.002821f
C1474 XM1/a_100_54686# XM2/a_n158_n100050# 0.116862f
C1475 XM1/a_100_n42962# XM3/a_n100_8309# 5.71e-20
C1476 XM1/a_n100_n11467# m1_1634_n2388# 1.3e-19
C1477 XM1/a_100_73354# XM2/a_n158_n81598# 0.102062f
C1478 XM4/w_n358_n132787# XM2/a_100_n281934# 0.103342f
C1479 XM2/a_100_n258210# XM3/a_n158_n53754# 0.044422f
C1480 XM3/a_n158_75746# m1_1634_n2388# 6.1e-20
C1481 XM1/a_n100_14381# XM2/a_100_n139590# 1.45e-19
C1482 XM2/a_n100_n263579# XM4/a_100_n58934# 2.56e-20
C1483 XM3/a_n100_107765# m1_1634_n2388# 0.072015f
C1484 XM1/a_n158_n173638# XM2/a_n100_n329479# 7.26e-20
C1485 XM2/a_100_n300386# XM3/a_n100_n95291# 0.010147f
C1486 XM3/a_n100_n71463# XM4/a_n100_n71463# 0.009521f
C1487 XM1/a_100_15914# XM2/a_n100_n137051# 0.005074f
C1488 XM4/a_n100_64253# m1_1634_n2388# 0.072015f
C1489 XM2/a_n158_n144862# XM3/a_n100_59073# 7.26e-20
C1490 XM1/a_100_n144918# XM3/a_n158_n93122# 0.003891f
C1491 XM1/a_n100_10073# XM2/a_100_n142226# 6.96e-20
C1492 XM4/w_n358_n132787# XM3/a_n100_n84931# 0.009186f
C1493 XM4/a_100_n70330# m1_1634_n2388# 6.1e-20
C1494 XM3/a_n158_20838# m1_1634_n2388# 6.1e-20
C1495 XM1/a_100_126486# XM2/a_100_n26242# 4.64e-21
C1496 XM1/a_n158_48942# XM2/a_n158_n105322# 9.28e-21
C1497 XM1/a_100_34582# m1_1634_n2388# 0.001152f
C1498 XM1/a_n100_5765# XM2/a_n158_n150134# 0.005074f
C1499 XM1/a_100_n55886# XM3/a_n158_n4026# 0.001549f
C1500 XM1/a_100_69046# XM2/a_n158_n86870# 0.008202f
C1501 XM1/a_100_46070# XM3/a_n100_97405# 5.71e-20
C1502 XM3/a_n158_n114878# m1_1634_n2388# 6.1e-20
C1503 XM1/a_n100_n78959# XM2/a_100_n234486# 7.26e-20
C1504 XM1/a_n158_n71682# XM2/a_n100_n226675# 7.18e-20
C1505 XM1/a_100_n8498# XM2/a_n158_n163314# 0.115304f
C1506 XM1/a_n100_41665# XM3/a_n100_93261# 6.79e-19
C1507 XM2/a_n158_n337290# XM3/a_n100_n130515# 7.26e-20
C1508 XM1/a_n158_54686# XM2/a_n158_n100050# 9.28e-21
C1509 XM1/a_n158_n124814# XM3/a_n100_n73535# 3.89e-20
C1510 XM4/w_n358_n132787# XM3/a_n158_n20602# 0.032295f
C1511 XM4/a_n100_n7231# m1_1634_n2388# 0.072015f
C1512 XM1/a_n158_n12806# XM2/a_n158_n165950# 4.64e-21
C1513 XM1/a_n158_n2754# XM2/a_n158_n155406# 4.64e-21
C1514 XM1/a_100_148026# XM2/a_100_n7790# 4.64e-21
C1515 XM1/a_n100_54589# XM3/a_n158_106826# 8.85e-19
C1516 XM3/a_n100_n91147# XM4/a_n100_n91147# 0.009521f
C1517 XM4/w_n358_n132787# XM2/a_n100_n221403# 0.025855f
C1518 XM1/a_100_n47270# XM3/a_n100_3129# 2.85e-20
C1519 XM1/a_100_41762# XM2/a_n158_n113230# 0.098168f
C1520 XM1/a_100_37454# XM4/w_n358_n132787# 0.054609f
C1521 XM4/a_n100_24885# m1_1634_n2388# 0.072015f
C1522 XM2/a_n158_n10426# XM1/a_n158_145154# 4.64e-21
C1523 XM2/a_100_n10426# XM1/a_100_145154# 4.64e-21
C1524 XM1/a_n158_n91786# XM2/a_n100_n245127# 7.26e-20
C1525 XM1/a_100_n35782# XM3/a_n100_14525# 2.85e-20
C1526 XM1/a_n158_n34346# XM2/a_n100_n187135# 7.26e-20
C1527 XM4/w_n358_n132787# XM3/a_n100_n124299# 0.009186f
C1528 XM1/a_n158_n163586# XM2/a_n100_n318935# 7.26e-20
C1529 XM4/a_100_n109698# m1_1634_n2388# 6.1e-20
C1530 XM2/a_n158_n131682# XM3/a_n100_73577# 1.45e-19
C1531 XM1/a_n158_n160714# XM2/a_n158_n316202# 4.64e-21
C1532 XM4/w_n358_n132787# XM3/a_n100_105693# 0.009014f
C1533 XM1/a_100_n131994# XM2/a_n100_n287303# 0.005074f
C1534 XM1/a_100_155206# XM2/a_100_2754# 4.64e-21
C1535 XM2/a_n158_n15698# XM1/a_n100_137877# 0.00864f
C1536 XM2/a_n158_n173858# XM3/a_n100_31101# 1.45e-19
C1537 XM2/a_100_n281934# XM3/a_n100_n77679# 0.005074f
C1538 XM4/w_n358_n132787# XM4/a_n100_119161# -0.004445f
C1539 XM1/a_n100_n146451# XM3/a_n100_n95291# 6.76e-19
C1540 XM2/a_100_n126410# XM3/a_n158_78854# 0.077916f
C1541 XM1/a_n158_n50142# XM2/a_n158_n202854# 4.64e-21
C1542 XM1/a_100_110690# XM2/a_n158_n44694# 0.06f
C1543 XM2/a_100_n102686# XM3/a_n100_102585# 0.010147f
C1544 XM3/a_n100_24885# XM4/a_n100_24885# 0.009521f
C1545 XM1/a_100_10170# XM3/a_n100_61145# 2.85e-20
C1546 XM1/a_n100_n139271# XM3/a_n100_n88039# 8.46e-19
C1547 XM1/a_n158_n144918# XM3/a_n100_n94255# 1.94e-20
C1548 XM4/w_n358_n132787# XM3/a_n158_n59970# 0.032295f
C1549 XM4/a_n100_n46599# m1_1634_n2388# 0.072015f
C1550 XM2/a_100_n168586# XM3/a_n158_36378# 0.077916f
C1551 XM1/a_100_n110454# XM2/a_n100_n266215# 0.005074f
C1552 XM1/a_n158_176746# XM2/a_n158_23842# 4.64e-21
C1553 XM2/a_100_n89506# m1_1634_n2388# 0.017213f
C1554 XM4/w_n358_n132787# XM3/a_n100_86009# 0.008206f
C1555 XM3/a_n100_n110831# XM4/a_n100_n110831# 0.009521f
C1556 XM2/a_n100_n131779# XM4/a_100_72638# 2.56e-20
C1557 XM1/a_100_n81734# XM2/a_100_n237122# 4.64e-21
C1558 XM1/a_n158_2990# XM3/a_n100_54929# 1.94e-20
C1559 XM4/w_n358_n132787# XM2/a_n158_n158042# 0.107093f
C1560 XM2/a_n158_n318838# XM3/a_n100_n112903# 1.45e-19
C1561 XM4/w_n358_n132787# XM3/a_n100_31101# 0.008928f
C1562 XM1/a_n158_156642# XM2/a_n158_2754# 9.28e-21
C1563 XM1/a_n158_67610# XM3/a_n100_119161# 1.94e-20
C1564 XM2/a_n158_n118502# XM3/a_n100_88081# 7.26e-20
C1565 XM1/a_n158_n96094# XM3/a_n100_n44527# 1.94e-20
C1566 XM1/a_n158_n80298# XM3/a_n100_n27951# 1.06e-20
C1567 XM4/w_n358_n132787# XM3/a_n158_130654# 0.038462f
C1568 XM1/a_100_n15678# XM3/a_n100_35245# 0.001161f
C1569 XM1/a_100_160950# XM2/a_n158_5390# 0.042864f
C1570 XM4/w_n358_n132787# XM4/a_n100_79793# -0.004445f
C1571 XM1/a_n100_n50239# XM3/a_n158_2190# 2.85e-20
C1572 XM2/a_n158_n160678# XM3/a_n100_45605# 8.75e-20
C1573 XM2/a_n100_n313663# XM3/a_n158_n106590# 0.005074f
C1574 XM3/a_n100_n26915# m1_1634_n2388# 0.072015f
C1575 XM1/a_n100_91925# XM2/a_100_n63146# 7.26e-20
C1576 XM2/a_100_n113230# XM3/a_n158_93358# 0.059611f
C1577 XM1/a_n158_n123378# XM2/a_n100_n279395# 7.26e-20
C1578 XM2/a_n158_n226578# XM3/a_n100_n19663# 7.26e-20
C1579 XM2/a_100_n84234# XM3/a_n158_120294# 0.051432f
C1580 XM4/w_n358_n132787# XM3/a_n158_n99338# 0.032295f
C1581 XM4/a_n100_n85967# m1_1634_n2388# 0.072015f
C1582 XM2/a_100_n202854# XM3/a_n100_3129# 0.010147f
C1583 XM2/a_n158_n44694# XM4/w_n358_n132787# 0.107093f
C1584 XM1/a_n158_n74554# XM2/a_n158_n229214# 9.28e-21
C1585 XM1/a_n100_40229# m1_1634_n2388# 9.41e-20
C1586 XM1/a_100_n154970# XM2/a_100_n310930# 4.64e-21
C1587 XM1/a_n100_n50239# XM4/w_n358_n132787# 0.013468f
C1588 XM2/a_100_n155406# XM3/a_n158_50882# 0.077916f
C1589 XM1/a_n100_150801# XM4/w_n358_n132787# 0.011694f
C1590 XM3/a_n100_n130515# XM4/a_n100_n130515# 0.009521f
C1591 XM1/a_100_20222# XM2/a_n158_n134318# 0.116862f
C1592 XM1/a_n158_150898# XM2/a_n158_n2518# 4.64e-21
C1593 XM1/a_n158_n88914# XM2/a_n158_n242394# 4.64e-21
C1594 XM1/a_n100_n66035# m1_1634_n2388# 9.07e-20
C1595 XM3/a_n100_69433# m1_1634_n2388# 0.072015f
C1596 XM3/a_n100_8309# XM4/a_n100_8309# 0.009521f
C1597 XM1/a_n100_152237# XM2/a_n100_n2615# 0.001471f
C1598 XM1/a_n100_89053# XM4/w_n358_n132787# 0.011583f
C1599 XM4/w_n358_n132787# XM2/a_100_n94778# 0.103342f
C1600 XM1/a_100_18786# XM2/a_n158_n136954# 0.025338f
C1601 XM2/a_100_n213398# m1_1634_n2388# 0.022596f
C1602 XM4/a_100_114078# m1_1634_n2388# 6.1e-20
C1603 XM3/a_n100_14525# m1_1634_n2388# 0.072015f
C1604 XM1/a_100_73354# XM2/a_n100_n81695# 0.005074f
C1605 XM4/w_n358_n132787# XM2/a_n158_n281934# 0.107093f
C1606 XM2/a_n158_n258210# XM3/a_n158_n53754# 4.64e-21
C1607 XM4/w_n358_n132787# XM4/a_n100_40425# -0.004445f
C1608 XM1/a_n100_14381# XM2/a_n158_n139590# 0.010147f
C1609 XM2/a_n158_n300386# XM3/a_n100_n95291# 1.45e-19
C1610 XM1/a_n158_n140610# XM3/a_n100_n89075# 1.94e-20
C1611 XM3/a_n100_n66283# m1_1634_n2388# 0.072015f
C1612 XM1/a_n100_45973# XM4/w_n358_n132787# 0.013401f
C1613 XM4/w_n358_n132787# XM3/a_n158_56062# 0.032295f
C1614 XM1/a_n100_47409# XM2/a_100_n107958# 7.26e-20
C1615 XM1/a_n100_10073# XM2/a_n158_n142226# 0.004998f
C1616 XM4/a_n100_n125335# m1_1634_n2388# 0.072014f
C1617 XM2/a_100_n255574# XM3/a_n158_n48574# 0.019496f
C1618 XM1/a_100_n126250# XM4/w_n358_n132787# 0.055048f
C1619 XM2/a_n100_n260943# XM4/a_100_n53754# 2.56e-20
C1620 XM1/a_100_69046# XM2/a_n100_n86967# 0.005074f
C1621 XM1/a_n100_n162247# XM3/a_n100_n111867# 2.6e-19
C1622 XM1/a_n100_n78959# XM2/a_n158_n234486# 0.005074f
C1623 XM1/a_100_37454# XM3/a_n158_88178# 0.00544f
C1624 XM1/a_100_n8498# XM2/a_n100_n163411# 3.27e-19
C1625 XM1/a_100_84842# XM2/a_n100_n71151# 0.005074f
C1626 XM4/w_n358_n132787# XM4/a_n100_n31059# -0.004445f
C1627 XM1/a_100_n19986# XM2/a_n158_n173858# 0.116862f
C1628 XM1/a_n100_n14339# XM2/a_100_n168586# 1.45e-19
C1629 XM1/a_100_7298# XM4/w_n358_n132787# 0.048442f
C1630 XM4/a_100_74710# m1_1634_n2388# 6.1e-20
C1631 XM1/a_n158_n12806# XM2/a_n100_n166047# 7.26e-20
C1632 XM1/a_n158_n2754# XM2/a_n100_n155503# 7.26e-20
C1633 XM2/a_n100_n152867# m1_1634_n2388# 7.61e-19
C1634 XM3/a_n100_2093# m1_1634_n2388# 0.072015f
C1635 XM1/a_n100_n94755# XM3/a_n158_n42358# 2.85e-20
C1636 XM3/a_n100_n105651# m1_1634_n2388# 0.072015f
C1637 XM4/w_n358_n132787# XM2/a_100_n218670# 0.103791f
C1638 XM2/a_n158_n18334# XM1/a_100_136538# 0.109852f
C1639 XM2/a_n100_n18431# XM1/a_n158_136538# 5.78e-20
C1640 XM2/a_100_n18334# XM1/a_n100_135005# 7.26e-20
C1641 XM1/a_100_41762# XM2/a_n100_n113327# 0.005074f
C1642 XM3/a_n158_94394# m1_1634_n2388# 6.1e-20
C1643 XM2/a_100_n337290# m1_1634_n2388# 0.017213f
C1644 XM1/a_n100_n48803# m1_1634_n2388# 1.3e-19
C1645 XM2/a_100_n329382# XM3/a_n158_n124202# 0.077916f
C1646 XM3/a_n100_77721# XM4/a_n100_77721# 0.009521f
C1647 XM1/a_n158_27402# XM3/a_n100_79793# 1.8e-21
C1648 XM1/a_n158_n160714# XM2/a_n100_n316299# 7.26e-20
C1649 XM3/a_n158_39486# m1_1634_n2388# 6.1e-20
C1650 XM4/w_n358_n132787# XM1/a_100_132230# 0.053546f
C1651 XM1/a_100_n131994# XM2/a_100_n284570# 4.64e-21
C1652 XM1/a_100_n19986# XM4/w_n358_n132787# 0.048442f
C1653 XM1/a_100_25966# XM3/a_n100_77721# 2.85e-20
C1654 XM4/w_n358_n132787# XM3/a_n100_n11375# 0.009836f
C1655 XM1/a_n100_n165119# m1_1634_n2388# 7.81e-20
C1656 XM1/a_n100_n139271# XM2/a_100_n292478# 7.26e-20
C1657 XM2/a_n158_n281934# XM3/a_n100_n77679# 7.26e-20
C1658 XM1/a_n158_160950# XM2/a_n158_5390# 4.64e-21
C1659 XM4/w_n358_n132787# XM4/a_n100_n70427# -0.004445f
C1660 XM1/a_n100_4329# XM3/a_n158_56062# 1.14e-20
C1661 XM1/a_n158_23094# XM3/a_n100_73577# 1.94e-20
C1662 XM1/a_n100_17253# XM3/a_n158_69530# 2.85e-20
C1663 XM3/a_n158_n41322# m1_1634_n2388# 6.1e-20
C1664 XM1/a_n158_n50142# XM2/a_n100_n202951# 7.26e-20
C1665 XM2/a_n158_n102686# XM3/a_n100_102585# 1.45e-19
C1666 XM4/a_100_35342# m1_1634_n2388# 6.1e-20
C1667 XM2/a_100_n237122# XM3/a_n158_n30962# 0.077916f
C1668 XM1/a_n100_n41623# XM2/a_100_n197582# 3.46e-20
C1669 XM2/a_100_n73690# XM4/a_n100_131593# 2.76e-19
C1670 XM2/a_100_n279298# XM3/a_n100_n72499# 0.005074f
C1671 XM1/a_n158_173874# XM2/a_n158_21206# 4.64e-21
C1672 XM1/a_100_n110454# XM2/a_100_n263482# 4.64e-21
C1673 XM1/a_100_n9934# XM3/a_n100_40425# 0.001413f
C1674 XM1/a_100_2990# XM3/a_n100_53893# 2.85e-20
C1675 XM1/a_100_n81734# XM2/a_n158_n237122# 0.059611f
C1676 XM1/a_100_n162150# XM3/a_n100_n110831# 5.71e-20
C1677 XM1/a_n100_n70343# m1_1634_n2388# 1.29e-19
C1678 XM4/w_n358_n132787# XM2/a_n100_n158139# 0.024482f
C1679 XM2/a_n100_n276759# m1_1634_n2388# 0.003031f
C1680 XM4/a_n100_98441# m1_1634_n2388# 0.072015f
C1681 XM4/w_n358_n132787# XM3/a_n100_n50743# 0.008928f
C1682 XM4/a_100_n36142# m1_1634_n2388# 6.1e-20
C1683 XM1/a_100_103510# XM2/a_n158_n49966# 0.104789f
C1684 XM4/w_n358_n132787# XM3/a_n100_130557# 0.009017f
C1685 XM2/a_n100_n129143# XM4/a_100_77818# 2.56e-20
C1686 XM2/a_n100_n60607# XM4/w_n358_n132787# 0.012279f
C1687 XM4/w_n358_n132787# XM4/a_n100_n109795# -0.004445f
C1688 XM1/a_100_n101838# XM3/a_n100_n49707# 2.85e-20
C1689 XM1/a_100_n64502# XM2/a_n158_n218670# 0.116862f
C1690 XM1/a_n158_n58758# XM3/a_n100_n8267# 1.94e-20
C1691 XM2/a_n100_n160775# XM3/a_n100_45605# 0.004501f
C1692 XM2/a_100_n310930# XM3/a_n158_n106590# 0.033127f
C1693 XM3/a_n158_n80690# m1_1634_n2388# 6.1e-20
C1694 XM2/a_n100_n316299# XM4/a_100_n111770# 2.56e-20
C1695 XM2/a_n158_n113230# XM3/a_n158_93358# 4.64e-21
C1696 XM1/a_n158_130794# XM2/a_n158_n23606# 9.28e-21
C1697 XM2/a_100_n84234# XM3/a_n100_120197# 0.005074f
C1698 XM2/a_n158_n84234# XM3/a_n158_120294# 4.64e-21
C1699 XM2/a_n158_n202854# XM3/a_n100_3129# 1.45e-19
C1700 XM1/a_n100_71821# XM4/w_n358_n132787# 0.013852f
C1701 XM1/a_100_n154970# XM2/a_n158_n310930# 0.003918f
C1702 XM1/a_n158_n121942# XM3/a_n100_n71463# 1.94e-20
C1703 XM1/a_100_n65938# XM4/w_n358_n132787# 0.054609f
C1704 XM1/a_100_160950# XM4/w_n358_n132787# 0.053546f
C1705 XM1/a_100_n150662# XM4/w_n358_n132787# 0.053768f
C1706 XM1/a_n158_n88914# XM2/a_n100_n242491# 7.26e-20
C1707 XM1/a_100_94894# XM2/a_100_n57874# 4.64e-21
C1708 XM1/a_n100_n167991# XM3/a_n158_n116950# 8.48e-19
C1709 XM2/a_100_n218670# XM3/a_n158_n13350# 0.077916f
C1710 XM1/a_n100_132133# XM2/a_100_n20970# 7.26e-20
C1711 XM1/a_100_123614# XM4/w_n358_n132787# 0.053546f
C1712 XM4/w_n358_n132787# XM2/a_n158_n94778# 0.10594f
C1713 XM1/a_100_18786# XM2/a_n100_n137051# 0.005074f
C1714 XM1/a_n100_17253# XM4/w_n358_n132787# 0.0135f
C1715 XM2/a_n158_n213398# m1_1634_n2388# 2.36e-21
C1716 XM4/w_n358_n132787# XM3/a_n100_49749# 0.009036f
C1717 XM4/a_n100_59073# m1_1634_n2388# 0.072015f
C1718 XM2/a_100_n260846# XM3/a_n100_n54887# 0.010147f
C1719 XM1/a_n100_127825# XM2/a_100_n26242# 1.45e-19
C1720 XM4/w_n358_n132787# XM3/a_n100_n90111# 0.009186f
C1721 XM4/a_100_n75510# m1_1634_n2388# 6.1e-20
C1722 XM1/a_n158_47506# XM3/a_n100_99477# 1.92e-20
C1723 XM4/w_n358_n132787# XM2/a_n100_n282031# 0.024576f
C1724 XM2/a_n100_n258307# XM3/a_n158_n53754# 0.005074f
C1725 XM3/a_n158_108898# m1_1634_n2388# 6.1e-20
C1726 XM1/a_n158_n173638# XM2/a_n158_n326746# 4.64e-21
C1727 XM3/a_n158_n120058# m1_1634_n2388# 6.1e-20
C1728 XM1/a_100_n21422# XM3/a_n158_30162# 0.00544f
C1729 XM1/a_n158_44634# XM3/a_n100_95333# 1.94e-20
C1730 XM1/a_n100_38793# XM3/a_n158_91286# 0.001486f
C1731 XM1/a_n100_80437# XM2/a_n158_n73690# 0.010147f
C1732 XM1/a_n100_47409# XM2/a_n158_n107958# 0.005074f
C1733 XM1/a_n100_10073# XM2/a_n100_n142323# 1.24e-19
C1734 XM2/a_n158_n255574# XM3/a_n158_n48574# 4.64e-21
C1735 XM1/a_100_116434# XM2/a_n158_n36786# 0.079863f
C1736 XM1/a_n100_5765# XM2/a_100_n147498# 7.26e-20
C1737 XM1/a_100_n60194# XM4/w_n358_n132787# 0.054609f
C1738 XM1/a_100_69046# XM2/a_100_n84234# 4.64e-21
C1739 XM1/a_100_n111890# XM3/a_n100_n60067# 2.85e-20
C1740 XM1/a_n100_n99063# XM3/a_n100_n48671# 1.04e-19
C1741 XM4/w_n358_n132787# XM3/a_n158_n25782# 0.032295f
C1742 XM4/a_n100_n12411# m1_1634_n2388# 0.072014f
C1743 XM1/a_n100_n10031# m1_1634_n2388# 7.24e-20
C1744 XM2/a_n100_n139687# XM3/a_n158_64350# 0.002589f
C1745 XM1/a_n100_153673# XM2/a_100_118# 1.15e-19
C1746 XM2/a_100_n334654# XM3/a_n100_n130515# 0.005074f
C1747 XM1/a_n100_n68907# XM2/a_100_n223942# 7.26e-20
C1748 XM1/a_n100_n14339# XM2/a_n158_n168586# 0.010147f
C1749 XM1/a_100_41762# XM4/w_n358_n132787# 0.053325f
C1750 XM3/a_n100_88081# m1_1634_n2388# 0.072015f
C1751 XM4/a_n100_19705# m1_1634_n2388# 0.072015f
C1752 XM3/a_n100_45605# XM4/a_n100_45605# 0.009521f
C1753 XM1/a_n100_146493# XM2/a_n158_n7790# 0.010147f
C1754 XM1/a_n158_n42962# XM2/a_n158_n197582# 9.28e-21
C1755 XM4/w_n358_n132787# XM3/a_n100_n129479# 0.009186f
C1756 XM4/a_100_n114878# m1_1634_n2388# 6.1e-20
C1757 XM1/a_n158_n15678# XM3/a_n100_36281# 1.94e-20
C1758 XM2/a_100_n150134# m1_1634_n2388# 0.02391f
C1759 XM3/a_n100_33173# m1_1634_n2388# 0.072015f
C1760 XM1/a_n100_58897# m1_1634_n2388# 1.3e-19
C1761 XM1/a_n158_n177946# XM2/a_n158_n332018# 9.28e-21
C1762 XM1/a_n100_n162247# XM4/w_n358_n132787# 0.013401f
C1763 XM4/w_n358_n132787# XM2/a_n158_n218670# 0.107093f
C1764 XM1/a_n158_79098# XM3/a_n100_129521# 1.94e-20
C1765 XM2/a_n100_n184499# XM4/a_100_19802# 2.56e-20
C1766 XM1/a_100_113562# XM2/a_n158_n39422# 0.056885f
C1767 XM4/w_n358_n132787# XM4/a_n100_113981# -0.004445f
C1768 XM1/a_n158_n163586# XM2/a_n158_n316202# 4.64e-21
C1769 XM1/a_n100_n54547# XM2/a_100_n208126# 1.33e-19
C1770 XM4/w_n358_n132787# XM3/a_n158_74710# 0.032295f
C1771 XM2/a_100_n242394# XM3/a_n100_n37275# 0.010147f
C1772 XM1/a_100_n1318# XM4/w_n358_n132787# 0.048442f
C1773 XM1/a_n100_110593# XM4/w_n358_n132787# 0.012279f
C1774 XM1/a_n100_107721# XM2/a_n158_n44694# 0.005074f
C1775 XM4/w_n358_n132787# XM3/a_n158_106826# 0.038862f
C1776 XM1/a_100_n131994# XM2/a_n158_n284570# 0.017159f
C1777 XM1/a_100_77662# XM3/a_n100_128485# 2.85e-20
C1778 XM4/w_n358_n132787# XM3/a_n158_n65150# 0.032295f
C1779 XM4/a_n100_n51779# m1_1634_n2388# 0.072015f
C1780 XM2/a_100_n197582# XM3/a_n100_8309# 0.010147f
C1781 XM1/a_n100_n139271# XM2/a_n158_n292478# 0.005074f
C1782 XM4/w_n358_n132787# XM3/a_n158_19802# 0.038462f
C1783 XM1/a_n100_21561# m1_1634_n2388# 1.3e-19
C1784 XM1/a_100_n176510# XM2/a_100_n332018# 4.64e-21
C1785 XM1/a_100_173874# XM2/a_100_21206# 4.64e-21
C1786 XM2/a_100_n102686# XM3/a_n158_103718# 0.077526f
C1787 XM1/a_n100_n180915# m1_1634_n2388# 8.14e-20
C1788 XM1/a_100_n103274# XM2/a_n100_n255671# 1.17e-21
C1789 XM1/a_n100_n41623# XM2/a_n158_n197582# 0.002941f
C1790 XM1/a_n100_n43059# XM2/a_100_n197582# 1.45e-19
C1791 XM2/a_n158_n279298# XM3/a_n100_n72499# 7.26e-20
C1792 XM1/a_100_n110454# XM2/a_n158_n263482# 0.061169f
C1793 XM1/a_100_158078# XM2/a_100_2754# 4.64e-21
C1794 XM2/a_n100_n89603# m1_1634_n2388# 7.61e-19
C1795 XM1/a_100_n131994# XM3/a_n100_n79751# 2.85e-20
C1796 XM1/a_100_n77426# XM3/a_n100_n25879# 2.85e-20
C1797 XM1/a_100_n81734# XM2/a_n100_n237219# 0.005074f
C1798 XM2/a_100_n73690# XM4/w_n358_n132787# 0.084379f
C1799 XM1/a_n100_n107679# XM2/a_100_n263482# 7.26e-20
C1800 XM4/w_n358_n132787# XM2/a_100_n155406# 0.10476f
C1801 XM4/w_n358_n132787# XM4/a_n100_74613# -0.004445f
C1802 XM2/a_100_n274026# m1_1634_n2388# 0.017213f
C1803 XM1/a_n158_n4190# XM3/a_n100_46641# 1.94e-20
C1804 XM3/a_n100_n32095# m1_1634_n2388# 0.072015f
C1805 XM1/a_100_n17114# XM3/a_n100_33173# 2.46e-20
C1806 XM1/a_100_133666# XM4/w_n358_n132787# 0.048442f
C1807 XM1/a_n100_71821# XM3/a_n100_124341# 9.63e-19
C1808 XM1/a_100_58994# XM3/a_n100_110873# 2.85e-20
C1809 XM2/a_100_n115866# XM3/a_n100_88081# 0.005074f
C1810 XM3/a_n158_58134# m1_1634_n2388# 6.1e-20
C1811 XM4/w_n358_n132787# XM3/a_n158_n104518# 0.032641f
C1812 XM4/a_n100_n91147# m1_1634_n2388# 0.072015f
C1813 XM1/a_n100_n110551# XM3/a_n100_n59031# 1.19e-19
C1814 XM1/a_100_n86042# XM3/a_n100_n34167# 2.85e-20
C1815 XM1/a_n158_n63066# XM3/a_n100_n11375# 9.62e-21
C1816 XM2/a_n158_n310930# XM3/a_n158_n106590# 4.64e-21
C1817 XM2/a_n100_n113327# XM3/a_n158_93358# 0.005074f
C1818 XM1/a_n158_n123378# XM2/a_n158_n276662# 4.64e-21
C1819 XM2/a_100_n223942# XM3/a_n100_n19663# 0.005074f
C1820 XM2/a_n158_n84234# XM3/a_n100_120197# 7.26e-20
C1821 XM2/a_n100_n84331# XM3/a_n158_120294# 0.005074f
C1822 XM1/a_100_n47270# XM3/a_n158_4262# 0.00544f
C1823 XM1/a_100_61866# XM3/a_n100_112945# 2.85e-20
C1824 XM1/a_100_n154970# XM2/a_n100_n311027# 0.005074f
C1825 XM4/a_100_108898# m1_1634_n2388# 6.1e-20
C1826 XM1/a_n158_n177946# XM3/a_n100_n126371# 1.94e-20
C1827 XM2/a_100_n308294# XM3/a_n158_n101410# 0.030791f
C1828 XM1/a_n100_n47367# XM3/a_n158_3226# 2.85e-20
C1829 XM2/a_n100_n313663# XM4/a_100_n106590# 2.56e-20
C1830 XM2/a_n100_n205587# XM4/a_100_1154# 2.56e-20
C1831 XM4/w_n358_n132787# XM4/a_n100_35245# -0.004445f
C1832 XM1/a_n158_n81734# XM3/a_n100_n31059# 1.94e-20
C1833 XM1/a_n100_159417# XM2/a_n158_5390# 0.010147f
C1834 XM3/a_n100_n71463# m1_1634_n2388# 0.072015f
C1835 XM1/a_n100_84745# XM2/a_100_n71054# 7.26e-20
C1836 XM4/w_n358_n132787# XM2/a_n100_n94875# 0.025034f
C1837 XM1/a_100_18786# XM2/a_100_n134318# 4.64e-21
C1838 XM1/a_100_n140610# XM4/w_n358_n132787# 0.048442f
C1839 XM2/a_n100_n213495# m1_1634_n2388# 0.002141f
C1840 pbias sw_b 0.001381f
C1841 XM1/a_n100_n145015# XM3/a_n158_n94158# 2.85e-20
C1842 XM2/a_n158_n260846# XM3/a_n100_n54887# 1.45e-19
C1843 XM1/a_100_89150# XM2/a_n158_n65782# 0.10401f
C1844 XM4/a_n100_n130515# m1_1634_n2388# 0.072015f
C1845 XM3/a_n100_n17591# XM4/a_n100_n17591# 0.009521f
C1846 XM4/w_n358_n132787# XM2/a_100_n279298# 0.103579f
C1847 XM1/a_100_n113326# XM3/a_n100_n61103# 2.85e-20
C1848 XM1/a_n158_n107582# XM2/a_n158_n263482# 4.64e-21
C1849 XM2/a_n100_n13159# XM4/w_n358_n132787# 0.012279f
C1850 XM3/a_n100_108801# m1_1634_n2388# 0.072015f
C1851 XM1/a_n158_n173638# XM2/a_n100_n326843# 7.26e-20
C1852 XM1/a_n158_155206# XM2/a_n100_2657# 7.26e-20
C1853 XM1/a_n158_10170# XM2/a_n158_n144862# 4.64e-21
C1854 XM1/a_100_166694# XM2/a_n100_13201# 0.005074f
C1855 XM2/a_100_n144862# XM3/a_n100_60109# 0.010147f
C1856 XM1/a_n100_n120603# XM2/a_n100_n276759# 0.002448f
C1857 XM1/a_n158_n19986# XM3/a_n100_32137# 1.94e-20
C1858 XM1/a_n158_126486# XM2/a_n100_n28975# 7.26e-20
C1859 XM4/w_n358_n132787# XM4/a_n100_n36239# -0.004445f
C1860 XM1/a_n100_n83267# XM3/a_n158_n30962# 2.85e-20
C1861 XM3/a_n100_13489# XM4/a_n100_13489# 0.009521f
C1862 XM3/a_n100_98441# XM4/a_n100_98441# 0.009521f
C1863 XM2/a_n100_n255671# XM3/a_n158_n48574# 0.005074f
C1864 XM3/a_n158_n7134# m1_1634_n2388# 6.1e-20
C1865 XM1/a_n100_5765# XM2/a_n158_n147498# 0.005074f
C1866 XM1/a_100_n81734# XM4/w_n358_n132787# 0.054609f
C1867 XM2/a_100_n187038# XM3/a_n100_17633# 0.005074f
C1868 XM1/a_n158_77662# XM3/a_n100_128485# 1.94e-20
C1869 XM1/a_100_69046# XM2/a_n158_n84234# 0.085705f
C1870 XM4/a_100_69530# m1_1634_n2388# 6.1e-20
C1871 XM1/a_100_n101838# XM2/a_n158_n255574# 0.116862f
C1872 XM1/a_n100_n78959# XM2/a_100_n231850# 7.26e-20
C1873 XM1/a_n100_n122039# XM3/a_n158_n70330# 4.33e-21
C1874 XM2/a_n158_n334654# XM3/a_n100_n130515# 7.26e-20
C1875 XM3/a_n100_n110831# m1_1634_n2388# 0.072015f
C1876 XM1/a_n100_n68907# XM2/a_n158_n223942# 0.005074f
C1877 XM4/w_n358_n132787# XM3/a_n100_7273# 0.008969f
C1878 XM1/a_100_160950# XM2/a_100_8026# 4.64e-21
C1879 XM3/a_n100_n37275# XM4/a_n100_n37275# 0.009521f
C1880 XM1/a_n100_86181# XM4/w_n358_n132787# 0.012279f
C1881 XM4/w_n358_n132787# XM3/a_n100_68397# 0.009141f
C1882 XM2/a_n158_n150134# m1_1634_n2388# 2.36e-21
C1883 XM2/a_100_n289842# XM3/a_n158_n83798# 0.077916f
C1884 XM1/a_100_n180818# XM3/a_n100_n129479# 5.71e-20
C1885 XM2/a_100_n332018# XM3/a_n100_n125335# 0.005074f
C1886 XM1/a_n100_n143579# XM3/a_n158_n93122# 1.76e-20
C1887 XM4/w_n358_n132787# XM3/a_n100_n16555# 0.009161f
C1888 XM4/w_n358_n132787# XM2/a_n100_n218767# 0.025775f
C1889 XM4/a_100_n1954# m1_1634_n2388# 6.1e-20
C1890 XM2/a_100_n202854# XM3/a_n158_4262# 0.008202f
C1891 XM2/a_n158_29114# XM1/a_n158_182490# 4.64e-21
C1892 XM2/a_100_29114# XM1/a_n100_182393# 7.26e-20
C1893 XM2/a_n100_29017# XM1/a_100_182490# 0.005074f
C1894 XM2/a_n100_n337387# m1_1634_n2388# 3.8e-19
C1895 XM4/w_n358_n132787# XM3/a_n100_13489# 0.009186f
C1896 XM1/a_n158_n163586# XM2/a_n100_n316299# 7.26e-20
C1897 XM4/w_n358_n132787# XM4/a_n100_n75607# -0.004445f
C1898 XM1/a_n100_n54547# XM2/a_n158_n208126# 0.008992f
C1899 XM2/a_100_n131682# XM3/a_n100_74613# 0.00524f
C1900 XM1/a_n158_n160714# XM2/a_n158_n313566# 4.64e-21
C1901 XM3/a_n158_n46502# m1_1634_n2388# 6.1e-20
C1902 XM2/a_n158_n242394# XM3/a_n100_n37275# 1.45e-19
C1903 XM4/w_n358_n132787# XM3/a_n100_106729# 0.009186f
C1904 XM1/a_100_n131994# XM2/a_n100_n284667# 0.005074f
C1905 XM4/a_100_30162# m1_1634_n2388# 6.1e-20
C1906 XM1/a_n158_73354# XM3/a_n100_124341# 1.94e-20
C1907 XM2/a_n158_n197582# XM3/a_n100_8309# 1.45e-19
C1908 XM1/a_n158_107818# XM2/a_n100_n47427# 7.26e-20
C1909 XM2/a_100_n173858# XM3/a_n100_32137# 0.010147f
C1910 XM1/a_n100_n140707# XM3/a_n158_n90014# 2.85e-20
C1911 XM1/a_n100_n116295# XM4/w_n358_n132787# 0.01363f
C1912 XM2/a_n100_n181863# XM4/a_100_24982# 2.56e-20
C1913 XM1/a_n158_100638# XM2/a_n100_n52699# 7.26e-20
C1914 XM1/a_100_38890# XM2/a_n158_n115866# 0.116862f
C1915 XM1/a_100_n176510# XM2/a_n158_n332018# 0.047927f
C1916 XM1/a_100_n104710# XM3/a_n158_n53754# 0.002042f
C1917 XM2/a_n158_n102686# XM3/a_n158_103718# 4.64e-21
C1918 XM2/a_100_n102686# XM3/a_n100_103621# 0.005074f
C1919 XM1/a_n100_10073# XM3/a_n158_61242# 2.85e-20
C1920 XM1/a_100_n136302# m1_1634_n2388# 8.49e-19
C1921 XM1/a_n100_n41623# XM2/a_n100_n197679# 0.002209f
C1922 XM3/a_n100_n56959# XM4/a_n100_n56959# 0.009521f
C1923 XM1/a_n100_n43059# XM2/a_n158_n197582# 0.010147f
C1924 XM1/a_n100_109157# XM2/a_n158_n44694# 0.010147f
C1925 XM1/a_100_n110454# XM2/a_n100_n263579# 0.005074f
C1926 XM2/a_100_n86870# m1_1634_n2388# 0.025819f
C1927 XM4/a_n100_93261# m1_1634_n2388# 0.072015f
C1928 XM4/w_n358_n132787# XM3/a_n100_n55923# 0.008931f
C1929 XM4/a_100_n41322# m1_1634_n2388# 6.1e-20
C1930 XM3/a_n100_51821# m1_1634_n2388# 0.072015f
C1931 XM1/a_100_n81734# XM2/a_100_n234486# 4.64e-21
C1932 XM3/a_n100_131593# XM4/a_n100_131593# 0.01485f
C1933 XM1/a_n100_n107679# XM2/a_n158_n263482# 0.005074f
C1934 XM4/w_n358_n132787# XM2/a_n158_n155406# 0.107093f
C1935 XM4/w_n358_n132787# XM4/a_n100_n114975# -0.004445f
C1936 XM1/a_n158_n63066# XM2/a_n158_n218670# 4.64e-21
C1937 XM3/a_n158_n85870# m1_1634_n2388# 6.1e-20
C1938 XM1/a_100_60430# XM4/w_n358_n132787# 0.054609f
C1939 XM1/a_n158_146590# XM2/a_n158_n7790# 9.28e-21
C1940 XM4/w_n358_n132787# XM3/a_n158_93358# 0.037143f
C1941 XM2/a_n158_n115866# XM3/a_n100_88081# 7.26e-20
C1942 XM1/a_n100_n179479# m1_1634_n2388# 1.3e-19
C1943 XM2/a_100_n271390# XM3/a_n158_n66186# 0.077916f
C1944 XM1/a_100_97766# XM2/a_n100_n55335# 0.005074f
C1945 XM4/w_n358_n132787# XM3/a_n158_131690# 0.032295f
C1946 XM1/a_n100_74693# XM4/w_n358_n132787# 0.01363f
C1947 XM2/a_100_n313566# XM3/a_n100_n107723# 0.010147f
C1948 XM4/w_n358_n132787# XM3/a_n158_38450# 0.038462f
C1949 XM2/a_n100_n311027# XM3/a_n158_n106590# 0.005074f
C1950 XM3/a_n158_3226# m1_1634_n2388# 6.1e-20
C1951 XM1/a_100_n38654# XM3/a_n100_13489# 2.85e-20
C1952 XM1/a_n100_n31571# XM2/a_100_n187038# 7.26e-20
C1953 XM4/w_n358_n132787# XM1/a_100_n134866# 0.053188f
C1954 XM1/a_n158_n123378# XM2/a_n100_n276759# 7.26e-20
C1955 XM2/a_n158_n223942# XM3/a_n100_n19663# 7.26e-20
C1956 XM2/a_100_n84234# XM3/a_n158_121330# 0.077916f
C1957 XM3/a_n100_n76643# XM4/a_n100_n76643# 0.009521f
C1958 XM1/a_100_n154970# XM2/a_100_n308294# 4.64e-21
C1959 XM4/a_n100_53893# m1_1634_n2388# 0.072015f
C1960 XM2/a_n158_n308294# XM3/a_n158_n101410# 4.64e-21
C1961 XM4/w_n358_n132787# XM3/a_n100_n95291# 0.009036f
C1962 XM4/a_100_n80690# m1_1634_n2388# 6.1e-20
C1963 XM1/a_100_76226# XM2/a_100_n78962# 4.64e-21
C1964 XM2/a_100_n221306# XM3/a_n100_n14483# 0.005074f
C1965 XM1/a_n100_n61727# XM3/a_n100_n11375# 6.24e-19
C1966 XM4/a_n100_3129# m1_1634_n2388# 0.072015f
C1967 XM3/a_n158_n125238# m1_1634_n2388# 6.1e-20
C1968 XM2/a_n100_n15795# XM1/a_n158_139410# 7.26e-20
C1969 XM2/a_n158_n15698# XM1/a_100_139410# 0.086873f
C1970 XM4/w_n358_n132787# XM2/a_100_n92142# 0.106018f
C1971 XM1/a_100_18786# XM2/a_n158_n134318# 0.068569f
C1972 XM1/a_n158_n182254# avdd 0.011771f
C1973 XM1/a_100_n104710# XM2/a_100_n258210# 4.64e-21
C1974 XM2/a_100_n210762# m1_1634_n2388# 0.017213f
C1975 XM3/a_n100_66325# XM4/a_n100_66325# 0.009521f
C1976 XM1/a_100_73354# XM2/a_n100_n79059# 4.8e-19
C1977 XM4/w_n358_n132787# XM2/a_n158_n279298# 0.107093f
C1978 XM1/a_n100_149365# XM2/a_n158_n5154# 0.010147f
C1979 XM1/a_n100_87617# XM2/a_n100_n68515# 0.004948f
C1980 XM3/a_n158_76782# m1_1634_n2388# 6.1e-20
C1981 XM1/a_n158_n107582# XM2/a_n100_n263579# 7.26e-20
C1982 XM1/a_n100_159417# XM4/w_n358_n132787# 0.012279f
C1983 XM1/a_n100_n163683# XM3/a_n158_n111770# 2.85e-20
C1984 XM4/w_n358_n132787# XM3/a_n158_n30962# 0.032295f
C1985 XM4/a_n100_n17591# m1_1634_n2388# 0.072015f
C1986 XM1/a_n158_10170# XM2/a_n100_n144959# 7.26e-20
C1987 XM1/a_100_n5626# m1_1634_n2388# 0.002547f
C1988 XM2/a_n158_n144862# XM3/a_n100_60109# 1.45e-19
C1989 XM1/a_n100_n120603# XM2/a_100_n274026# 7.26e-20
C1990 XM3/a_n158_21874# m1_1634_n2388# 6.1e-20
C1991 XM1/a_n100_47409# XM2/a_100_n105322# 7.26e-20
C1992 XM1/a_n158_n100402# XM3/a_n100_n48671# 1.94e-20
C1993 XM1/a_n100_67513# XM2/a_100_n86870# 1.45e-19
C1994 XM3/a_n100_115017# XM4/a_n100_115017# 0.009521f
C1995 XM3/a_n100_n96327# XM4/a_n100_n96327# 0.009521f
C1996 XM2/a_100_n252938# XM3/a_n158_n48574# 0.035464f
C1997 XM2/a_n100_n258307# XM4/a_100_n53754# 2.56e-20
C1998 XM4/a_n100_14525# m1_1634_n2388# 0.072015f
C1999 XM2/a_n158_n187038# XM3/a_n100_17633# 7.26e-20
C2000 XM1/a_100_69046# XM2/a_n100_n84331# 0.005074f
C2001 XM1/a_100_46070# XM3/a_n100_98441# 9.33e-21
C2002 XM2/a_100_n295114# XM3/a_n100_n90111# 0.010147f
C2003 XM1/a_n100_n78959# XM2/a_n158_n231850# 0.005074f
C2004 XM1/a_n100_45973# XM2/a_100_n107958# 1.45e-19
C2005 XM4/a_100_n120058# m1_1634_n2388# 6.1e-20
C2006 XM1/a_n158_158078# XM2/a_n100_5293# 7.26e-20
C2007 XM1/a_n100_64641# XM2/a_100_n89506# 1.45e-19
C2008 XM2/a_100_n139590# XM3/a_n158_65386# 0.077916f
C2009 XM1/a_n100_n94755# XM4/w_n358_n132787# 0.013474f
C2010 XM1/a_n100_21# XM2/a_100_n155406# 7.26e-20
C2011 XM2/a_100_n181766# XM3/a_n158_22910# 0.065842f
C2012 XM4/w_n358_n132787# XM4/a_n100_108801# -0.004445f
C2013 XM1/a_100_148026# XM2/a_100_n5154# 4.64e-21
C2014 XM2/a_n100_n150231# m1_1634_n2388# 9.17e-19
C2015 XM1/a_n100_n57419# XM2/a_100_n213398# 1.97e-20
C2016 XM1/a_n100_40229# XM2/a_100_n113230# 7.26e-20
C2017 XM2/a_n158_n332018# XM3/a_n100_n125335# 7.26e-20
C2018 XM1/a_100_n165022# XM4/w_n358_n132787# 0.048442f
C2019 XM4/w_n358_n132787# XM3/a_n158_n70330# 0.032295f
C2020 XM4/a_n100_n56959# m1_1634_n2388# 0.072015f
C2021 XM4/w_n358_n132787# XM2/a_100_n216034# 0.103341f
C2022 XM2/a_n158_n202854# XM3/a_n158_4262# 4.64e-21
C2023 XM1/a_100_41762# XM2/a_n100_n110691# 0.003994f
C2024 XM2/a_100_n334654# m1_1634_n2388# 0.019967f
C2025 XM1/a_n158_n172202# XM2/a_n158_n326746# 9.28e-21
C2026 XM1/a_n100_n101935# XM2/a_100_n255574# 1.45e-19
C2027 XM2/a_n158_n7790# XM1/a_n158_145154# 4.64e-21
C2028 XM2/a_100_n7790# XM1/a_100_145154# 4.64e-21
C2029 XM1/a_n100_25869# m1_1634_n2388# 1.13e-19
C2030 XM1/a_100_n57322# XM4/w_n358_n132787# 0.053079f
C2031 XM1/a_100_n35782# XM3/a_n100_15561# 5.71e-20
C2032 XM1/a_100_n96094# XM3/a_n100_n44527# 2.85e-20
C2033 XM1/a_n100_n54547# XM2/a_n100_n208223# 5.53e-19
C2034 XM2/a_n158_n131682# XM3/a_n100_74613# 7.85e-20
C2035 XM3/a_n100_n116011# XM4/a_n100_n116011# 0.009521f
C2036 XM1/a_n158_n160714# XM2/a_n100_n313663# 7.26e-20
C2037 XM1/a_100_n34346# XM2/a_100_n189674# 4.64e-21
C2038 XM1/a_100_n12806# XM3/a_n100_38353# 4.58e-20
C2039 XM1/a_n158_n35782# XM3/a_n100_14525# 1.94e-20
C2040 XM2/a_100_n13062# XM1/a_100_142282# 4.64e-21
C2041 XM1/a_100_54686# XM3/a_n100_105693# 2.85e-20
C2042 XM2/a_n158_n173858# XM3/a_n100_32137# 1.45e-19
C2043 XM2/a_100_23842# XM1/a_100_179618# 4.64e-21
C2044 XM1/a_n100_152237# XM2/a_n100_21# 3.11e-19
C2045 XM1/a_100_80534# XM4/w_n358_n132787# 0.048442f
C2046 XM1/a_100_n176510# XM2/a_n100_n332115# 0.005074f
C2047 XM1/a_n100_165161# XM4/w_n358_n132787# 0.012279f
C2048 XM2/a_100_n126410# XM3/a_n158_79890# 0.077916f
C2049 XM1/a_100_110690# XM2/a_n158_n42058# 0.033906f
C2050 XM2/a_n100_n102783# XM3/a_n158_103718# 8.54e-20
C2051 XM2/a_n158_n102686# XM3/a_n100_103621# 7.26e-20
C2052 XM1/a_100_10170# XM3/a_n100_62181# 2.85e-20
C2053 XM1/a_n100_n41623# XM2/a_100_n194946# 7.26e-20
C2054 XM4/w_n358_n132787# XM4/a_n100_69433# -0.004445f
C2055 XM1/a_100_n61630# XM3/a_n100_n10339# 5.71e-20
C2056 XM2/a_100_n168586# XM3/a_n158_37414# 0.077916f
C2057 XM1/a_100_150898# XM2/a_n158_n2518# 0.098947f
C2058 XM2/a_100_n276662# XM3/a_n100_n72499# 0.005074f
C2059 XM3/a_n100_n37275# m1_1634_n2388# 0.072015f
C2060 XM1/a_n158_n9934# XM3/a_n158_40522# 1.14e-21
C2061 XM1/a_n100_2893# XM3/a_n158_53990# 2.85e-20
C2062 XM4/w_n358_n132787# XM3/a_n100_87045# 0.009077f
C2063 XM4/w_n358_n132787# XM3/a_n158_n109698# 0.034634f
C2064 XM4/a_n100_n96327# m1_1634_n2388# 0.072015f
C2065 XM1/a_100_n81734# XM2/a_n158_n234486# 0.034296f
C2066 XM4/w_n358_n132787# XM2/a_n100_n155503# 0.024598f
C2067 XM1/a_n100_28741# XM2/a_100_n126410# 7.26e-20
C2068 XM2/a_n100_n274123# m1_1634_n2388# 0.001787f
C2069 XM1/a_n158_n63066# XM2/a_n100_n218767# 7.26e-20
C2070 XM4/w_n358_n132787# XM3/a_n100_32137# 0.009186f
C2071 XM1/a_n158_54686# XM3/a_n100_105693# 1.94e-20
C2072 XM2/a_n100_n126507# XM4/a_100_77818# 2.56e-20
C2073 XM4/w_n358_n132787# XM3/a_n100_131593# 0.013085f
C2074 XM4/w_n358_n132787# XM4/a_n100_n2051# -0.004445f
C2075 XM2/a_n158_n313566# XM3/a_n100_n107723# 1.45e-19
C2076 XM1/a_100_n15678# XM3/a_n100_36281# 2.85e-20
C2077 XM1/a_n158_n175074# XM3/a_n100_n123263# 1.94e-20
C2078 XM1/a_100_152334# XM2/a_100_n2518# 4.64e-21
C2079 XM4/a_100_103718# m1_1634_n2388# 6.1e-20
C2080 XM1/a_n100_n31571# XM2/a_n158_n187038# 0.005074f
C2081 XM1/a_n100_91925# XM2/a_100_n60510# 7.26e-20
C2082 XM2/a_100_n84234# XM3/a_n100_121233# 0.010147f
C2083 XM4/w_n358_n132787# XM4/a_n100_30065# -0.004445f
C2084 XM3/a_n100_34209# XM4/a_n100_34209# 0.009521f
C2085 XM2/a_n158_n42058# XM4/w_n358_n132787# 0.107093f
C2086 XM3/a_n100_n76643# m1_1634_n2388# 0.072015f
C2087 XM1/a_100_n154970# XM2/a_n158_n308294# 0.089989f
C2088 XM2/a_n100_n308391# XM3/a_n158_n101410# 0.005074f
C2089 XM1/a_n100_n122039# XM2/a_100_n276662# 1.36e-19
C2090 XM1/a_100_76226# XM2/a_n158_n78962# 0.079084f
C2091 XM2/a_n158_n221306# XM3/a_n100_n14483# 7.26e-20
C2092 XM1/a_n158_94894# XM2/a_n100_n60607# 7.26e-20
C2093 XM3/a_n100_70469# m1_1634_n2388# 0.072015f
C2094 XM1/a_100_n119070# XM2/a_100_n274026# 4.64e-21
C2095 XM2/a_100_n197582# XM3/a_n158_9442# 0.017159f
C2096 XM1/a_n158_n47270# XM3/a_n100_3129# 1.94e-20
C2097 XM4/w_n358_n132787# XM2/a_n158_n92142# 0.107093f
C2098 XM1/a_100_18786# XM2/a_n100_n134415# 0.005074f
C2099 XM1/a_100_n104710# XM2/a_n158_n258210# 0.107125f
C2100 XM1/a_n100_77565# m1_1634_n2388# 1.3e-19
C2101 XM1/a_100_n160714# XM3/a_n100_n108759# 2.85e-20
C2102 XM3/a_n100_15561# m1_1634_n2388# 0.072014f
C2103 XM4/w_n358_n132787# XM4/a_n100_n41419# -0.004445f
C2104 XM3/a_n158_n12314# m1_1634_n2388# 6.1e-20
C2105 XM4/w_n358_n132787# XM2/a_n100_n279395# 0.024842f
C2106 XM1/a_100_14478# XM4/w_n358_n132787# 0.048442f
C2107 XM1/a_100_n144918# XM3/a_n100_n94255# 2.85e-20
C2108 XM3/a_n158_109934# m1_1634_n2388# 6.1e-20
C2109 XM4/a_100_64350# m1_1634_n2388# 6.1e-20
C2110 XM1/a_n100_n173735# XM3/a_n100_n121191# 6.5e-19
C2111 XM1/a_100_n142046# XM2/a_100_n297750# 4.64e-21
C2112 XM4/w_n358_n132787# XM3/a_n158_57098# 0.037486f
C2113 XM1/a_n100_n120603# XM2/a_n158_n274026# 0.005074f
C2114 XM1/a_n100_47409# XM2/a_n158_n105322# 0.005074f
C2115 XM1/a_n158_n123378# XM3/a_n100_n71463# 1.94e-20
C2116 XM1/a_100_n55886# XM3/a_n100_n5159# 2.85e-20
C2117 XM1/a_n100_67513# XM2/a_n158_n86870# 0.010147f
C2118 XM3/a_n100_n116011# m1_1634_n2388# 0.072014f
C2119 XM2/a_n158_n252938# XM3/a_n158_n48574# 4.64e-21
C2120 XM1/a_100_n143482# XM3/a_n100_n91147# 1.99e-20
C2121 XM2/a_n100_n187135# XM3/a_n100_17633# 0.003522f
C2122 XM1/a_n158_n160714# XM3/a_n100_n109795# 9.42e-21
C2123 XM2/a_n158_n295114# XM3/a_n100_n90111# 1.45e-19
C2124 XM1/a_n100_45973# XM2/a_n158_n107958# 0.010147f
C2125 XM1/a_n100_64641# XM2/a_n158_n89506# 0.010147f
C2126 XM1/a_100_84842# XM2/a_n100_n68515# 0.005074f
C2127 XM1/a_n158_n129122# XM3/a_n100_n78715# 1.94e-20
C2128 XM1/a_n100_n114859# XM4/w_n358_n132787# 0.013589f
C2129 XM1/a_n158_n98966# XM3/a_n100_n47635# 3.89e-20
C2130 XM4/a_n100_127449# m1_1634_n2388# 0.072015f
C2131 XM2/a_100_n250302# XM3/a_n158_n43394# 0.028454f
C2132 XM4/w_n358_n132787# XM3/a_n100_n21735# 0.009186f
C2133 XM1/a_n100_n68907# XM2/a_100_n221306# 7.26e-20
C2134 XM4/a_100_n7134# m1_1634_n2388# 6.1e-20
C2135 XM1/a_n100_21# XM2/a_n158_n155406# 0.005074f
C2136 XM2/a_n100_n255671# XM4/a_100_n48574# 2.56e-20
C2137 XM2/a_n158_n181766# XM3/a_n158_22910# 4.64e-21
C2138 XM1/a_n100_n53111# m1_1634_n2388# 1.3e-19
C2139 XM1/a_100_119306# XM2/a_n100_n36883# 1.06e-19
C2140 XM1/a_n158_58994# XM3/a_n100_109837# 1.94e-20
C2141 XM4/w_n358_n132787# XM4/a_n100_n80787# -0.004445f
C2142 XM2/a_100_n147498# m1_1634_n2388# 0.017213f
C2143 XM3/a_n158_n51682# m1_1634_n2388# 6.1e-20
C2144 XM1/a_n100_n57419# XM2/a_n158_n213398# 0.001183f
C2145 XM1/a_n100_40229# XM2/a_n158_n113230# 0.005074f
C2146 XM4/a_100_24982# m1_1634_n2388# 6.1e-20
C2147 XM1/a_100_28838# XM3/a_n158_80926# 0.002042f
C2148 XM4/w_n358_n132787# XM2/a_n158_n216034# 0.107093f
C2149 XM2/a_n100_n202951# XM3/a_n158_4262# 0.005074f
C2150 XM3/a_n158_95430# m1_1634_n2388# 6.1e-20
C2151 XM2/a_n158_n334654# m1_1634_n2388# 2.36e-21
C2152 XM1/a_n100_n101935# XM2/a_n158_n255574# 0.010147f
C2153 XM1/a_n158_79098# XM3/a_n100_130557# 2.83e-20
C2154 XM1/a_100_n175074# XM3/a_n100_n123263# 2.85e-20
C2155 XM1/a_n158_n83170# XM3/a_n100_n32095# 1.94e-20
C2156 XM2/a_n100_n131779# XM3/a_n100_74613# 0.005829f
C2157 XM3/a_n158_40522# m1_1634_n2388# 6.1e-20
C2158 XM4/w_n358_n132787# XM3/a_n158_107862# 0.032295f
C2159 XM1/a_100_n34346# XM2/a_n158_n189674# 0.065453f
C2160 XM1/a_100_77662# XM3/a_n100_129521# 2.85e-20
C2161 XM2/a_100_n324110# XM3/a_n158_n119022# 0.077916f
C2162 XM1/a_100_n176510# XM2/a_100_n329382# 4.64e-21
C2163 XM1/a_100_n63066# XM4/w_n358_n132787# 0.05487f
C2164 XM2/a_n100_n102783# XM3/a_n100_103621# 0.006262f
C2165 XM4/a_n100_88081# m1_1634_n2388# 0.072015f
C2166 XM1/a_n158_23094# XM3/a_n100_74613# 1.94e-20
C2167 XM4/w_n358_n132787# XM3/a_n100_n61103# 0.009186f
C2168 XM4/a_100_n46502# m1_1634_n2388# 6.1e-20
C2169 XM1/a_n158_33146# XM2/a_n158_n121138# 9.28e-21
C2170 XM1/a_100_8734# XM3/a_n100_59073# 2.85e-20
C2171 XM1/a_n100_n41623# XM2/a_n158_n194946# 0.005074f
C2172 XM4/w_n358_n132787# XM4/a_n100_n120155# -0.004445f
C2173 XM3/a_n158_n91050# m1_1634_n2388# 6.1e-20
C2174 XM2/a_n158_n276662# XM3/a_n100_n72499# 7.26e-20
C2175 XM1/a_100_n9934# XM3/a_n100_41461# 6.29e-19
C2176 XM1/a_100_2990# XM3/a_n100_54929# 2.85e-20
C2177 XM2/a_n100_n23703# XM1/a_100_132230# 0.005074f
C2178 XM2/a_n158_n23606# XM1/a_n100_130697# 0.010147f
C2179 XM2/a_n100_n86967# m1_1634_n2388# 7.61e-19
C2180 XM1/a_n158_n22858# XM3/a_n100_27993# 1.94e-20
C2181 XM1/a_100_n81734# XM2/a_n100_n234583# 0.005074f
C2182 XM1/a_100_n2754# XM3/a_n158_48810# 0.00544f
C2183 XM1/a_n158_71918# XM3/a_n158_122366# 2.84e-22
C2184 XM1/a_n100_n107679# XM2/a_100_n260846# 7.26e-20
C2185 XM2/a_100_n231850# XM3/a_n158_n25782# 0.077916f
C2186 XM4/w_n358_n132787# XM2/a_100_n152770# 0.103342f
C2187 XM1/a_n100_28741# XM2/a_n158_n126410# 0.005074f
C2188 XM2/a_100_n271390# m1_1634_n2388# 0.023368f
C2189 XM2/a_100_n274026# XM3/a_n100_n67319# 0.005074f
C2190 XM1/a_n100_n67471# XM2/a_100_n221306# 1.45e-19
C2191 XM3/a_n100_87045# XM4/a_n100_87045# 0.009521f
C2192 XM1/a_n100_n67471# XM3/a_n158_n15422# 2.85e-20
C2193 XM1/a_n100_n17211# XM3/a_n100_35245# 7.28e-19
C2194 XM2/a_n100_n57971# XM4/w_n358_n132787# 0.012279f
C2195 XM4/w_n358_n132787# XM3/a_n158_8406# 0.032295f
C2196 XM2/a_100_23842# XM1/a_n100_178085# 1.45e-19
C2197 XM4/a_n100_48713# m1_1634_n2388# 0.072015f
C2198 XM4/w_n358_n132787# XM3/a_n100_n100471# 0.009026f
C2199 XM4/a_100_n85870# m1_1634_n2388# 6.1e-20
C2200 XM1/a_n158_n80298# XM2/a_n158_n234486# 9.28e-21
C2201 XM1/a_n100_76129# XM2/a_100_n78962# 7.26e-20
C2202 XM2/a_n158_n84234# XM3/a_n100_121233# 1.45e-19
C2203 XM2/a_n100_n110691# XM3/a_n158_93358# 0.003644f
C2204 XM2/a_n100_n123871# XM4/a_100_82998# 2.56e-20
C2205 XM1/a_n158_n176510# XM3/a_n100_n125335# 3.39e-20
C2206 XM1/a_100_n60194# XM3/a_n100_n9303# 2.85e-20
C2207 XM1/a_100_163822# XM2/a_n158_8026# 0.019886f
C2208 XM1/a_100_61866# XM3/a_n100_113981# 2.85e-20
C2209 sw_bn XM4/w_n358_n132787# 0.003128f
C2210 XM3/a_n158_n130418# m1_1634_n2388# 6.1e-20
C2211 XM1/a_100_n147790# XM3/a_n100_n96327# 4.11e-20
C2212 XM1/a_n158_97766# XM2/a_n100_n57971# 7.26e-20
C2213 XM1/a_100_n154970# XM2/a_n100_n308391# 0.005074f
C2214 XM1/a_100_n147790# XM2/a_100_n303022# 4.64e-21
C2215 XM2/a_100_n305658# XM3/a_n158_n101410# 0.02417f
C2216 XM1/a_n100_n122039# XM2/a_n158_n276662# 0.009343f
C2217 XM2/a_n100_n311027# XM4/a_100_n106590# 2.56e-20
C2218 XM1/a_100_n142046# XM4/w_n358_n132787# 0.054609f
C2219 XM1/a_100_76226# XM2/a_n100_n79059# 0.005074f
C2220 XM2/a_n100_n202951# XM4/a_100_1154# 2.56e-20
C2221 XM1/a_100_n119070# XM2/a_n158_n274026# 0.101673f
C2222 XM2/a_n158_n197582# XM3/a_n158_9442# 4.64e-21
C2223 XM4/w_n358_n132787# XM3/a_n158_n36142# 0.032295f
C2224 XM4/a_n100_n22771# m1_1634_n2388# 0.072015f
C2225 XM4/w_n358_n132787# XM2/a_n100_n92239# 0.024666f
C2226 XM1/a_100_n104710# XM2/a_n100_n258307# 0.005074f
C2227 XM2/a_n100_n210859# m1_1634_n2388# 7.61e-19
C2228 XM1/a_n100_n2851# m1_1634_n2388# 9.43e-20
C2229 XM4/w_n358_n132787# XM3/a_n100_50785# 0.009186f
C2230 XM1/a_n158_n131994# XM2/a_n158_n287206# 4.64e-21
C2231 XM1/a_100_n24294# XM3/a_n158_28090# 6.08e-19
C2232 XM4/w_n358_n132787# XM2/a_100_n276662# 0.103997f
C2233 XM1/a_n158_n107582# XM2/a_n158_n260846# 4.64e-21
C2234 XM4/a_n100_9345# m1_1634_n2388# 0.072015f
C2235 XM3/a_n100_109837# m1_1634_n2388# 0.072015f
C2236 XM4/a_100_n125238# m1_1634_n2388# 6.1e-20
C2237 XM2/a_100_n213398# XM3/a_n158_n8170# 0.077916f
C2238 XM1/a_100_n142046# XM2/a_n158_n297750# 0.028843f
C2239 XM1/a_n158_44634# XM3/a_n100_96369# 1.94e-20
C2240 XM1/a_n100_n120603# XM2/a_n100_n274123# 6.38e-19
C2241 XM2/a_100_n255574# XM3/a_n100_n49707# 0.010147f
C2242 XM1/a_n100_n60291# XM2/a_100_n216034# 7.26e-20
C2243 XM2/a_n100_n253035# XM3/a_n158_n48574# 0.005074f
C2244 XM1/a_100_n140610# XM2/a_n158_n295114# 0.116862f
C2245 XM1/a_n158_77662# XM3/a_n100_129521# 1.94e-20
C2246 XM1/a_100_n134866# XM3/a_n100_n82859# 2.85e-20
C2247 XM1/a_100_n54450# XM2/a_n158_n208126# 0.116862f
C2248 XM1/a_n100_n20083# XM3/a_n158_31198# 5.5e-21
C2249 XM4/w_n358_n132787# XM4/a_n100_103621# -0.004445f
C2250 XM1/a_n158_n179382# XM2/a_n158_n334654# 4.64e-21
C2251 XM1/a_n158_n143482# XM2/a_n158_n297750# 9.28e-21
C2252 XM1/a_100_n28602# XM4/w_n358_n132787# 0.054853f
C2253 XM1/a_n100_31613# XM3/a_n158_84034# 2.85e-20
C2254 XM4/w_n358_n132787# XM3/a_n158_n75510# 0.033018f
C2255 XM4/a_n100_n62139# m1_1634_n2388# 0.072015f
C2256 XM2/a_n158_n250302# XM3/a_n158_n43394# 4.64e-21
C2257 XM1/a_n100_n68907# XM2/a_n158_n221306# 0.005074f
C2258 XM3/a_n100_89117# m1_1634_n2388# 0.072015f
C2259 XM1/a_n100_n167991# XM2/a_100_n321474# 7.26e-20
C2260 XM2/a_n100_n181863# XM3/a_n158_22910# 0.005074f
C2261 XM1/a_n100_30177# m1_1634_n2388# 1.23e-19
C2262 XM1/a_n158_n24294# XM3/a_n158_28090# 1.14e-21
C2263 XM1/a_n100_n94755# XM3/a_n100_n43491# 4.29e-19
C2264 XM1/a_n158_n65938# XM3/a_n100_n14483# 2.91e-20
C2265 XM1/a_n100_n57419# XM2/a_n100_n213495# 0.003456f
C2266 XM3/a_n100_34209# m1_1634_n2388# 0.072015f
C2267 XM1/a_n100_40229# XM2/a_n100_n113327# 0.002599f
C2268 XM2/a_100_n329382# XM3/a_n100_n125335# 0.005074f
C2269 XM4/w_n358_n132787# XM2/a_n100_n216131# 0.024993f
C2270 XM2/a_100_n200218# XM3/a_n158_4262# 0.046759f
C2271 XM1/a_n158_80534# XM2/a_n158_n73690# 9.28e-21
C2272 XM2/a_n100_n334751# m1_1634_n2388# 0.001789f
C2273 XM1/a_n158_n14242# XM3/a_n100_36281# 1.94e-20
C2274 XM1/a_n100_n11467# XM4/w_n358_n132787# 0.01363f
C2275 XM1/a_n158_n180818# XM3/a_n100_n128443# 5.01e-21
C2276 XM1/a_100_n163586# XM3/a_n100_n111867# 2.85e-20
C2277 XM4/w_n358_n132787# XM3/a_n158_75746# 0.032515f
C2278 XM4/w_n358_n132787# XM3/a_n100_107765# 0.00888f
C2279 XM1/a_100_n34346# XM2/a_n100_n189771# 0.005074f
C2280 XM1/a_n158_73354# XM3/a_n100_125377# 1.94e-20
C2281 XM1/a_n100_n132091# m1_1634_n2388# 9.25e-20
C2282 XM1/a_n100_n124911# m1_1634_n2388# 8.14e-20
C2283 XM1/a_n158_n64502# XM3/a_n100_n13447# 1.94e-20
C2284 XM1/a_n100_157981# XM2/a_100_2754# 7.26e-20
C2285 XM4/w_n358_n132787# XM4/a_n100_64253# -0.004445f
C2286 XM3/a_n100_n42455# m1_1634_n2388# 0.072015f
C2287 XM4/w_n358_n132787# XM3/a_n158_20838# 0.032295f
C2288 XM2/a_n100_n179227# XM4/a_100_24982# 2.56e-20
C2289 XM1/a_100_n7062# XM3/a_n100_43533# 2.85e-20
C2290 XM1/a_100_34582# XM4/w_n358_n132787# 0.054715f
C2291 XM1/a_n100_31613# XM2/a_100_n123774# 7.26e-20
C2292 XM1/a_100_n176510# XM2/a_n158_n329382# 0.04598f
C2293 XM1/a_n100_n89011# XM2/a_n100_n245127# 0.00473f
C2294 XM4/w_n358_n132787# XM3/a_n158_n114878# 0.037235f
C2295 XM4/a_n100_n101507# m1_1634_n2388# 0.072015f
C2296 XM2/a_100_n237122# XM3/a_n100_n32095# 0.010147f
C2297 XM2/a_100_n73690# XM4/a_100_131690# 1.51e-21
C2298 XM1/a_n100_27305# XM2/a_100_n126410# 1.45e-19
C2299 XM1/a_100_n107582# XM3/a_n100_n56959# 8.73e-20
C2300 XM1/a_n100_1457# XM3/a_n100_53893# 4.68e-19
C2301 XM3/a_n100_54929# XM4/a_n100_54929# 0.009521f
C2302 XM1/a_n158_n42962# XM3/a_n100_8309# 3.89e-20
C2303 XM1/a_100_n37218# XM3/a_n100_13489# 2.85e-20
C2304 XM1/a_n100_74693# XM3/a_n158_125474# 2.85e-20
C2305 XM2/a_100_n84234# m1_1634_n2388# 0.017213f
C2306 XM4/w_n358_n132787# XM4/a_n100_n7231# -0.004445f
C2307 XM1/a_n158_71918# XM3/a_n100_122269# 1.22e-20
C2308 XM1/a_n158_n116198# XM2/a_n158_n271390# 4.64e-21
C2309 XM1/a_n100_n107679# XM2/a_n158_n260846# 0.005074f
C2310 XM1/a_n100_n28699# XM3/a_n100_22813# 5.85e-20
C2311 XM4/w_n358_n132787# XM2/a_n158_n152770# 0.107093f
C2312 XM2/a_n100_5293# XM4/w_n358_n132787# 0.012279f
C2313 XM1/a_n158_n63066# XM2/a_n158_n216034# 4.64e-21
C2314 XM1/a_n158_n4190# XM3/a_n100_47677# 1.94e-20
C2315 XM4/a_100_98538# m1_1634_n2388# 6.1e-20
C2316 XM1/a_n158_n130558# XM2/a_n158_n284570# 9.28e-21
C2317 XM2/a_n158_n274026# XM3/a_n100_n67319# 7.26e-20
C2318 XM1/a_n100_n67471# XM2/a_n158_n221306# 0.010147f
C2319 XM1/a_100_n17114# XM3/a_n100_34209# 5.71e-20
C2320 XM2/a_100_n115866# XM3/a_n100_89117# 0.010147f
C2321 XM4/w_n358_n132787# XM4/a_n100_24885# -0.004445f
C2322 XM1/a_n158_99202# XM2/a_n158_n55238# 9.28e-21
C2323 XM3/a_n158_59170# m1_1634_n2388# 6.1e-20
C2324 XM3/a_n100_n81823# m1_1634_n2388# 0.072015f
C2325 XM1/a_100_56122# XM4/w_n358_n132787# 0.049898f
C2326 XM2/a_100_n158042# XM3/a_n100_46641# 0.005074f
C2327 XM1/a_n100_n31571# XM2/a_100_n184402# 7.26e-20
C2328 XM3/a_n100_n22771# XM4/a_n100_n22771# 0.009521f
C2329 XM1/a_n100_76129# XM2/a_n158_n78962# 0.005074f
C2330 XM2/a_100_n84234# XM3/a_n158_122366# 0.058442f
C2331 XM1/a_n100_126389# XM2/a_n158_n28878# 0.005074f
C2332 XM1/a_n158_n182254# XM4/w_n358_n132787# 1.14e-31
C2333 XM1/a_n100_n61727# XM2/a_100_n216034# 1.45e-19
C2334 XM1/a_n158_171002# XM2/a_n158_15934# 4.64e-21
C2335 avdd XM2/a_n100_n337387# 1.41e-20
C2336 XM1/a_n158_n130558# XM3/a_n100_n79751# 1.94e-20
C2337 XM1/a_100_n147790# XM2/a_n158_n303022# 0.0748f
C2338 XM2/a_n158_n305658# XM3/a_n158_n101410# 4.64e-21
C2339 XM1/a_n100_n122039# XM2/a_n100_n276759# 6.38e-19
C2340 XM1/a_n100_n20083# m1_1634_n2388# 7.54e-20
C2341 XM4/w_n358_n132787# XM4/a_n100_n46599# -0.004445f
C2342 XM3/a_n158_n17494# m1_1634_n2388# 6.1e-20
C2343 XM1/a_100_76226# XM2/a_100_n76326# 4.64e-21
C2344 XM2/a_100_n218670# XM3/a_n100_n14483# 0.005074f
C2345 XM1/a_100_n119070# XM2/a_n100_n274123# 0.005074f
C2346 XM2/a_n100_n197679# XM3/a_n158_9442# 0.005074f
C2347 XM4/a_100_59170# m1_1634_n2388# 6.1e-20
C2348 XM1/a_n100_84745# XM2/a_100_n68418# 7.26e-20
C2349 XM4/w_n358_n132787# XM2/a_100_n89506# 0.103342f
C2350 XM1/a_100_57558# XM2/a_100_n97414# 4.64e-21
C2351 XM1/a_n100_12945# XM2/a_100_n142226# 7.26e-20
C2352 XM2/a_100_n208126# m1_1634_n2388# 0.025343f
C2353 XM2/a_100_n303022# XM3/a_n158_n96230# 0.039748f
C2354 XM1/a_n158_n131994# XM2/a_n100_n287303# 7.26e-20
C2355 XM1/a_100_n70246# XM4/w_n358_n132787# 0.048442f
C2356 XM2/a_n100_n308391# XM4/a_100_n101410# 2.56e-20
C2357 XM3/a_n100_n121191# m1_1634_n2388# 0.072015f
C2358 XM4/w_n358_n132787# XM2/a_n158_n276662# 0.103279f
C2359 XM1/a_n158_129358# XM2/a_n158_n26242# 4.64e-21
C2360 XM1/a_n158_n107582# XM2/a_n100_n260943# 7.26e-20
C2361 XM2/a_n100_n10523# XM4/w_n358_n132787# 0.012279f
C2362 XM1/a_n158_47506# XM2/a_n158_n107958# 4.64e-21
C2363 XM1/a_n158_10170# XM2/a_n100_n142323# 6.96e-20
C2364 XM1/a_100_n142046# XM2/a_n100_n297847# 0.005074f
C2365 XM3/a_n100_n42455# XM4/a_n100_n42455# 0.009521f
C2366 XM2/a_100_n144862# XM3/a_n100_61145# 0.010147f
C2367 XM1/a_n100_n175171# XM2/a_100_n329382# 1.45e-19
C2368 XM2/a_n158_n255574# XM3/a_n100_n49707# 1.45e-19
C2369 XM1/a_n100_n60291# XM2/a_n158_n216034# 0.005074f
C2370 XM1/a_n158_126486# XM2/a_n100_n26339# 7.26e-20
C2371 XM1/a_n158_163822# XM2/a_n158_8026# 4.64e-21
C2372 XM4/a_n100_122269# m1_1634_n2388# 0.072015f
C2373 XM4/w_n358_n132787# XM3/a_n100_n26915# 0.009186f
C2374 XM4/a_100_n12314# m1_1634_n2388# 6.1e-20
C2375 XM1/a_n100_122081# XM2/a_n100_n31611# 7.77e-20
C2376 XM2/a_100_n187038# XM3/a_n100_18669# 0.010147f
C2377 XM1/a_n158_n179382# XM2/a_n100_n334751# 7.26e-20
C2378 XM4/w_n358_n132787# XM4/a_n100_n85967# -0.004445f
C2379 XM3/a_n158_n56862# m1_1634_n2388# 6.1e-20
C2380 XM1/a_n100_40229# XM4/w_n358_n132787# 0.014345f
C2381 XM4/a_100_19802# m1_1634_n2388# 6.1e-20
C2382 XM1/a_n100_21# XM2/a_100_n152770# 7.26e-20
C2383 XM2/a_n100_n250399# XM3/a_n158_n43394# 0.005074f
C2384 XM1/a_n100_n167991# XM2/a_n158_n321474# 0.005074f
C2385 XM1/a_n100_n66035# XM4/w_n358_n132787# 0.013462f
C2386 XM4/w_n358_n132787# XM3/a_n100_69433# 0.009643f
C2387 XM2/a_n100_n147595# m1_1634_n2388# 7.61e-19
C2388 XM1/a_n100_n57419# XM2/a_100_n210762# 7.26e-20
C2389 XM1/a_100_79098# XM3/a_n100_129521# 2.85e-20
C2390 XM2/a_n158_n329382# XM3/a_n100_n125335# 7.26e-20
C2391 XM1/a_100_n107582# m1_1634_n2388# 4.86e-19
C2392 XM4/w_n358_n132787# XM2/a_100_n213398# 0.105544f
C2393 XM2/a_n158_n200218# XM3/a_n158_4262# 4.64e-21
C2394 XM2/a_100_n332018# m1_1634_n2388# 0.017213f
C2395 XM3/a_n100_n62139# XM4/a_n100_n62139# 0.009521f
C2396 XM4/w_n358_n132787# XM3/a_n100_14525# 0.009186f
C2397 XM1/a_n100_n4287# XM2/a_100_n158042# 1.45e-19
C2398 XM1/a_n158_n139174# XM3/a_n100_n87003# 1.94e-20
C2399 XM4/a_n100_82901# m1_1634_n2388# 0.072015f
C2400 XM1/a_n100_22997# XM3/a_n100_74613# 4.37e-19
C2401 XM2/a_100_n284570# XM3/a_n158_n78618# 0.077916f
C2402 XM4/w_n358_n132787# XM3/a_n100_n66283# 0.009186f
C2403 XM4/a_100_n51682# m1_1634_n2388# 6.1e-20
C2404 XM1/a_100_n34346# XM2/a_100_n187038# 4.64e-21
C2405 XM3/a_n100_22813# XM4/a_n100_22813# 0.009521f
C2406 XM2/a_100_n326746# XM3/a_n100_n120155# 0.005074f
C2407 XM1/a_100_n83170# XM2/a_n158_n237122# 0.116862f
C2408 XM1/a_100_n67374# XM4/w_n358_n132787# 0.048442f
C2409 XM1/a_n158_107818# XM2/a_n100_n44791# 7.26e-20
C2410 XM1/a_100_54686# XM3/a_n100_106729# 2.85e-20
C2411 XM4/w_n358_n132787# XM4/a_n100_n125335# -0.004445f
C2412 XM1/a_100_n65938# XM3/a_n100_n14483# 4.35e-20
C2413 XM2/a_100_n173858# XM3/a_n100_33173# 0.005074f
C2414 XM3/a_n158_n96230# m1_1634_n2388# 6.1e-20
C2415 XM1/a_100_n58758# XM2/a_n158_n213398# 0.116862f
C2416 XM1/a_n100_31613# XM2/a_n158_n123774# 0.005074f
C2417 XM1/a_100_n176510# XM2/a_n100_n329479# 0.005074f
C2418 XM1/a_n100_n89011# XM2/a_100_n242394# 7.26e-20
C2419 XM2/a_n158_n237122# XM3/a_n100_n32095# 1.45e-19
C2420 XM1/a_n100_10073# XM3/a_n158_62278# 4.32e-20
C2421 XM4/w_n358_n132787# XM1/a_100_n163586# 0.054609f
C2422 XM1/a_100_107818# XM2/a_100_n47330# 4.64e-21
C2423 XM1/a_n100_27305# XM2/a_n158_n126410# 0.010147f
C2424 XM2/a_n100_n176591# XM4/a_100_30162# 2.56e-20
C2425 XM1/a_n100_n48803# XM3/a_n158_2190# 2.85e-20
C2426 XM3/a_n100_52857# m1_1634_n2388# 0.072015f
C2427 XM1/a_n158_106382# XM2/a_n158_n47330# 9.28e-21
C2428 XM3/a_n100_n81823# XM4/a_n100_n81823# 0.009521f
C2429 XM1/a_n100_n28699# XM2/a_100_n184402# 7.26e-20
C2430 XM1/a_100_67610# XM3/a_n100_118125# 2.85e-20
C2431 XM1/a_n158_n116198# XM2/a_n100_n271487# 7.26e-20
C2432 XM4/w_n358_n132787# XM3/a_n100_2093# 0.009186f
C2433 XM4/w_n358_n132787# XM2/a_n100_n152867# 0.025738f
C2434 XM1/a_n100_28741# XM2/a_100_n123774# 7.26e-20
C2435 XM2/a_n100_n271487# m1_1634_n2388# 0.002452f
C2436 XM1/a_n158_n63066# XM2/a_n100_n216131# 7.26e-20
C2437 XM4/a_n100_43533# m1_1634_n2388# 0.072015f
C2438 XM4/w_n358_n132787# XM3/a_n100_n105651# 0.009186f
C2439 XM4/a_100_n91050# m1_1634_n2388# 6.1e-20
C2440 XM2/a_n158_n115866# XM3/a_n100_89117# 1.45e-19
C2441 XM1/a_n158_54686# XM3/a_n100_106729# 1.94e-20
C2442 XM1/a_n100_44537# m1_1634_n2388# 1.3e-19
C2443 XM4/w_n358_n132787# XM3/a_n158_94394# 0.032295f
C2444 XM4/w_n358_n132787# XM2/a_100_n337290# 0.103341f
C2445 XM1/a_n100_n48803# XM4/w_n358_n132787# 0.01363f
C2446 XM1/a_100_n98966# XM2/a_n158_n252938# 0.116862f
C2447 XM3/a_n100_4165# XM4/a_n100_4165# 0.009521f
C2448 XM4/w_n358_n132787# XM3/a_n158_39486# 0.032295f
C2449 XM2/a_n158_n158042# XM3/a_n100_46641# 7.26e-20
C2450 XM1/a_n100_n31571# XM2/a_n158_n184402# 0.005074f
C2451 XM2/a_100_n110594# XM3/a_n158_94394# 0.077916f
C2452 XM4/w_n358_n132787# XM1/a_n100_n165119# 0.013385f
C2453 XM2/a_100_n84234# XM3/a_n100_122269# 0.005074f
C2454 XM2/a_n158_n84234# XM3/a_n158_122366# 4.64e-21
C2455 XM2/a_100_n266118# XM3/a_n158_n61006# 0.077916f
C2456 XM1/a_n158_n38654# XM2/a_n158_n192310# 9.28e-21
C2457 XM1/a_n100_n61727# XM2/a_n158_n216034# 0.010147f
C2458 XM2/a_100_n308294# XM3/a_n100_n102543# 0.010147f
C2459 XM4/w_n358_n132787# XM3/a_n158_n41322# 0.032295f
C2460 XM4/a_n100_n27951# m1_1634_n2388# 0.072015f
C2461 XM1/a_100_n147790# XM2/a_n100_n303119# 0.005074f
C2462 XM2/a_100_n152770# XM3/a_n158_51918# 0.067011f
C2463 XM2/a_n100_n305755# XM3/a_n158_n101410# 0.005074f
C2464 XM1/a_100_n127686# XM3/a_n100_n75607# 2.85e-20
C2465 XM1/a_n100_n71779# m1_1634_n2388# 9.35e-20
C2466 XM3/a_n100_n101507# XM4/a_n100_n101507# 0.009521f
C2467 XM1/a_100_76226# XM2/a_n158_n76326# 0.014823f
C2468 XM2/a_n158_n218670# XM3/a_n100_n14483# 7.26e-20
C2469 XM1/a_100_n73118# m1_1634_n2388# 5.46e-19
C2470 XM2/a_100_n194946# XM3/a_n158_9442# 0.037801f
C2471 XM4/w_n358_n132787# XM2/a_n158_n89506# 0.107093f
C2472 XM1/a_n100_12945# XM2/a_n158_n142226# 0.005074f
C2473 XM1/a_n100_n27263# XM3/a_n158_23946# 2.67e-20
C2474 XM2/a_n158_n13062# XM1/a_100_139410# 0.007033f
C2475 XM2/a_n100_n13159# XM1/a_n158_139410# 7.26e-20
C2476 XM1/a_100_57558# XM2/a_n158_n97414# 0.100115f
C2477 XM2/a_n158_n208126# m1_1634_n2388# 2.36e-21
C2478 XM2/a_n158_n303022# XM3/a_n158_n96230# 4.64e-21
C2479 XM1/a_n100_n70343# XM4/w_n358_n132787# 0.013608f
C2480 XM1/a_n100_160853# XM2/a_100_5390# 7.26e-20
C2481 XM1/a_n100_43101# XM3/a_n100_94297# 0.001134f
C2482 XM4/w_n358_n132787# XM2/a_n100_n276759# 0.026749f
C2483 XM2/a_100_n216034# XM3/a_n100_n9303# 0.005074f
C2484 XM3/a_n158_77818# m1_1634_n2388# 6.1e-20
C2485 XM3/a_n158_110970# m1_1634_n2388# 6.1e-20
C2486 XM4/w_n358_n132787# XM4/a_n100_98441# -0.004445f
C2487 XM1/a_n158_47506# XM2/a_n100_n108055# 7.26e-20
C2488 XM2/a_n158_n144862# XM3/a_n100_61145# 1.45e-19
C2489 XM1/a_100_n142046# XM2/a_100_n295114# 4.64e-21
C2490 XM1/a_n100_n83267# XM3/a_n100_n32095# 7.68e-19
C2491 XM3/a_n100_n8267# m1_1634_n2388# 0.072015f
C2492 XM1/a_n100_n175171# XM2/a_n158_n329382# 0.010147f
C2493 XM3/a_n158_22910# m1_1634_n2388# 6.1e-20
C2494 XM1/a_100_10170# XM4/w_n358_n132787# 0.054514f
C2495 XM4/w_n358_n132787# XM3/a_n158_n80690# 0.035272f
C2496 XM4/a_n100_n67319# m1_1634_n2388# 0.072015f
C2497 XM1/a_n100_n155067# XM3/a_n158_n104518# 2.85e-20
C2498 XM2/a_n158_n187038# XM3/a_n100_18669# 1.45e-19
C2499 XM1/a_n100_150801# XM2/a_n158_n5154# 0.003292f
C2500 XM2/a_100_n139590# XM3/a_n158_66422# 0.077916f
C2501 XM1/a_100_n75990# XM3/a_n158_n24746# 0.00544f
C2502 XM3/a_n100_n121191# XM4/a_n100_n121191# 0.009521f
C2503 XM1/a_n100_21# XM2/a_n158_n152770# 0.005074f
C2504 XM1/a_n158_n159278# XM3/a_n100_n107723# 1.94e-20
C2505 XM2/a_100_n247666# XM3/a_n158_n43394# 0.026507f
C2506 XM1/a_n100_n167991# XM2/a_n100_n321571# 0.004872f
C2507 XM2/a_n100_n253035# XM4/a_100_n48574# 2.56e-20
C2508 XM2/a_100_n181766# XM3/a_n158_23946# 0.077916f
C2509 XM2/a_100_n289842# XM3/a_n100_n84931# 0.010147f
C2510 XM1/a_n158_58994# XM3/a_n100_110873# 1.94e-20
C2511 XM3/a_n100_75649# XM4/a_n100_75649# 0.009521f
C2512 XM1/a_100_n121942# XM3/a_n100_n70427# 2.85e-20
C2513 XM2/a_100_n144862# m1_1634_n2388# 0.025819f
C2514 XM1/a_100_n152098# XM3/a_n158_n101410# 0.001512f
C2515 XM1/a_n100_n57419# XM2/a_n158_n210762# 0.005074f
C2516 XM3/a_n100_122269# XM4/a_n100_122269# 0.009521f
C2517 XM1/a_n100_24433# XM3/a_n100_75649# 4.67e-19
C2518 XM4/w_n358_n132787# XM2/a_n158_n213398# 0.105837f
C2519 XM2/a_n100_n200315# XM3/a_n158_4262# 0.005074f
C2520 XM4/w_n358_n132787# XM4/a_n100_59073# -0.004445f
C2521 XM3/a_n100_n47635# m1_1634_n2388# 0.072015f
C2522 XM1/a_100_n35782# XM3/a_n100_16597# 6.97e-21
C2523 XM1/a_n100_n4287# XM2/a_n158_n158042# 0.010147f
C2524 XM1/a_n100_n152195# XM3/a_n158_n100374# 2.85e-20
C2525 XM1/a_100_38890# XM4/w_n358_n132787# 0.048442f
C2526 XM1/a_n100_n173735# XM2/a_100_n329382# 7.26e-20
C2527 XM4/w_n358_n132787# XM3/a_n158_n120058# 0.038462f
C2528 XM4/a_n100_n106687# m1_1634_n2388# 0.072015f
C2529 XM1/a_100_n34346# XM2/a_n158_n187038# 0.028454f
C2530 XM1/a_n100_155109# XM2/a_n158_2754# 0.005074f
C2531 XM4/w_n358_n132787# XM3/a_n158_108898# 0.032295f
C2532 XM1/a_100_n12806# XM3/a_n100_39389# 2.85e-20
C2533 XM1/a_n100_50281# m1_1634_n2388# 9.55e-20
C2534 XM2/a_n158_n326746# XM3/a_n100_n120155# 7.26e-20
C2535 XM1/a_n158_n149226# XM3/a_n100_n97363# 1.94e-20
C2536 XM1/a_n158_n35782# XM3/a_n100_15561# 3.89e-20
C2537 XM2/a_100_26478# XM1/a_100_179618# 4.64e-21
C2538 XM2/a_100_n10426# XM1/a_100_142282# 4.64e-21
C2539 XM2/a_n158_n13062# XM1/a_n158_140846# 9.28e-21
C2540 XM1/a_n100_103413# XM2/a_n100_n52699# 0.004582f
C2541 XM2/a_n158_n173858# XM3/a_n100_33173# 7.26e-20
C2542 XM1/a_n100_n152195# XM2/a_100_n305658# 7.26e-20
C2543 XM1/a_n100_n103371# XM2/a_100_n258210# 7.26e-20
C2544 XM1/a_n100_n89011# XM2/a_n158_n242394# 0.005074f
C2545 XM2/a_100_n100050# XM3/a_n158_104754# 0.077916f
C2546 XM1/a_n158_14478# XM3/a_n100_65289# 1.94e-20
C2547 XM1/a_100_n183690# XM2/a_n158_n337290# 0.11685f
C2548 XM4/w_n358_n132787# XM4/a_n100_n12411# -0.004445f
C2549 XM1/a_n100_100541# XM4/w_n358_n132787# 0.012279f
C2550 XM1/a_n100_n10031# XM4/w_n358_n132787# 0.013065f
C2551 XM2/a_100_n168586# XM3/a_n158_38450# 0.015991f
C2552 XM1/a_100_172438# XM4/w_n358_n132787# 0.048442f
C2553 XM4/a_100_93358# m1_1634_n2388# 6.1e-20
C2554 XM1/a_n158_n5626# XM3/a_n100_45605# 2.34e-20
C2555 XM1/a_n100_2893# XM3/a_n158_55026# 2.85e-20
C2556 XM2/a_n100_n84331# m1_1634_n2388# 7.61e-19
C2557 XM4/w_n358_n132787# XM3/a_n100_88081# 0.009186f
C2558 XM1/a_100_13042# m1_1634_n2388# 6.67e-19
C2559 XM1/a_n158_n88914# XM3/a_n100_n38311# 1.94e-20
C2560 XM4/w_n358_n132787# XM4/a_n100_19705# -0.004445f
C2561 XM3/a_n100_n87003# m1_1634_n2388# 0.072015f
C2562 XM1/a_n100_n28699# XM2/a_n158_n184402# 0.005074f
C2563 XM1/a_n100_28741# XM2/a_n158_n123774# 0.005074f
C2564 XM4/w_n358_n132787# XM2/a_100_n150134# 0.106245f
C2565 XM1/a_n100_58897# XM4/w_n358_n132787# 0.01363f
C2566 XM1/a_n100_n129219# m1_1634_n2388# 1.11e-19
C2567 XM2/a_100_n268754# m1_1634_n2388# 0.017213f
C2568 XM4/w_n358_n132787# XM3/a_n100_33173# 0.009135f
C2569 XM2/a_100_n271390# XM3/a_n100_n67319# 0.005074f
C2570 XM1/a_100_100638# XM2/a_n100_n55335# 0.005074f
C2571 XM4/w_n358_n132787# XM2/a_n158_n337290# 0.101988f
C2572 XM1/a_n100_57461# XM2/a_100_n97414# 7.26e-20
C2573 XM1/a_100_n116198# XM3/a_n100_n64211# 0.001288f
C2574 XM1/a_n100_n106243# XM3/a_n100_n55923# 0.001041f
C2575 XM1/a_n158_n67374# XM3/a_n100_n15519# 1.94e-20
C2576 XM2/a_100_n205490# XM3/a_n158_118# 0.077916f
C2577 XM1/a_n100_170905# XM2/a_n158_15934# 0.005074f
C2578 XM1/a_n158_89150# XM2/a_n100_n65879# 7.26e-20
C2579 XM2/a_n100_n158139# XM3/a_n100_46641# 0.004501f
C2580 XM1/a_100_n73118# XM3/a_n100_n22771# 0.001222f
C2581 XM1/a_n100_n38751# m1_1634_n2388# 2.01e-19
C2582 XM4/w_n358_n132787# XM4/a_n100_n51779# -0.004445f
C2583 XM3/a_n158_n22674# m1_1634_n2388# 6.1e-20
C2584 XM1/a_n100_76129# XM2/a_100_n76326# 7.26e-20
C2585 XM2/a_n100_n84331# XM3/a_n158_122366# 0.005074f
C2586 XM2/a_n158_n84234# XM3/a_n100_122269# 7.26e-20
C2587 XM3/a_n100_105693# XM4/a_n100_105693# 0.009521f
C2588 XM2/a_n100_n121235# XM4/a_100_82998# 2.56e-20
C2589 XM1/a_n100_n130655# XM3/a_n158_n78618# 2.85e-20
C2590 XM1/a_n100_21561# XM4/w_n358_n132787# 0.01363f
C2591 XM4/a_100_53990# m1_1634_n2388# 6.1e-20
C2592 XM2/a_n158_n39422# XM4/w_n358_n132787# 0.107093f
C2593 XM1/a_n158_23094# XM2/a_n158_n131682# 9.28e-21
C2594 XM2/a_n158_n308294# XM3/a_n100_n102543# 1.45e-19
C2595 XM2/a_n158_n152770# XM3/a_n158_51918# 4.64e-21
C2596 XM1/a_100_96330# XM2/a_n158_n57874# 0.116862f
C2597 XM1/a_100_n147790# XM2/a_100_n300386# 4.64e-21
C2598 XM1/a_n100_n180915# XM4/w_n358_n132787# 0.013401f
C2599 XM4/a_100_3226# m1_1634_n2388# 6.1e-20
C2600 XM1/a_100_76226# XM2/a_n100_n76423# 0.005074f
C2601 XM3/a_n100_n126371# m1_1634_n2388# 0.072015f
C2602 XM1/a_n158_94894# XM2/a_n100_n57971# 7.26e-20
C2603 XM3/a_n100_71505# m1_1634_n2388# 0.072015f
C2604 XM2/a_n158_n194946# XM3/a_n158_9442# 4.64e-21
C2605 XM1/a_100_n21422# XM2/a_100_n176494# 4.64e-21
C2606 XM4/w_n358_n132787# XM2/a_n100_n89603# 0.025738f
C2607 XM1/a_100_n133430# XM3/a_n100_n81823# 2.85e-20
C2608 XM1/a_100_n83170# XM4/w_n358_n132787# 0.048442f
C2609 XM1/a_100_57558# XM2/a_n100_n97511# 0.005074f
C2610 XM1/a_100_n139174# XM3/a_n158_n87942# 0.00544f
C2611 XM2/a_n100_n208223# m1_1634_n2388# 8e-19
C2612 XM2/a_n100_n303119# XM3/a_n158_n96230# 0.005074f
C2613 XM1/a_n158_n131994# XM2/a_n158_n284570# 4.64e-21
C2614 XM3/a_n100_16597# m1_1634_n2388# 0.072015f
C2615 XM1/a_100_n110454# XM3/a_n158_n58934# 0.00544f
C2616 XM4/a_n100_117089# m1_1634_n2388# 0.072015f
C2617 XM4/w_n358_n132787# XM2/a_100_n274026# 0.103341f
C2618 XM4/w_n358_n132787# XM3/a_n100_n32095# 0.009036f
C2619 XM4/a_100_n17494# m1_1634_n2388# 6.1e-20
C2620 XM2/a_n158_n216034# XM3/a_n100_n9303# 7.26e-20
C2621 XM1/a_n100_4329# XM2/a_100_n150134# 1.45e-19
C2622 XM3/a_n100_110873# m1_1634_n2388# 0.072015f
C2623 XM1/a_100_n142046# XM2/a_n158_n295114# 0.065063f
C2624 XM4/w_n358_n132787# XM4/a_n100_n91147# -0.004445f
C2625 XM3/a_n158_n62042# m1_1634_n2388# 6.1e-20
C2626 XM1/a_n100_n45931# XM3/a_n100_5201# 2.09e-19
C2627 XM1/a_100_158078# XM2/a_n100_5293# 0.005074f
C2628 XM4/w_n358_n132787# XM3/a_n158_58134# 0.032295f
C2629 XM1/a_n100_n60291# XM2/a_100_n213398# 7.26e-20
C2630 XM1/a_100_46070# XM4/w_n358_n132787# 0.048442f
C2631 XM4/a_100_14622# m1_1634_n2388# 6.1e-20
C2632 XM2/a_n158_8026# XM4/w_n358_n132787# 0.107093f
C2633 XM1/a_100_n44398# XM3/a_n100_6237# 0.001477f
C2634 XM3/a_n100_43533# XM4/a_n100_43533# 0.009521f
C2635 XM4/w_n358_n132787# XM1/a_n100_137877# 0.01219f
C2636 XM2/a_100_n337290# XM3/a_n158_n131454# 0.077916f
C2637 XM1/a_100_n129122# XM4/w_n358_n132787# 0.054609f
C2638 XM1/a_n158_n179382# XM2/a_n158_n332018# 4.64e-21
C2639 XM4/w_n358_n132787# XM1/a_100_n137738# 0.048442f
C2640 XM1/a_n158_n131994# XM3/a_n100_n79751# 1.94e-20
C2641 XM1/a_100_n80298# XM3/a_n100_n28987# 5.71e-20
C2642 XM1/a_100_n53014# m1_1634_n2388# 2.43e-19
C2643 XM2/a_n158_n247666# XM3/a_n158_n43394# 4.64e-21
C2644 XM1/a_n158_n73118# XM3/a_n158_n22674# 1.14e-21
C2645 XM2/a_n158_n289842# XM3/a_n100_n84931# 1.45e-19
C2646 XM1/a_100_119306# XM2/a_n100_n34247# 0.005074f
C2647 XM4/a_n100_77721# m1_1634_n2388# 0.072015f
C2648 XM4/w_n358_n132787# XM3/a_n100_n71463# 0.009186f
C2649 XM4/a_100_n56862# m1_1634_n2388# 6.1e-20
C2650 XM4/w_n358_n132787# XM2/a_n100_n213495# 0.023697f
C2651 XM1/a_100_79098# XM3/a_n158_130654# 0.00544f
C2652 XM2/a_100_n245030# XM3/a_n158_n38214# 0.037411f
C2653 XM3/a_n158_96466# m1_1634_n2388# 6.1e-20
C2654 XM4/w_n358_n132787# XM4/a_n100_n130515# -0.004445f
C2655 XM2/a_n100_n332115# m1_1634_n2388# 7.85e-19
C2656 XM3/a_n158_n101410# m1_1634_n2388# 6.1e-20
C2657 XM2/a_n100_n250399# XM4/a_100_n43394# 2.56e-20
C2658 XM1/a_n100_n41623# XM3/a_n158_9442# 6.54e-19
C2659 XM1/a_n100_n14339# XM3/a_n158_36378# 2.85e-20
C2660 XM1/a_n100_15817# XM3/a_n158_66422# 2.85e-20
C2661 XM1/a_n100_n173735# XM2/a_n158_n329382# 0.005074f
C2662 XM1/a_n158_165258# XM2/a_n158_10662# 9.28e-21
C2663 XM1/a_n100_37357# XM2/a_100_n118502# 7.26e-20
C2664 XM1/a_n158_25966# XM3/a_n158_77818# 1.14e-21
C2665 XM1/a_100_n34346# XM2/a_n100_n187135# 0.005074f
C2666 XM3/a_n158_41558# m1_1634_n2388# 6.1e-20
C2667 XM4/w_n358_n132787# XM3/a_n100_108801# 0.008986f
C2668 pcbias sw_b 0.0465f
C2669 pbias sw_bn 0.001128f
C2670 XM1/a_n100_31613# XM2/a_100_n121138# 7.26e-20
C2671 XM1/a_n100_n152195# XM2/a_n158_n305658# 0.005074f
C2672 XM1/a_n100_n103371# XM2/a_n158_n258210# 0.005074f
C2673 XM4/w_n358_n132787# XM3/a_n158_n7134# 0.032295f
C2674 XM1/a_n158_n136302# XM2/a_n158_n289842# 4.64e-21
C2675 XM2/a_100_n100050# XM3/a_n100_104657# 0.005159f
C2676 XM1/a_100_n183690# XM2/a_n100_n337387# 4.68e-21
C2677 XM1/a_n100_n117731# m1_1634_n2388# 7.34e-20
C2678 XM1/a_n100_n80395# XM3/a_n158_n29926# 2.11e-20
C2679 XM1/a_100_8734# XM3/a_n100_60109# 5.71e-20
C2680 XM1/a_n100_n22955# XM3/a_n158_28090# 0.001324f
C2681 XM2/a_n158_n168586# XM3/a_n158_38450# 4.64e-21
C2682 XM4/a_n100_38353# m1_1634_n2388# 0.072015f
C2683 XM2/a_100_n318838# XM3/a_n158_n113842# 0.077916f
C2684 XM4/w_n358_n132787# XM3/a_n100_n110831# 0.009186f
C2685 XM4/a_100_n96230# m1_1634_n2388# 6.1e-20
C2686 XM1/a_n100_104849# XM2/a_n100_n47427# 0.005548f
C2687 XM2/a_n100_n21067# XM1/a_100_132230# 0.005074f
C2688 XM1/a_n100_74693# XM3/a_n158_126510# 2.85e-20
C2689 XM2/a_100_n81598# m1_1634_n2388# 0.023671f
C2690 XM1/a_n100_48845# m1_1634_n2388# 1.1e-19
C2691 XM1/a_n158_n173638# XM3/a_n100_n123263# 1.94e-20
C2692 XM1/a_100_n129122# XM3/a_n100_n77679# 4.7e-20
C2693 XM1/a_100_n88914# XM3/a_n100_n37275# 2.85e-20
C2694 XM1/a_n158_n22858# XM3/a_n100_29029# 1.94e-20
C2695 XM1/a_100_165258# XM4/w_n358_n132787# 0.048442f
C2696 XM1/a_n158_n109018# XM3/a_n100_n57995# 1.94e-20
C2697 XM1/a_n158_71918# XM3/a_n100_123305# 3.89e-20
C2698 XM4/w_n358_n132787# XM2/a_n158_n150134# 0.107093f
C2699 XM1/a_n158_n116198# XM2/a_n158_n268754# 4.64e-21
C2700 XM1/a_n100_n89011# m1_1634_n2388# 9.61e-20
C2701 XM1/a_n158_n11370# XM3/a_n100_39389# 1.94e-20
C2702 XM1/a_n100_24433# XM2/a_100_n129046# 7.26e-20
C2703 XM2/a_n158_n271390# XM3/a_n100_n67319# 7.26e-20
C2704 XM4/w_n358_n132787# XM2/a_n100_n337387# 0.02288f
C2705 XM2/a_n100_n55335# XM4/w_n358_n132787# 0.012279f
C2706 XM1/a_n100_57461# XM2/a_n158_n97414# 0.005074f
C2707 XM1/a_n100_22997# XM2/a_100_n131682# 9.05e-20
C2708 XM4/w_n358_n132787# XM3/a_n158_n46502# 0.033396f
C2709 XM4/a_n100_n33131# m1_1634_n2388# 0.072015f
C2710 XM2/a_100_n226578# XM3/a_n158_n20602# 0.077916f
C2711 XM1/a_100_5862# m1_1634_n2388# 9.71e-19
C2712 XM1/a_n158_n117634# XM3/a_n100_n66283# 3.89e-20
C2713 XM2/a_100_n268754# XM3/a_n100_n62139# 0.005074f
C2714 XM1/a_n100_76129# XM2/a_n158_n76326# 0.005074f
C2715 XM1/a_100_163822# XM2/a_n158_10662# 0.074021f
C2716 XM2/a_n100_n152867# XM3/a_n158_51918# 0.005074f
C2717 XM1/a_n158_97766# XM2/a_n100_n55335# 7.26e-20
C2718 XM1/a_100_n147790# XM2/a_n158_n300386# 0.019107f
C2719 XM1/a_n100_165161# XM2/a_100_10662# 1.45e-19
C2720 XM1/a_100_n136302# XM4/w_n358_n132787# 0.049932f
C2721 XM1/a_n100_n114859# XM3/a_n158_n63078# 2.55e-20
C2722 XM2/a_n100_n118599# XM4/a_100_88178# 2.56e-20
C2723 XM1/a_100_n150662# XM3/a_n100_n98399# 0.001158f
C2724 XM1/a_100_n119070# XM2/a_n100_n271487# 8.32e-19
C2725 XM2/a_n100_n195043# XM3/a_n158_9442# 0.005074f
C2726 XM1/a_100_n21422# XM2/a_n158_n176494# 0.090379f
C2727 XM4/w_n358_n132787# XM2/a_100_n86870# 0.10657f
C2728 XM4/w_n358_n132787# XM4/a_n100_93261# -0.004445f
C2729 XM1/a_n100_12945# XM2/a_100_n139590# 7.26e-20
C2730 XM3/a_n100_n13447# m1_1634_n2388# 0.072015f
C2731 XM2/a_100_n205490# m1_1634_n2388# 0.017213f
C2732 XM4/w_n358_n132787# XM3/a_n100_51821# 0.007942f
C2733 XM2/a_100_n300386# XM3/a_n158_n96230# 0.015212f
C2734 XM1/a_n158_n131994# XM2/a_n100_n284667# 7.26e-20
C2735 XM3/a_n100_96369# XM4/a_n100_96369# 0.009521f
C2736 XM2/a_n100_n305755# XM4/a_100_n101410# 2.56e-20
C2737 XM4/w_n358_n132787# XM2/a_n158_n274026# 0.101988f
C2738 XM1/a_n158_n96094# XM2/a_n158_n250302# 9.28e-21
C2739 XM3/a_n100_11417# XM4/a_n100_11417# 0.009521f
C2740 XM4/w_n358_n132787# XM3/a_n158_n85870# 0.037964f
C2741 XM4/a_n100_n72499# m1_1634_n2388# 0.072015f
C2742 XM1/a_n158_47506# XM2/a_n158_n105322# 4.64e-21
C2743 XM1/a_n100_4329# XM2/a_n158_n150134# 0.010147f
C2744 XM1/a_n100_n179479# XM4/w_n358_n132787# 0.01363f
C2745 XM1/a_100_n142046# XM2/a_n100_n295211# 0.005074f
C2746 XM1/a_n100_n60291# XM2/a_n158_n213398# 0.005074f
C2747 XM1/a_n100_n81831# m1_1634_n2388# 1.3e-19
C2748 XM1/a_100_n50142# XM3/a_n100_2093# 2.85e-20
C2749 XM4/w_n358_n132787# XM3/a_n158_3226# 0.032295f
C2750 XM1/a_n100_n20083# XM3/a_n158_32234# 2.85e-20
C2751 XM1/a_n158_64738# XM2/a_n158_n89506# 9.28e-21
C2752 XM4/a_100_127546# m1_1634_n2388# 6.1e-20
C2753 XM1/a_n158_n179382# XM2/a_n100_n332115# 7.26e-20
C2754 XM2/a_100_n250302# XM3/a_n100_n44527# 0.010147f
C2755 XM4/w_n358_n132787# XM4/a_n100_53893# -0.004445f
C2756 XM2/a_n100_n247763# XM3/a_n158_n43394# 0.005074f
C2757 XM3/a_n100_90153# m1_1634_n2388# 0.072015f
C2758 XM1/a_100_n167894# XM4/w_n358_n132787# 0.04904f
C2759 XM1/a_100_n130558# XM3/a_n100_n78715# 2.85e-20
C2760 XM3/a_n100_n52815# m1_1634_n2388# 0.072015f
C2761 XM1/a_n100_n24391# XM3/a_n158_26018# 3.44e-21
C2762 XM1/a_100_31710# XM3/a_n158_82998# 0.00544f
C2763 XM2/a_n100_n144959# m1_1634_n2388# 7.61e-19
C2764 XM4/w_n358_n132787# XM3/a_n158_n125238# 0.038462f
C2765 XM4/a_n100_n111867# m1_1634_n2388# 0.072015f
C2766 XM4/w_n358_n132787# XM4/a_n100_3129# -0.004445f
C2767 XM3/a_n100_35245# m1_1634_n2388# 0.072015f
C2768 XM3/a_n100_n8267# XM4/a_n100_n8267# 0.009521f
C2769 XM4/w_n358_n132787# XM2/a_100_n210762# 0.103341f
C2770 XM1/a_100_79098# XM3/a_n100_130557# 4.23e-20
C2771 XM1/a_n100_60333# m1_1634_n2388# 9.43e-20
C2772 XM1/a_100_n154970# m1_1634_n2388# 0.003275f
C2773 XM2/a_n158_n245030# XM3/a_n158_n38214# 4.64e-21
C2774 XM1/a_n158_n14242# XM3/a_n100_37317# 1.94e-20
C2775 XM2/a_100_n329382# m1_1634_n2388# 0.023368f
C2776 XM1/a_n100_n43059# XM3/a_n158_9442# 2.82e-20
C2777 XM1/a_100_71918# m1_1634_n2388# 0.001092f
C2778 XM2/a_100_n129046# XM3/a_n100_75649# 0.005074f
C2779 XM1/a_n100_37357# XM2/a_n158_n118502# 0.005074f
C2780 XM4/w_n358_n132787# XM3/a_n158_76782# 0.032295f
C2781 XM4/w_n358_n132787# XM4/a_n100_n17591# -0.004445f
C2782 XM1/a_n158_n182254# pbias 0.011406f
C2783 XM2/a_100_n324110# XM3/a_n100_n120155# 0.005074f
C2784 XM2/a_100_n171222# XM3/a_n100_33173# 0.005074f
C2785 XM1/a_100_n7062# XM3/a_n100_44569# 2.85e-20
C2786 XM1/a_100_n5626# XM4/w_n358_n132787# 0.055087f
C2787 XM4/w_n358_n132787# XM3/a_n158_21874# 0.032295f
C2788 XM1/a_100_169566# XM4/w_n358_n132787# 0.048442f
C2789 XM4/a_100_88178# m1_1634_n2388# 6.1e-20
C2790 XM1/a_n100_31613# XM2/a_n158_n121138# 0.005074f
C2791 XM1/a_n100_8637# XM3/a_n100_61145# 0.001119f
C2792 XM1/a_n100_n152195# XM2/a_n100_n305755# 0.003018f
C2793 XM1/a_n158_n136302# XM2/a_n100_n289939# 4.89e-20
C2794 XM2/a_n158_n100050# XM3/a_n100_104657# 7.56e-20
C2795 XM1/a_n100_n70343# XM3/a_n158_n18530# 2.85e-20
C2796 XM4/w_n358_n132787# XM4/a_n100_14525# -0.004445f
C2797 XM1/a_n100_100541# XM2/a_n158_n55238# 0.005074f
C2798 XM3/a_n100_n92183# m1_1634_n2388# 0.072015f
C2799 XM2/a_n100_n168683# XM3/a_n158_38450# 0.005074f
C2800 XM2/a_n100_n173955# XM4/a_100_30162# 2.56e-20
C2801 XM1/a_100_n37218# XM3/a_n100_14525# 2.85e-20
C2802 XM3/a_n100_n27951# XM4/a_n100_n27951# 0.009521f
C2803 XM2/a_n158_n81598# m1_1634_n2388# 2.36e-21
C2804 XM1/a_100_71918# XM3/a_n158_122366# 1.91e-19
C2805 XM1/a_n158_28838# XM2/a_n158_n126410# 4.64e-21
C2806 XM2/a_100_n231850# XM3/a_n100_n26915# 0.010147f
C2807 XM1/a_n100_n28699# XM2/a_100_n181766# 7.26e-20
C2808 XM1/a_n100_n77523# XM3/a_n100_n25879# 6.89e-19
C2809 XM1/a_100_67610# XM3/a_n100_119161# 2.85e-20
C2810 XM4/w_n358_n132787# XM2/a_n100_n150231# 0.025056f
C2811 XM1/a_n158_n116198# XM2/a_n100_n268851# 7.26e-20
C2812 XM1/a_n100_n28699# XM3/a_n100_23849# 5.98e-19
C2813 XM1/a_n100_101977# XM2/a_100_n52602# 1.45e-19
C2814 XM2/a_n100_n268851# m1_1634_n2388# 7.61e-19
C2815 XM1/a_n100_24433# XM2/a_n158_n129046# 0.005074f
C2816 XM1/a_100_n17114# XM3/a_n100_35245# 1.29e-20
C2817 XM2/a_100_n115866# XM3/a_n100_90153# 0.010147f
C2818 XM4/w_n358_n132787# XM2/a_100_n334654# 0.104215f
C2819 XM4/w_n358_n132787# XM4/a_n100_n56959# -0.004445f
C2820 XM3/a_n158_n27854# m1_1634_n2388# 6.1e-20
C2821 XM1/a_n100_25869# XM4/w_n358_n132787# 0.013098f
C2822 XM3/a_n158_60206# m1_1634_n2388# 6.1e-20
C2823 XM1/a_n100_n38751# XM3/a_n158_13586# 2.85e-20
C2824 XM4/a_100_48810# m1_1634_n2388# 6.1e-20
C2825 XM1/a_n100_22997# XM2/a_n158_n131682# 0.005563f
C2826 XM2/a_100_n158042# XM3/a_n100_47677# 0.010147f
C2827 XM2/a_n158_n268754# XM3/a_n100_n62139# 7.26e-20
C2828 XM3/a_n100_n131551# m1_1634_n2388# 0.072015f
C2829 XM2/a_n158_21206# XM1/a_n100_176649# 0.005074f
C2830 XM2/a_100_n81598# XM3/a_n100_122269# 0.004352f
C2831 XM1/a_n100_n140707# m1_1634_n2388# 8.61e-20
C2832 XM1/a_n100_126389# XM2/a_n158_n26242# 0.005074f
C2833 XM1/a_n158_171002# XM2/a_n158_18570# 4.64e-21
C2834 XM1/a_n158_n97530# XM2/a_n158_n252938# 4.64e-21
C2835 XM3/a_n100_64253# XM4/a_n100_64253# 0.009521f
C2836 XM1/a_n158_n157842# XM2/a_n158_n313566# 4.64e-21
C2837 XM1/a_100_n147790# XM2/a_n100_n300483# 0.005074f
C2838 XM1/a_n158_n134866# XM3/a_n100_n83895# 1.94e-20
C2839 XM3/a_n100_n47635# XM4/a_n100_n47635# 0.009521f
C2840 XM1/a_n100_n33007# XM3/a_n158_17730# 2.85e-20
C2841 XM1/a_100_96330# XM4/w_n358_n132787# 0.048442f
C2842 XM1/a_n158_17350# XM2/a_n158_n136954# 9.28e-21
C2843 XM4/a_n100_111909# m1_1634_n2388# 0.072015f
C2844 XM1/a_n100_56025# XM2/a_n100_n100147# 9.65e-19
C2845 XM1/a_n100_n90447# XM2/a_100_n245030# 1.45e-19
C2846 XM4/w_n358_n132787# XM3/a_n100_n37275# 0.009026f
C2847 XM4/a_100_n22674# m1_1634_n2388# 6.1e-20
C2848 XM1/a_100_n21422# XM2/a_n100_n176591# 0.005074f
C2849 XM4/w_n358_n132787# XM2/a_n158_n86870# 0.107093f
C2850 XM1/a_n100_12945# XM2/a_n158_n139590# 0.005074f
C2851 XM1/a_100_n167894# XM3/a_n100_n117047# 2.85e-20
C2852 XM4/w_n358_n132787# XM4/a_n100_n96327# -0.004445f
C2853 XM3/a_n158_n67222# m1_1634_n2388# 6.1e-20
C2854 XM1/a_100_n97530# XM2/a_100_n252938# 4.64e-21
C2855 XM2/a_n158_n300386# XM3/a_n158_n96230# 4.64e-21
C2856 XM4/w_n358_n132787# XM2/a_n100_n274123# 0.025142f
C2857 XM4/a_100_9442# m1_1634_n2388# 6.1e-20
C2858 XM2/a_100_n213398# XM3/a_n100_n9303# 0.005074f
C2859 XM2/a_n100_n7887# XM4/w_n358_n132787# 0.012279f
C2860 XM1/a_n158_129358# XM2/a_n158_n23606# 4.64e-21
C2861 XM1/a_n158_n133430# XM3/a_n100_n82859# 1.94e-20
C2862 XM3/a_n158_112006# m1_1634_n2388# 6.1e-20
C2863 XM1/a_n158_47506# XM2/a_n100_n105419# 7.26e-20
C2864 XM2/a_100_n144862# XM3/a_n100_62181# 0.005074f
C2865 XM1/a_100_43198# XM3/a_n100_94297# 2.85e-20
C2866 XM1/a_100_n166458# XM3/a_n158_n114878# 0.003931f
C2867 XM2/a_100_n297750# XM3/a_n158_n91050# 0.048706f
C2868 XM1/a_n100_73257# m1_1634_n2388# 7.34e-20
C2869 XM1/a_100_63302# XM2/a_100_n92142# 4.64e-21
C2870 XM2/a_n100_n303119# XM4/a_100_n96230# 2.56e-20
C2871 XM1/a_n158_163822# XM2/a_n158_10662# 4.64e-21
C2872 XM2/a_100_n187038# XM3/a_n100_19705# 0.005074f
C2873 XM3/a_n100_n67319# XM4/a_n100_n67319# 0.009521f
C2874 XM4/a_n100_72541# m1_1634_n2388# 0.072015f
C2875 XM4/w_n358_n132787# XM3/a_n100_n76643# 0.009128f
C2876 XM4/a_100_n62042# m1_1634_n2388# 6.1e-20
C2877 XM2/a_n158_n250302# XM3/a_n100_n44527# 1.45e-19
C2878 XM1/a_n100_n89011# XM3/a_n158_n37178# 2.85e-20
C2879 XM1/a_n158_n25730# XM2/a_n100_n181863# 4.56e-20
C2880 XM1/a_100_79098# XM2/a_100_n73690# 4.64e-21
C2881 XM3/a_n158_n106590# m1_1634_n2388# 6.1e-20
C2882 XM4/w_n358_n132787# XM3/a_n100_70469# 0.008782f
C2883 XM2/a_100_n142226# m1_1634_n2388# 0.017213f
C2884 XM1/a_n100_63205# XM3/a_n158_114078# 2.85e-20
C2885 XM4/w_n358_n132787# XM2/a_n158_n210762# 0.101988f
C2886 XM1/a_100_n7062# XM4/w_n358_n132787# 0.048442f
C2887 XM1/a_n100_77565# XM4/w_n358_n132787# 0.01363f
C2888 XM2/a_n100_n245127# XM3/a_n158_n38214# 0.005074f
C2889 XM1/a_n100_n124911# XM3/a_n100_n72499# 1.56e-19
C2890 XM4/w_n358_n132787# XM3/a_n100_15561# 0.009186f
C2891 XM4/w_n358_n132787# XM3/a_n158_n12314# 0.032295f
C2892 XM2/a_n158_n129046# XM3/a_n100_75649# 7.26e-20
C2893 XM1/a_n100_n173735# XM2/a_100_n326746# 7.26e-20
C2894 XM1/a_100_n159278# XM2/a_n158_n313566# 0.116862f
C2895 XM4/w_n358_n132787# XM3/a_n158_109934# 0.034136f
C2896 XM3/a_n100_n87003# XM4/a_n100_n87003# 0.009521f
C2897 XM2/a_n158_n324110# XM3/a_n100_n120155# 7.26e-20
C2898 XM2/a_n158_n171222# XM3/a_n100_33173# 7.26e-20
C2899 XM4/a_n100_33173# m1_1634_n2388# 0.072015f
C2900 XM1/a_100_n170766# XM3/a_n100_n119119# 2.85e-20
C2901 XM4/w_n358_n132787# XM3/a_n100_n116011# 0.009186f
C2902 XM4/a_100_n101410# m1_1634_n2388# 6.1e-20
C2903 XM2/a_100_n123774# XM3/a_n158_80926# 0.068179f
C2904 XM2/a_100_n100050# XM3/a_n158_105790# 0.077916f
C2905 XM2/a_n100_n100147# XM3/a_n100_104657# 0.006262f
C2906 XM2/a_100_n279298# XM3/a_n158_n73438# 0.077916f
C2907 XM1/a_n100_n91883# XM3/a_n100_n39347# 7.54e-19
C2908 XM1/a_n100_n54547# XM3/a_n158_n4026# 4.57e-19
C2909 XM2/a_100_n321474# XM3/a_n100_n114975# 0.005074f
C2910 XM2/a_100_n165950# XM3/a_n158_38450# 0.038969f
C2911 XM1/a_100_107818# XM2/a_100_n44694# 4.64e-21
C2912 XM4/w_n358_n132787# XM4/a_n100_127449# -0.004445f
C2913 XM1/a_n100_n45931# XM3/a_n158_6334# 2.85e-20
C2914 XM1/a_n100_n1415# XM3/a_n100_49749# 7.07e-19
C2915 XM1/a_100_102074# XM4/w_n358_n132787# 0.048442f
C2916 XM2/a_n100_n81695# m1_1634_n2388# 9.37e-19
C2917 XM1/a_100_71918# XM3/a_n100_122269# 1.61e-19
C2918 XM1/a_n158_28838# XM2/a_n100_n126507# 7.26e-20
C2919 XM2/a_n158_n231850# XM3/a_n100_n26915# 1.45e-19
C2920 XM1/a_n100_n28699# XM2/a_n158_n181766# 0.005074f
C2921 XM3/a_n100_53893# m1_1634_n2388# 0.072015f
C2922 XM1/a_n100_n53111# XM4/w_n358_n132787# 0.01363f
C2923 XM4/w_n358_n132787# XM2/a_100_n147498# 0.103341f
C2924 XM4/w_n358_n132787# XM3/a_n158_n51682# 0.03591f
C2925 XM4/a_n100_n38311# m1_1634_n2388# 0.072015f
C2926 XM2/a_100_n266118# m1_1634_n2388# 0.025819f
C2927 XM2/a_n100_n171319# XM4/a_100_35342# 2.56e-20
C2928 XM1/a_100_66174# XM3/a_n158_117186# 0.00544f
C2929 XM1/a_n100_24433# XM2/a_n100_n129143# 0.004501f
C2930 XM1/a_n100_8637# m1_1634_n2388# 9.16e-21
C2931 XM2/a_n158_n115866# XM3/a_n100_90153# 1.45e-19
C2932 XM4/w_n358_n132787# XM2/a_n158_n334654# 0.107093f
C2933 XM3/a_n100_n106687# XM4/a_n100_n106687# 0.009521f
C2934 XM1/a_n100_57461# XM2/a_100_n94778# 2.87e-20
C2935 XM4/w_n358_n132787# XM3/a_n158_95430# 0.032295f
C2936 XM3/a_n100_32137# XM4/a_n100_32137# 0.009521f
C2937 XM1/a_100_171002# XM2/a_100_15934# 4.64e-21
C2938 XM1/a_n100_22997# XM2/a_n100_n131779# 0.004501f
C2939 XM2/a_n158_n158042# XM3/a_n100_47677# 1.45e-19
C2940 XM4/w_n358_n132787# XM3/a_n158_40522# 0.03391f
C2941 XM1/a_n158_n120506# XM3/a_n100_n69391# 1.94e-20
C2942 XM2/a_100_n110594# XM3/a_n158_95430# 0.077916f
C2943 XM2/a_n100_n81695# XM3/a_n158_122366# 0.004352f
C2944 XM2/a_n158_n81598# XM3/a_n100_122269# 4.56e-20
C2945 XM1/a_n158_n146354# XM3/a_n100_n94255# 1.94e-20
C2946 XM4/w_n358_n132787# XM4/a_n100_88081# -0.004445f
C2947 XM1/a_n158_n97530# XM2/a_n100_n253035# 7.26e-20
C2948 XM2/a_100_n152770# XM3/a_n158_52954# 0.077916f
C2949 XM1/a_n158_n157842# XM2/a_n100_n313663# 7.26e-20
C2950 XM3/a_n100_n18627# m1_1634_n2388# 0.072015f
C2951 XM1/a_n100_n47367# XM3/a_n100_5201# 3.38e-19
C2952 XM1/a_n100_n126347# XM2/a_100_n281934# 7.26e-20
C2953 XM1/a_n158_70482# XM2/a_n158_n84234# 9.28e-21
C2954 XM1/a_100_17350# XM4/w_n358_n132787# 0.048442f
C2955 XM1/a_n100_56025# XM2/a_100_n97414# 7.26e-20
C2956 XM4/w_n358_n132787# XM3/a_n158_n91050# 0.038462f
C2957 XM4/a_n100_n77679# m1_1634_n2388# 0.072015f
C2958 XM2/a_100_n260846# XM3/a_n158_n55826# 0.077916f
C2959 XM1/a_n100_n90447# XM2/a_n158_n245030# 0.010147f
C2960 XM2/a_100_n194946# XM3/a_n158_10478# 0.077916f
C2961 XM1/a_n100_n152195# m1_1634_n2388# 9.15e-20
C2962 XM1/a_100_n21422# XM2/a_100_n173858# 4.64e-21
C2963 XM4/w_n358_n132787# XM2/a_n100_n86967# 0.025738f
C2964 XM1/a_100_57558# XM2/a_n100_n94875# 0.002238f
C2965 XM1/a_n100_37357# m1_1634_n2388# 1.3e-19
C2966 XM2/a_100_n303022# XM3/a_n100_n97363# 0.010147f
C2967 XM1/a_100_n97530# XM2/a_n158_n252938# 0.057664f
C2968 XM1/a_n100_n96191# XM3/a_n158_n44430# 1.96e-20
C2969 XM1/a_n100_n27263# XM3/a_n158_24982# 2.85e-20
C2970 XM1/a_n158_92022# XM2/a_n158_n63146# 4.64e-21
C2971 XM3/a_n100_n126371# XM4/a_n100_n126371# 0.009521f
C2972 XM1/a_100_n134866# XM2/a_100_n289842# 4.64e-21
C2973 XM1/a_n158_n55886# XM3/a_n100_n5159# 1.94e-20
C2974 XM2/a_n100_n205587# m1_1634_n2388# 7.61e-19
C2975 XM2/a_n100_n300483# XM3/a_n158_n96230# 0.005074f
C2976 XM1/a_n100_n55983# XM2/a_100_n210762# 7.26e-20
C2977 XM4/w_n358_n132787# XM2/a_100_n271390# 0.105846f
C2978 XM2/a_n158_n213398# XM3/a_n100_n9303# 7.26e-20
C2979 XM1/a_n100_n20083# XM2/a_100_n173858# 1.45e-19
C2980 XM3/a_n158_78854# m1_1634_n2388# 6.1e-20
C2981 XM1/a_100_86278# XM4/w_n358_n132787# 0.048442f
C2982 XM3/a_n100_111909# m1_1634_n2388# 0.072015f
C2983 XM1/a_n100_n47367# XM2/a_100_n202854# 7.26e-20
C2984 XM1/a_100_149462# XM4/w_n358_n132787# 0.048442f
C2985 XM4/a_100_122366# m1_1634_n2388# 6.1e-20
C2986 XM2/a_n158_n144862# XM3/a_n100_62181# 7.26e-20
C2987 XM2/a_n158_n297750# XM3/a_n158_n91050# 4.64e-21
C2988 XM3/a_n158_23946# m1_1634_n2388# 6.1e-20
C2989 XM1/a_100_63302# XM2/a_n158_n92142# 0.054158f
C2990 XM2/a_100_n210762# XM3/a_n100_n4123# 0.005074f
C2991 XM1/a_100_n9934# m1_1634_n2388# 0.001577f
C2992 XM4/w_n358_n132787# XM4/a_n100_48713# -0.004445f
C2993 XM2/a_n158_n187038# XM3/a_n100_19705# 7.26e-20
C2994 XM3/a_n100_n57995# m1_1634_n2388# 0.072015f
C2995 XM1/a_n100_150801# XM2/a_n158_n2518# 0.005074f
C2996 XM2/a_100_n139590# XM3/a_n158_67458# 0.014823f
C2997 XM1/a_n158_n143482# XM3/a_n100_n93219# 1.14e-20
C2998 XM1/a_n100_n137835# XM3/a_n158_n85870# 0.001028f
C2999 XM4/w_n358_n132787# XM3/a_n158_n130418# 0.038462f
C3000 XM4/a_n100_n117047# m1_1634_n2388# 0.072015f
C3001 XM1/a_n100_175213# XM2/a_n158_21206# 0.010147f
C3002 XM2/a_100_n181766# XM3/a_n158_24982# 0.044032f
C3003 XM1/a_n100_n1415# XM2/a_100_n155406# 1.45e-19
C3004 XM1/a_n100_n45931# XM2/a_100_n200218# 1.45e-19
C3005 iout_n XM4/w_n358_n132787# 0.003297f
C3006 XM1/a_n100_n136399# XM3/a_n158_n85870# 0.00173f
C3007 XM4/w_n358_n132787# XM4/a_n100_n22771# -0.004445f
C3008 XM4/w_n358_n132787# XM2/a_n100_n210859# 0.025625f
C3009 XM1/a_n100_n2851# XM4/w_n358_n132787# 0.013481f
C3010 XM2/a_n100_n247763# XM4/a_100_n43394# 2.56e-20
C3011 XM2/a_100_n242394# XM3/a_n158_n38214# 0.017549f
C3012 XM4/a_100_82998# m1_1634_n2388# 6.1e-20
C3013 XM2/a_n100_n329479# m1_1634_n2388# 0.001432f
C3014 XM2/a_100_n284570# XM3/a_n100_n79751# 0.010147f
C3015 XM2/a_n100_n129143# XM3/a_n100_75649# 0.005829f
C3016 XM1/a_n100_n173735# XM2/a_n158_n326746# 0.005074f
C3017 XM4/w_n358_n132787# XM4/a_n100_9345# -0.004445f
C3018 XM1/a_100_70482# XM3/a_n100_121233# 2.85e-20
C3019 XM4/w_n358_n132787# XM3/a_n100_109837# 0.009108f
C3020 XM1/a_n100_37357# XM2/a_100_n115866# 7.26e-20
C3021 XM1/a_n158_21658# XM3/a_n100_72541# 1.94e-20
C3022 XM1/a_n100_20125# m1_1634_n2388# 8.14e-20
C3023 XM1/a_n100_n111987# XM3/a_n158_n61006# 2.85e-20
C3024 XM1/a_n158_n183690# sw_bn 0.010925f
C3025 XM3/a_n100_n97363# m1_1634_n2388# 0.072015f
C3026 XM1/a_n100_n93319# XM2/a_100_n247666# 1.45e-19
C3027 XM1/a_n158_n37218# XM3/a_n100_13489# 1.94e-20
C3028 XM1/a_n158_n35782# XM3/a_n100_16597# 4.21e-21
C3029 XM1/a_n100_n103371# XM2/a_n158_n255574# 1.17e-21
C3030 XM2/a_n158_n123774# XM3/a_n158_80926# 4.64e-21
C3031 XM1/a_100_74790# XM4/w_n358_n132787# 0.048442f
C3032 XM2/a_100_n100050# XM3/a_n100_105693# 0.010147f
C3033 XM1/a_n158_14478# XM3/a_n100_66325# 1.94e-20
C3034 XM1/a_n158_10170# XM3/a_n158_62278# 1.14e-21
C3035 XM1/a_n158_n17114# XM2/a_n158_n171222# 9.28e-21
C3036 XM1/a_n100_179521# XM4/w_n358_n132787# 0.012279f
C3037 XM1/a_100_n131994# XM3/a_n158_n80690# 0.002646f
C3038 XM3/a_n100_129521# XM4/a_n100_129521# 0.009521f
C3039 XM2/a_n158_n321474# XM3/a_n100_n114975# 7.26e-20
C3040 XM1/a_100_n113326# XM2/a_100_n268754# 4.64e-21
C3041 XM2/a_n158_n165950# XM3/a_n158_38450# 4.64e-21
C3042 XM1/a_n100_70385# XM3/a_n158_121330# 2.85e-20
C3043 XM1/a_n158_n5626# XM3/a_n100_46641# 1e-20
C3044 XM2/a_100_n78962# m1_1634_n2388# 0.017213f
C3045 XM4/w_n358_n132787# XM3/a_n100_89117# 0.008944f
C3046 XM3/a_n100_84973# XM4/a_n100_84973# 0.009521f
C3047 XM4/w_n358_n132787# XM4/a_n100_n62139# -0.004445f
C3048 XM3/a_n158_n33034# m1_1634_n2388# 6.1e-20
C3049 XM1/a_n100_n130655# XM2/a_100_n284570# 1.45e-19
C3050 XM1/a_n158_102074# XM2/a_n158_n52602# 9.28e-21
C3051 XM1/a_n100_30177# XM4/w_n358_n132787# 0.013602f
C3052 XM4/a_100_43630# m1_1634_n2388# 6.1e-20
C3053 XM4/w_n358_n132787# XM2/a_n158_n147498# 0.102053f
C3054 XM1/a_n100_96233# XM2/a_n158_n57874# 0.010147f
C3055 XM4/w_n358_n132787# XM3/a_n100_34209# 0.009186f
C3056 XM4/w_n358_n132787# XM1/a_100_139410# 0.053546f
C3057 XM1/a_100_66174# XM3/a_n100_117089# 2.85e-20
C3058 XM1/a_n100_n110551# XM3/a_n158_n59970# 2.85e-20
C3059 XM1/a_100_100638# XM2/a_n100_n52699# 0.005074f
C3060 XM4/w_n358_n132787# XM2/a_n100_n334751# 0.025163f
C3061 XM4/w_n358_n132787# XM1/a_100_n147790# 0.054609f
C3062 XM1/a_n100_57461# XM2/a_n158_n94778# 0.002238f
C3063 XM1/a_n100_n109115# m1_1634_n2388# 1.18e-19
C3064 XM1/a_n100_170905# XM2/a_n158_18570# 0.005074f
C3065 XM1/a_100_n180818# XM2/a_n158_n334654# 0.116862f
C3066 XM2/a_100_n266118# XM3/a_n100_n62139# 0.005074f
C3067 XM3/a_n100_5201# m1_1634_n2388# 0.072015f
C3068 XM4/a_n100_106729# m1_1634_n2388# 0.072015f
C3069 XM4/w_n358_n132787# XM1/a_n100_n132091# 0.013471f
C3070 XM1/a_n100_n124911# XM4/w_n358_n132787# 0.013401f
C3071 XM2/a_100_n81598# XM3/a_n158_123402# 0.077916f
C3072 XM2/a_n100_n81695# XM3/a_n100_122269# 0.001118f
C3073 XM4/w_n358_n132787# XM3/a_n100_n42455# 0.009186f
C3074 XM4/a_100_n27854# m1_1634_n2388# 6.1e-20
C3075 XM2/a_n158_n36786# XM4/w_n358_n132787# 0.105622f
C3076 XM1/a_n158_60430# XM2/a_n158_n94778# 4.64e-21
C3077 XM1/a_n100_n100499# m1_1634_n2388# 1.3e-19
C3078 XM1/a_n100_n66035# XM3/a_n100_n14483# 6.24e-19
C3079 XM4/w_n358_n132787# XM4/a_n100_n101507# -0.004445f
C3080 XM3/a_n158_n72402# m1_1634_n2388# 6.1e-20
C3081 XM1/a_n100_n126347# XM2/a_n158_n281934# 0.005074f
C3082 XM1/a_n100_n172299# m1_1634_n2388# 1.26e-19
C3083 XM1/a_n100_56025# XM2/a_n158_n97414# 0.005074f
C3084 XM2/a_n100_n115963# XM4/a_100_88178# 2.56e-20
C3085 XM1/a_n100_66077# XM2/a_100_n89506# 7.26e-20
C3086 XM3/a_n100_72541# m1_1634_n2388# 0.072015f
C3087 XM1/a_100_n21422# XM2/a_n158_n173858# 0.003528f
C3088 XM4/w_n358_n132787# XM2/a_100_n84234# 0.103342f
C3089 XM2/a_n158_n303022# XM3/a_n100_n97363# 1.45e-19
C3090 XM1/a_100_n113326# XM3/a_n158_n62042# 0.00544f
C3091 XM1/a_100_n106146# XM4/w_n358_n132787# 0.048442f
C3092 XM1/a_100_n97530# XM2/a_n100_n253035# 0.005074f
C3093 XM1/a_100_n134866# XM2/a_n158_n289842# 0.099726f
C3094 XM1/a_n100_n73215# XM3/a_n100_n20699# 0.001015f
C3095 XM1/a_n100_n55983# XM2/a_n158_n210762# 0.005074f
C3096 XM2/a_100_n202854# m1_1634_n2388# 0.025819f
C3097 XM3/a_n100_17633# m1_1634_n2388# 0.072015f
C3098 XM1/a_n100_79001# m1_1634_n2388# 9.31e-20
C3099 XM4/w_n358_n132787# XM2/a_n158_n271390# 0.105802f
C3100 XM3/a_n100_112945# XM4/a_n100_112945# 0.009521f
C3101 XM1/a_n100_n20083# XM2/a_n158_n173858# 0.010147f
C3102 XM1/a_100_n146354# XM3/a_n100_n94255# 2.85e-20
C3103 XM1/a_n100_114901# XM4/w_n358_n132787# 0.012279f
C3104 XM1/a_n100_n47367# XM2/a_n158_n202854# 0.005074f
C3105 XM1/a_100_120742# XM2/a_n100_n34247# 0.004978f
C3106 XM4/a_n100_67361# m1_1634_n2388# 0.072014f
C3107 XM4/w_n358_n132787# XM3/a_n158_59170# 0.039522f
C3108 XM2/a_n100_n297847# XM3/a_n158_n91050# 0.005074f
C3109 XM4/w_n358_n132787# XM3/a_n100_n81823# 0.009026f
C3110 XM4/a_100_n67222# m1_1634_n2388# 6.1e-20
C3111 XM1/a_100_63302# XM2/a_n100_n92239# 0.005074f
C3112 XM2/a_n158_n210762# XM3/a_n100_n4123# 7.26e-20
C3113 XM1/a_n158_n119070# XM2/a_n158_n274026# 4.64e-21
C3114 XM1/a_n158_n109018# XM2/a_n158_n263482# 9.28e-21
C3115 XM2/a_n158_10662# XM4/w_n358_n132787# 0.106353f
C3116 XM3/a_n158_n111770# m1_1634_n2388# 6.1e-20
C3117 XM1/a_100_n21422# XM4/w_n358_n132787# 0.054609f
C3118 XM1/a_100_n93222# XM2/a_n158_n247666# 0.116862f
C3119 XM2/a_n158_n139590# XM3/a_n158_67458# 4.64e-21
C3120 XM1/a_100_46070# XM2/a_n158_n107958# 0.116862f
C3121 XM1/a_n158_n25730# XM2/a_n158_n179130# 4.64e-21
C3122 XM1/a_n100_n163683# XM2/a_100_n318838# 7.26e-20
C3123 XM2/a_n158_n181766# XM3/a_n158_24982# 4.64e-21
C3124 XM1/a_n158_n25730# XM3/a_n100_24885# 1.94e-20
C3125 XM1/a_n100_n20083# XM4/w_n358_n132787# 0.013373f
C3126 XM1/a_100_n119070# XM3/a_n158_n67222# 0.003891f
C3127 XM1/a_n100_n1415# XM2/a_n158_n155406# 0.010147f
C3128 XM1/a_100_146590# XM4/w_n358_n132787# 0.048442f
C3129 XM2/a_100_n332018# XM3/a_n158_n126274# 0.077916f
C3130 XM4/w_n358_n132787# XM3/a_n158_n17494# 0.033613f
C3131 XM4/a_n100_n4123# m1_1634_n2388# 0.072015f
C3132 XM1/a_n100_n45931# XM2/a_n158_n200218# 0.010147f
C3133 XM1/a_n158_24530# XM3/a_n100_75649# 1.94e-20
C3134 XM2/a_n100_n142323# m1_1634_n2388# 7.61e-19
C3135 XM4/w_n358_n132787# XM2/a_100_n208126# 0.106508f
C3136 XM1/a_n158_n4190# XM2/a_n158_n158042# 9.28e-21
C3137 XM2/a_n100_n21067# XM1/a_n158_135102# 2.27e-20
C3138 XM2/a_n158_n242394# XM3/a_n158_n38214# 4.64e-21
C3139 XM1/a_n100_n14339# XM3/a_n158_37414# 1.73e-20
C3140 XM3/a_n158_97502# m1_1634_n2388# 6.1e-20
C3141 XM2/a_100_n326746# m1_1634_n2388# 0.017213f
C3142 XM1/a_n100_n41623# XM3/a_n158_10478# 2.85e-20
C3143 XM4/a_n100_27993# m1_1634_n2388# 0.072015f
C3144 XM4/w_n358_n132787# XM3/a_n100_n121191# 0.009026f
C3145 XM4/a_100_n106590# m1_1634_n2388# 6.1e-20
C3146 XM2/a_n158_n284570# XM3/a_n100_n79751# 1.45e-19
C3147 XM1/a_100_n90350# XM2/a_n158_n245030# 0.116862f
C3148 XM1/a_100_n153534# XM2/a_n158_n308294# 0.116862f
C3149 XM1/a_n100_173777# XM2/a_100_18570# 7.26e-20
C3150 XM1/a_n100_37357# XM2/a_n158_n115866# 0.005074f
C3151 XM1/a_100_n91786# XM3/a_n100_n40383# 0.00177f
C3152 XM3/a_n158_42594# m1_1634_n2388# 6.1e-20
C3153 XM1/a_n100_n93319# XM2/a_n158_n247666# 0.010147f
C3154 XM2/a_n100_n245127# XM4/a_100_n38214# 2.56e-20
C3155 XM2/a_100_n239758# XM3/a_n158_n33034# 0.046369f
C3156 XM3/a_n100_52857# XM4/a_n100_52857# 0.009521f
C3157 XM1/a_100_14478# XM3/a_n100_65289# 2.85e-20
C3158 XM4/w_n358_n132787# XM4/a_n100_122269# -0.004445f
C3159 XM1/a_n100_n103371# XM2/a_n100_n255671# 0.005189f
C3160 XM1/a_n158_n53014# XM2/a_n158_n208126# 4.64e-21
C3161 XM2/a_n100_n123871# XM3/a_n158_80926# 0.005074f
C3162 XM1/a_n100_n160811# XM3/a_n158_n109698# 2.85e-20
C3163 XM2/a_n158_n100050# XM3/a_n100_105693# 1.45e-19
C3164 XM1/a_n100_n22955# XM3/a_n158_29126# 2.85e-20
C3165 XM1/a_100_n113326# XM2/a_n158_n268754# 0.055716f
C3166 XM4/w_n358_n132787# XM3/a_n158_n56862# 0.03799f
C3167 XM4/a_n100_n43491# m1_1634_n2388# 0.072015f
C3168 XM2/a_n100_n166047# XM3/a_n158_38450# 0.005074f
C3169 XM1/a_100_n5626# XM3/a_n100_45605# 8.37e-19
C3170 XM1/a_100_n58758# XM3/a_n100_n8267# 2.85e-20
C3171 XM2/a_100_n18334# XM1/a_100_135102# 4.64e-21
C3172 XM1/a_n100_n130655# XM2/a_n158_n284570# 0.010147f
C3173 XM1/a_n158_28838# XM2/a_n158_n123774# 4.64e-21
C3174 XM1/a_n100_n31571# m1_1634_n2388# 1e-19
C3175 XM1/a_n158_n11370# XM3/a_n100_40425# 1.94e-20
C3176 XM4/w_n358_n132787# XM2/a_n100_n147595# 0.02472f
C3177 XM1/a_n158_n90350# XM2/a_n158_n245030# 9.28e-21
C3178 XM2/a_n100_n266215# m1_1634_n2388# 7.61e-19
C3179 XM2/a_100_n313566# XM3/a_n158_n108662# 0.077916f
C3180 XM1/a_100_n107582# XM4/w_n358_n132787# 0.054646f
C3181 XM1/a_100_n96094# XM2/a_n158_n250302# 0.116862f
C3182 XM3/a_n100_n1015# m1_1634_n2388# 0.072015f
C3183 XM4/w_n358_n132787# XM2/a_100_n332018# 0.103342f
C3184 XM1/a_n100_57461# XM2/a_n100_n94875# 0.002708f
C3185 XM2/a_100_n205490# XM3/a_n100_1057# 0.005074f
C3186 XM2/a_n100_n52699# XM4/w_n358_n132787# 0.012081f
C3187 XM1/a_n100_n51675# XM2/a_100_n205490# 1.45e-19
C3188 XM4/w_n358_n132787# XM4/a_n100_82901# -0.004445f
C3189 XM3/a_n100_n23807# m1_1634_n2388# 0.072015f
C3190 XM2/a_n158_n266118# XM3/a_n100_n62139# 7.26e-20
C3191 XM2/a_n100_n163411# XM4/a_n100_40425# 6.78e-21
C3192 XM2/a_100_n81598# XM3/a_n100_123305# 0.010147f
C3193 XM4/w_n358_n132787# XM3/a_n158_n96230# 0.038462f
C3194 XM4/a_n100_n82859# m1_1634_n2388# 0.072015f
C3195 XM1/a_n158_n97530# XM2/a_n158_n250302# 4.64e-21
C3196 XM2/a_100_n221306# XM3/a_n158_n15422# 0.077916f
C3197 XM1/a_n158_60430# XM2/a_n100_n94875# 7.26e-20
C3198 XM1/a_n100_n119167# XM2/a_100_n274026# 7.26e-20
C3199 XM1/a_100_n93222# XM3/a_n100_n41419# 2.85e-20
C3200 XM1/a_n158_n157842# XM2/a_n158_n310930# 4.64e-21
C3201 XM1/a_n100_n101935# XM3/a_n158_n50646# 3.15e-21
C3202 XM1/a_100_n143482# XM4/w_n358_n132787# 0.048442f
C3203 XM2/a_100_n263482# XM3/a_n100_n56959# 0.005074f
C3204 XM1/a_n158_n169330# XM3/a_n100_n117047# 1.94e-20
C3205 XM1/a_n100_56025# XM2/a_n100_n97511# 0.001385f
C3206 XM1/a_n100_66077# XM2/a_n158_n89506# 0.005074f
C3207 XM1/a_100_n21422# XM2/a_n100_n173955# 0.005074f
C3208 XM4/w_n358_n132787# XM2/a_n158_n84234# 0.103313f
C3209 XM1/a_100_n172202# XM3/a_n100_n121191# 2.85e-20
C3210 XM1/a_100_n134866# XM2/a_n100_n289939# 0.005074f
C3211 XM1/a_100_n97530# XM2/a_100_n250302# 4.64e-21
C3212 XM1/a_n100_n81831# XM2/a_100_n237122# 7.26e-20
C3213 XM4/w_n358_n132787# XM3/a_n100_52857# 0.009186f
C3214 XM4/a_100_117186# m1_1634_n2388# 6.1e-20
C3215 XM1/a_100_n110454# XM3/a_n100_n60067# 2.85e-20
C3216 XM1/a_n100_n55983# XM2/a_n100_n210859# 5.53e-19
C3217 XM4/w_n358_n132787# XM2/a_n100_n271487# 0.024015f
C3218 XM4/w_n358_n132787# XM4/a_n100_43533# -0.004445f
C3219 XM2/a_n100_n113327# XM4/a_100_93358# 2.56e-20
C3220 XM3/a_n100_n63175# m1_1634_n2388# 0.072015f
C3221 XM4/w_n358_n132787# XM1/a_100_136538# 0.049664f
C3222 XM3/a_n158_113042# m1_1634_n2388# 6.1e-20
C3223 XM1/a_100_n143482# XM2/a_n158_n297750# 0.116862f
C3224 XM1/a_n158_148026# XM2/a_n158_n7790# 4.64e-21
C3225 XM1/a_n100_44537# XM4/w_n358_n132787# 0.01363f
C3226 XM2/a_100_n142226# XM3/a_n100_62181# 0.005074f
C3227 XM4/a_n100_n122227# m1_1634_n2388# 0.072015f
C3228 XM2/a_n100_n300483# XM4/a_100_n96230# 2.56e-20
C3229 XM2/a_100_n295114# XM3/a_n158_n91050# 0.006254f
C3230 XM1/a_100_63302# XM2/a_100_n89506# 4.64e-21
C3231 XM3/a_n100_n13447# XM4/a_n100_n13447# 0.009521f
C3232 XM2/a_100_n337290# XM3/a_n100_n132587# 0.005078f
C3233 XM1/a_n158_n119070# XM2/a_n100_n274123# 7.26e-20
C3234 XM1/a_n158_n114762# XM3/a_n100_n64211# 1.94e-20
C3235 XM2/a_100_n184402# XM3/a_n100_19705# 0.005074f
C3236 XM1/a_n100_114901# XM2/a_100_n39422# 1.45e-19
C3237 XM1/a_100_n182254# sw_b 2.29e-21
C3238 XM1/a_n100_n11467# XM2/a_100_n165950# 1.45e-19
C3239 XM1/a_n100_44537# XM2/a_100_n110594# 7.26e-20
C3240 XM2/a_n100_n139687# XM3/a_n158_67458# 0.005074f
C3241 XM4/w_n358_n132787# XM4/a_n100_n27951# -0.004445f
C3242 XM1/a_n158_n25730# XM2/a_n100_n179227# 7.26e-20
C3243 XM1/a_100_1554# XM4/w_n358_n132787# 0.048442f
C3244 XM1/a_n100_n163683# XM2/a_n158_n318838# 0.005074f
C3245 XM2/a_n100_n181863# XM3/a_n158_24982# 0.005074f
C3246 XM1/a_n100_n18647# m1_1634_n2388# 1.3e-19
C3247 XM1/a_n100_120645# XM2/a_n100_n34247# 7.77e-20
C3248 XM3/a_n100_91189# m1_1634_n2388# 0.072014f
C3249 XM4/a_100_77818# m1_1634_n2388# 6.1e-20
C3250 XM1/a_n100_n71779# XM4/w_n358_n132787# 0.013059f
C3251 XM2/a_n100_n187135# XM4/a_100_17730# 8.43e-21
C3252 XM2/a_100_n139590# m1_1634_n2388# 0.023368f
C3253 XM2/a_100_n245030# XM3/a_n100_n39347# 0.010147f
C3254 XM1/a_100_n73118# XM4/w_n358_n132787# 0.052778f
C3255 XM3/a_n100_20741# XM4/a_n100_20741# 0.009521f
C3256 XM3/a_n100_36281# m1_1634_n2388# 0.072015f
C3257 XM1/a_n100_63205# XM3/a_n158_115114# 2.85e-20
C3258 XM3/a_n100_n102543# m1_1634_n2388# 0.072015f
C3259 XM2/a_n100_n242491# XM3/a_n158_n38214# 0.005074f
C3260 XM4/w_n358_n132787# XM2/a_n158_n208126# 0.103244f
C3261 XM1/a_n100_n104807# XM2/a_n100_n260943# 0.004742f
C3262 XM1/a_n100_30177# XM3/a_n100_81865# 1.17e-19
C3263 XM1/a_n100_n30135# XM2/a_100_n184402# 1.45e-19
C3264 XM4/w_n358_n132787# XM3/a_n158_77818# 0.038602f
C3265 XM2/a_100_n129046# XM3/a_n100_76685# 0.010147f
C3266 XM3/a_n100_n33131# XM4/a_n100_n33131# 0.009521f
C3267 XM4/w_n358_n132787# XM3/a_n158_110970# 0.032295f
C3268 XM1/a_100_n48706# XM4/w_n358_n132787# 0.048442f
C3269 XM1/a_n158_13042# XM3/a_n100_64253# 2.69e-20
C3270 XM2/a_n158_n239758# XM3/a_n158_n33034# 4.64e-21
C3271 XM1/a_100_n81734# XM3/a_n100_n30023# 2.85e-20
C3272 XM1/a_n100_34485# XM2/a_100_n121138# 7.26e-20
C3273 XM4/w_n358_n132787# XM3/a_n100_n8267# 0.009186f
C3274 XM2/a_100_n171222# XM3/a_n100_34209# 0.010147f
C3275 XM4/w_n358_n132787# XM3/a_n158_22910# 0.035697f
C3276 XM1/a_100_n70246# XM3/a_n100_n19663# 2.85e-20
C3277 XM1/a_n158_n53014# XM2/a_n100_n208223# 7.26e-20
C3278 XM1/a_n100_n28699# m1_1634_n2388# 9.49e-20
C3279 XM1/a_n158_n137738# XM2/a_n158_n292478# 9.28e-21
C3280 XM4/w_n358_n132787# XM4/a_n100_n67319# -0.004445f
C3281 XM3/a_n158_n38214# m1_1634_n2388# 6.1e-20
C3282 XM2/a_100_n100050# XM3/a_n158_106826# 0.03157f
C3283 XM1/a_100_31710# XM2/a_100_n123774# 4.64e-21
C3284 XM4/a_100_38450# m1_1634_n2388# 6.1e-20
C3285 XM1/a_n100_100541# XM2/a_n158_n52602# 0.005074f
C3286 XM1/a_n158_n162150# XM3/a_n100_n110831# 3.89e-20
C3287 XM3/a_n100_n2051# XM4/a_n100_n2051# 0.009521f
C3288 XM1/a_n100_166597# XM2/a_n100_10565# 9.94e-19
C3289 XM2/a_100_n318838# XM3/a_n100_n114975# 0.004271f
C3290 XM1/a_100_n113326# XM2/a_n100_n268851# 0.005074f
C3291 XM1/a_n100_n37315# XM2/a_100_n192310# 7.26e-20
C3292 XM1/a_100_28838# XM2/a_100_n126410# 4.64e-21
C3293 XM1/a_100_n177946# XM2/a_n158_n332018# 0.116862f
C3294 XM1/a_100_n126250# XM3/a_n100_n74571# 9.37e-19
C3295 XM3/a_n100_21# XM4/a_n100_21# 0.009521f
C3296 XM1/a_100_166694# XM4/w_n358_n132787# 0.052807f
C3297 XM2/a_n100_n79059# m1_1634_n2388# 7.61e-19
C3298 XM1/a_100_n11370# XM3/a_n100_39389# 2.85e-20
C3299 XM1/a_100_71918# XM3/a_n100_123305# 5.71e-20
C3300 XM1/a_n158_28838# XM2/a_n100_n123871# 7.26e-20
C3301 XM4/w_n358_n132787# XM2/a_100_n144862# 0.10657f
C3302 XM2/a_100_n263482# m1_1634_n2388# 0.017213f
C3303 XM1/a_n158_n77426# XM2/a_n158_n231850# 9.28e-21
C3304 XM3/a_n100_n52815# XM4/a_n100_n52815# 0.009521f
C3305 XM2/a_n100_n168683# XM4/a_100_35342# 6.59e-21
C3306 XM1/a_n100_96233# XM4/w_n358_n132787# 0.012279f
C3307 XM4/a_n100_101549# m1_1634_n2388# 0.072015f
C3308 XM2/a_100_n115866# XM3/a_n100_91189# 0.005074f
C3309 XM4/w_n358_n132787# XM2/a_n158_n332018# 0.107093f
C3310 XM2/a_100_n226578# XM3/a_n100_n21735# 0.010147f
C3311 XM4/w_n358_n132787# XM3/a_n100_n47635# 0.009186f
C3312 XM4/a_100_n33034# m1_1634_n2388# 6.1e-20
C3313 XM2/a_n158_n205490# XM3/a_n100_1057# 7.26e-20
C3314 XM3/a_n158_61242# m1_1634_n2388# 6.1e-20
C3315 XM1/a_n100_n51675# XM2/a_n158_n205490# 0.010147f
C3316 XM2/a_100_n158042# XM3/a_n100_48713# 0.005074f
C3317 XM4/w_n358_n132787# XM4/a_n100_n106687# -0.004445f
C3318 XM3/a_n158_n77582# m1_1634_n2388# 6.1e-20
C3319 XM2/a_n158_23842# XM1/a_n100_176649# 0.005074f
C3320 XM1/a_n100_50281# XM4/w_n358_n132787# 0.013487f
C3321 XM2/a_n158_n81598# XM3/a_n100_123305# 1.45e-19
C3322 XM1/a_n158_n97530# XM2/a_n100_n250399# 7.26e-20
C3323 XM1/a_n158_n157842# XM2/a_n100_n311027# 7.26e-20
C3324 XM1/a_n100_n119167# XM2/a_n158_n274026# 0.005074f
C3325 XM1/a_n100_n33007# XM3/a_n158_18766# 2.32e-20
C3326 XM1/a_n100_n104807# XM3/a_n158_n53754# 4.72e-19
C3327 XM1/a_n158_n70246# XM3/a_n100_n18627# 1.94e-20
C3328 XM1/a_n100_n126347# XM2/a_100_n279298# 7.26e-20
C3329 XM2/a_n158_n263482# XM3/a_n100_n56959# 7.26e-20
C3330 XM1/a_100_n160714# XM3/a_n158_n109698# 0.002193f
C3331 XM2/a_n100_n160775# XM4/a_n100_45605# 2.84e-20
C3332 XM1/a_100_n173638# m1_1634_n2388# 9.1e-19
C3333 XM3/a_n100_n72499# XM4/a_n100_n72499# 0.009521f
C3334 XM1/a_n100_122081# XM4/w_n358_n132787# 0.012203f
C3335 XM4/w_n358_n132787# XM2/a_n100_n84331# 0.026236f
C3336 XM1/a_100_13042# XM4/w_n358_n132787# 0.054705f
C3337 XM1/a_100_n97530# XM2/a_n158_n250302# 0.036243f
C3338 XM1/a_n100_n81831# XM2/a_n158_n237122# 0.005074f
C3339 XM2/a_n100_n202951# m1_1634_n2388# 7.61e-19
C3340 XM4/a_n100_62181# m1_1634_n2388# 0.072015f
C3341 XM4/w_n358_n132787# XM3/a_n100_n87003# 0.009186f
C3342 XM4/a_100_n72402# m1_1634_n2388# 6.1e-20
C3343 XM1/a_n100_129261# XM2/a_100_n26242# 7.26e-20
C3344 XM4/w_n358_n132787# XM2/a_100_n268754# 0.103341f
C3345 XM1/a_n100_31613# m1_1634_n2388# 1.07e-19
C3346 XM1/a_n100_n129219# XM4/w_n358_n132787# 0.013573f
C3347 XM1/a_100_n103274# XM3/a_n100_n51779# 6.34e-20
C3348 XM1/a_n100_169469# XM2/a_n158_15934# 0.005724f
C3349 XM2/a_n100_n5251# XM4/w_n358_n132787# 0.011694f
C3350 XM1/a_100_123614# XM2/a_100_n31514# 4.64e-21
C3351 XM3/a_n158_n116950# m1_1634_n2388# 6.1e-20
C3352 XM1/a_n100_n47367# XM2/a_100_n200218# 7.26e-20
C3353 XM3/a_n100_112945# m1_1634_n2388# 0.072015f
C3354 XM1/a_100_43198# XM3/a_n100_95333# 2.85e-20
C3355 XM2/a_n158_n142226# XM3/a_n100_62181# 7.26e-20
C3356 XM2/a_n158_n295114# XM3/a_n158_n91050# 4.64e-21
C3357 XM1/a_100_63302# XM2/a_n158_n89506# 0.039748f
C3358 XM2/a_100_n208126# XM3/a_n100_n4123# 0.005074f
C3359 XM2/a_n158_n337290# XM3/a_n100_n132587# 7.26e-20
C3360 XM1/a_n158_n86042# XM2/a_n158_n239758# 9.28e-21
C3361 XM1/a_n100_n38751# XM4/w_n358_n132787# 0.013441f
C3362 XM2/a_n158_n184402# XM3/a_n100_19705# 7.26e-20
C3363 XM1/a_100_n177946# XM3/a_n100_n126371# 2.85e-20
C3364 XM1/a_n100_n11467# XM2/a_n158_n165950# 0.010147f
C3365 XM1/a_n100_44537# XM2/a_n158_n110594# 0.005074f
C3366 XM4/w_n358_n132787# XM3/a_n158_n22674# 0.036692f
C3367 XM4/a_n100_n9303# m1_1634_n2388# 0.072015f
C3368 XM1/a_n100_34485# XM3/a_n158_85070# 2.85e-20
C3369 XM3/a_n100_73577# XM4/a_n100_73577# 0.009521f
C3370 XM2/a_100_n136954# XM3/a_n158_67458# 0.040138f
C3371 XM2/a_n100_n297847# XM4/a_100_n91050# 2.56e-20
C3372 XM2/a_100_n292478# XM3/a_n158_n85870# 0.057664f
C3373 XM3/a_n100_n92183# XM4/a_n100_n92183# 0.009521f
C3374 XM1/a_n158_40326# XM2/a_n158_n113230# 4.64e-21
C3375 XM4/a_n100_22813# m1_1634_n2388# 0.072015f
C3376 XM2/a_100_n179130# XM3/a_n158_24982# 0.010928f
C3377 XM1/a_n158_n183690# XM2/a_n158_n337290# 4.64e-21
C3378 XM4/w_n358_n132787# XM3/a_n100_n126371# 0.009055f
C3379 XM4/a_100_n111770# m1_1634_n2388# 6.1e-20
C3380 XM1/a_n158_n154970# XM3/a_n100_n104615# 2.4e-21
C3381 XM4/w_n358_n132787# XM3/a_n100_71505# 0.009186f
C3382 XM2/a_n158_n245030# XM3/a_n100_n39347# 1.45e-19
C3383 XM3/a_n158_6334# m1_1634_n2388# 6.1e-20
C3384 XM1/a_n158_38890# XM2/a_n158_n115866# 9.28e-21
C3385 XM4/w_n358_n132787# XM2/a_n100_n208223# 0.026252f
C3386 XM2/a_100_n200218# XM3/a_n100_6237# 0.005074f
C3387 XM2/a_n100_n326843# m1_1634_n2388# 7.61e-19
C3388 XM1/a_100_n137738# XM2/a_n158_n292478# 0.116862f
C3389 XM1/a_n100_n104807# XM2/a_100_n258210# 7.26e-20
C3390 XM1/a_n100_70385# m1_1634_n2388# 1.21e-19
C3391 XM4/w_n358_n132787# XM3/a_n100_16597# 0.0085f
C3392 XM1/a_n100_n30135# XM2/a_n158_n184402# 0.010147f
C3393 XM4/w_n358_n132787# XM4/a_n100_117089# -0.004445f
C3394 XM1/a_n158_37454# XM2/a_n158_n118502# 4.64e-21
C3395 XM4/a_n100_2093# m1_1634_n2388# 0.072015f
C3396 XM1/a_n100_n8595# XM3/a_n158_42594# 2.85e-20
C3397 XM1/a_n158_114998# XM2/a_n158_n39422# 9.28e-21
C3398 XM1/a_100_104946# XM2/a_100_n49966# 4.64e-21
C3399 XM2/a_n158_n129046# XM3/a_n100_76685# 1.45e-19
C3400 XM1/a_n158_8734# XM3/a_n158_59170# 1.14e-21
C3401 XM1/a_n158_n117634# XM2/a_n158_n271390# 9.28e-21
C3402 XM1/a_100_n2754# XM4/w_n358_n132787# 0.054609f
C3403 XM1/a_100_70482# XM3/a_n100_122269# 2.85e-20
C3404 XM4/w_n358_n132787# XM3/a_n100_110873# 0.009186f
C3405 XM1/a_100_57558# XM3/a_n100_107765# 1.09e-21
C3406 XM2/a_n100_n239855# XM3/a_n158_n33034# 0.005074f
C3407 XM1/a_n100_34485# XM2/a_n158_n121138# 0.005074f
C3408 XM4/w_n358_n132787# XM3/a_n158_n62042# 0.038462f
C3409 XM4/a_n100_n48671# m1_1634_n2388# 0.072015f
C3410 XM2/a_n158_n171222# XM3/a_n100_34209# 1.45e-19
C3411 XM1/a_n100_15817# m1_1634_n2388# 1.14e-19
C3412 XM1/a_n100_n129219# XM3/a_n100_n77679# 2.68e-19
C3413 XM2/a_100_n123774# XM3/a_n158_81962# 0.077916f
C3414 XM3/a_n100_n111867# XM4/a_n100_n111867# 0.009521f
C3415 XM2/a_100_n100050# XM3/a_n100_106729# 0.005074f
C3416 XM2/a_n158_n100050# XM3/a_n158_106826# 4.64e-21
C3417 XM1/a_100_31710# XM2/a_n158_n123774# 0.050264f
C3418 XM1/a_n158_143718# XM2/a_n158_n10426# 9.28e-21
C3419 XM2/a_n158_n318838# XM3/a_n100_n114975# 4.26e-20
C3420 XM1/a_100_n113326# XM2/a_100_n266118# 4.64e-21
C3421 XM2/a_100_n165950# XM3/a_n158_39486# 0.077916f
C3422 XM1/a_n100_70385# XM3/a_n158_122366# 1.72e-19
C3423 XM1/a_n100_n169427# XM3/a_n158_n116950# 8.08e-19
C3424 XM1/a_n100_n37315# XM2/a_n158_n192310# 0.005074f
C3425 XM1/a_100_28838# XM2/a_n158_n126410# 0.073242f
C3426 XM1/a_100_n53014# XM4/w_n358_n132787# 0.054624f
C3427 XM1/a_n100_106285# XM2/a_100_n47330# 1.45e-19
C3428 XM2/a_100_n76326# m1_1634_n2388# 0.020923f
C3429 XM1/a_n158_n80298# XM3/a_n100_n30023# 1.38e-20
C3430 XM2/a_100_n274026# XM3/a_n158_n68258# 0.077916f
C3431 XM3/a_n100_54929# m1_1634_n2388# 0.072015f
C3432 XM4/w_n358_n132787# XM4/a_n100_77721# -0.004445f
C3433 XM1/a_n158_24530# XM2/a_n158_n129046# 4.64e-21
C3434 XM4/w_n358_n132787# XM2/a_n158_n144862# 0.101988f
C3435 XM2/a_100_n316202# XM3/a_n100_n109795# 0.005074f
C3436 XM1/a_100_66174# XM3/a_n100_118125# 2.85e-20
C3437 XM3/a_n100_n28987# m1_1634_n2388# 0.072015f
C3438 XM1/a_100_25966# XM4/w_n358_n132787# 0.053885f
C3439 XM1/a_n100_142185# XM2/a_n158_n13062# 0.005074f
C3440 XM4/w_n358_n132787# XM3/a_n158_96466# 0.038462f
C3441 XM2/a_n158_n115866# XM3/a_n100_91189# 7.26e-20
C3442 XM4/w_n358_n132787# XM2/a_n100_n332115# 0.025632f
C3443 XM2/a_n158_n226578# XM3/a_n100_n21735# 1.45e-19
C3444 XM4/w_n358_n132787# XM3/a_n158_n101410# 0.038834f
C3445 XM4/a_n100_n88039# m1_1634_n2388# 0.072014f
C3446 XM1/a_n158_n48706# XM3/a_n100_2093# 1.94e-20
C3447 XM1/a_100_171002# XM2/a_100_18570# 4.64e-21
C3448 XM4/w_n358_n132787# XM3/a_n158_41558# 0.032295f
C3449 XM2/a_n158_n158042# XM3/a_n100_48713# 7.26e-20
C3450 XM1/a_n158_133666# XM2/a_n158_n20970# 9.28e-21
C3451 XM1/a_100_n64502# XM3/a_n100_n13447# 2.85e-20
C3452 XM2/a_n100_n166047# XM4/a_100_40522# 1.9e-20
C3453 XM2/a_100_n110594# XM3/a_n158_96466# 0.013654f
C3454 XM2/a_100_n81598# XM3/a_n158_124438# 0.077916f
C3455 XM1/a_n100_89053# XM2/a_n100_n63243# 0.005248f
C3456 XM1/a_n158_66174# XM2/a_n158_n89506# 4.64e-21
C3457 XM1/a_n158_60430# XM2/a_n158_n92142# 4.64e-21
C3458 XM1/a_n100_n117731# XM4/w_n358_n132787# 0.013363f
C3459 XM2/a_100_n152770# XM3/a_n158_53990# 0.042864f
C3460 XM4/a_100_112006# m1_1634_n2388# 6.1e-20
C3461 XM1/a_n100_n126347# XM2/a_n158_n279298# 0.005074f
C3462 XM1/a_n100_94797# XM2/a_100_n60510# 7.26e-20
C3463 XM1/a_100_47506# XM3/a_n158_98538# 0.001891f
C3464 XM4/w_n358_n132787# XM4/a_n100_38353# -0.004445f
C3465 XM1/a_n158_n54450# XM2/a_n158_n208126# 9.28e-21
C3466 XM2/a_100_n194946# XM3/a_n158_11514# 0.072074f
C3467 XM1/a_n100_66077# XM2/a_100_n86870# 7.26e-20
C3468 XM3/a_n100_n68355# m1_1634_n2388# 0.072015f
C3469 XM1/a_n158_92022# XM2/a_n158_n60510# 4.64e-21
C3470 XM4/w_n358_n132787# XM2/a_100_n81598# 0.106201f
C3471 XM1/a_n100_48845# XM4/w_n358_n132787# 0.013538f
C3472 XM1/a_100_n97530# XM2/a_n100_n250399# 0.005074f
C3473 XM2/a_100_n200218# m1_1634_n2388# 0.017213f
C3474 XM4/a_n100_n127407# m1_1634_n2388# 0.072015f
C3475 XM4/w_n358_n132787# XM2/a_n158_n268754# 0.107093f
C3476 XM2/a_100_n255574# XM3/a_n158_n50646# 0.077916f
C3477 XM1/a_n100_n89011# XM4/w_n358_n132787# 0.01311f
C3478 XM3/a_n100_41461# XM4/a_n100_41461# 0.009521f
C3479 XM3/a_n158_79890# m1_1634_n2388# 6.1e-20
C3480 XM1/a_n100_n47367# XM2/a_n158_n200218# 0.005074f
C3481 XM1/a_100_n166458# XM3/a_n100_n116011# 2.85e-20
C3482 XM2/a_100_n297750# XM3/a_n100_n92183# 0.010147f
C3483 XM2/a_n100_n295211# XM3/a_n158_n91050# 0.005074f
C3484 XM1/a_n100_n90447# m1_1634_n2388# 1.3e-19
C3485 XM4/w_n358_n132787# XM4/a_n100_n33131# -0.004445f
C3486 XM3/a_n158_24982# m1_1634_n2388# 6.1e-20
C3487 XM1/a_100_63302# XM2/a_n100_n89603# 0.005074f
C3488 XM2/a_n158_n208126# XM3/a_n100_n4123# 7.26e-20
C3489 XM3/a_n158_n4026# m1_1634_n2388# 6.1e-20
C3490 XM1/a_100_5862# XM4/w_n358_n132787# 0.054688f
C3491 XM2/a_n100_n337387# XM3/a_n100_n132587# 0.006572f
C3492 XM4/a_100_72638# m1_1634_n2388# 6.1e-20
C3493 XM1/a_100_n44398# XM4/w_n358_n132787# 0.05469f
C3494 XM1/a_n100_57461# XM3/a_n158_107862# 1.09e-21
C3495 XM1/a_100_n114762# XM2/a_n158_n268754# 0.116862f
C3496 XM1/a_n158_116434# XM2/a_n100_n39519# 7.26e-20
C3497 XM2/a_n158_n136954# XM3/a_n158_67458# 4.64e-21
C3498 XM1/a_n100_28741# m1_1634_n2388# 1.3e-19
C3499 XM2/a_n158_n292478# XM3/a_n158_n85870# 4.64e-21
C3500 XM1/a_n158_n75990# XM3/a_n100_n23807# 1.94e-20
C3501 XM3/a_n100_n107723# m1_1634_n2388# 0.072015f
C3502 XM1/a_n158_40326# XM2/a_n100_n113327# 3.69e-20
C3503 XM1/a_n100_n163683# XM2/a_100_n316202# 7.26e-20
C3504 XM2/a_n158_n179130# XM3/a_n158_24982# 4.64e-21
C3505 XM2/a_100_29114# XM4/w_n358_n132787# -5.68e-32
C3506 XM1/a_n100_n111987# m1_1634_n2388# 1.3e-19
C3507 XM2/a_n100_n139687# m1_1634_n2388# 0.001772f
C3508 XM1/a_100_n98966# XM3/a_n100_n46599# 1.05e-20
C3509 XM4/w_n358_n132787# XM2/a_100_n205490# 0.103342f
C3510 XM2/a_n158_n200218# XM3/a_n100_6237# 7.26e-20
C3511 XM1/a_n100_n10031# XM2/a_100_n165950# 6.06e-20
C3512 XM2/a_n158_n13062# XM1/a_100_140846# 0.116862f
C3513 XM2/a_n158_n15698# XM1/a_n100_139313# 0.005074f
C3514 XM2/a_100_n324110# m1_1634_n2388# 0.025819f
C3515 XM1/a_n100_n104807# XM2/a_n158_n258210# 0.005074f
C3516 XM4/w_n358_n132787# XM3/a_n100_n13447# 0.009017f
C3517 XM1/a_100_74790# XM3/a_n100_125377# 2.85e-20
C3518 XM1/a_n100_56025# XM3/a_n158_106826# 0.001667f
C3519 XM1/a_n158_37454# XM2/a_n100_n118599# 7.26e-20
C3520 XM4/w_n358_n132787# XM4/a_n100_n72499# -0.004445f
C3521 XM1/a_n158_21658# XM3/a_n100_73577# 1.94e-20
C3522 XM3/a_n158_n43394# m1_1634_n2388# 6.1e-20
C3523 XM4/a_100_33270# m1_1634_n2388# 6.1e-20
C3524 XM1/a_n158_153770# XM2/a_n158_118# 9.28e-21
C3525 XM1/a_n100_n134963# m1_1634_n2388# 8.95e-20
C3526 XM2/a_100_n237122# XM3/a_n158_n33034# 0.008591f
C3527 XM1/a_n158_n37218# XM3/a_n100_14525# 1.94e-20
C3528 XM2/a_n100_n242491# XM4/a_100_n38214# 2.56e-20
C3529 XM1/a_n158_18786# XM3/a_n100_69433# 1.36e-20
C3530 XM1/a_n100_14381# XM3/a_n158_65386# 2.85e-20
C3531 XM2/a_100_n279298# XM3/a_n100_n74571# 0.005563f
C3532 XM1/a_n100_n81831# XM4/w_n358_n132787# 0.01363f
C3533 XM1/a_n158_n53014# XM2/a_n158_n205490# 4.64e-21
C3534 XM1/a_100_64738# XM4/w_n358_n132787# 0.048442f
C3535 XM2/a_n158_n10426# XM1/a_n100_145057# 0.005074f
C3536 XM2/a_n100_n100147# XM3/a_n158_106826# 0.005074f
C3537 XM2/a_n158_n100050# XM3/a_n100_106729# 7.26e-20
C3538 XM1/a_100_31710# XM2/a_n100_n123871# 0.005074f
C3539 XM1/a_100_146590# XM2/a_n158_n7790# 0.116862f
C3540 XM2/a_n100_n318935# XM3/a_n100_n114975# 0.001243f
C3541 XM1/a_100_n113326# XM2/a_n158_n266118# 0.03819f
C3542 XM1/a_n100_n165119# XM3/a_n158_n112806# 2.85e-20
C3543 XM1/a_n158_n31474# XM3/a_n100_19705# 3.47e-20
C3544 XM1/a_100_28838# XM2/a_n100_n126507# 0.005074f
C3545 XM2/a_n158_n76326# m1_1634_n2388# 2.36e-21
C3546 XM4/a_n100_96369# m1_1634_n2388# 0.072015f
C3547 XM4/w_n358_n132787# XM3/a_n100_90153# 0.009186f
C3548 XM2/a_n100_n129143# XM4/a_100_75746# 2.11e-21
C3549 XM4/w_n358_n132787# XM3/a_n100_n52815# 0.009186f
C3550 XM4/a_100_n38214# m1_1634_n2388# 6.1e-20
C3551 XM1/a_n158_24530# XM2/a_n100_n129143# 1.8e-20
C3552 XM1/a_n100_11509# m1_1634_n2388# 1.3e-19
C3553 XM4/w_n358_n132787# XM2/a_n100_n144959# 0.02472f
C3554 XM2/a_n158_n316202# XM3/a_n100_n109795# 7.26e-20
C3555 XM1/a_n100_n113423# XM3/a_n158_n61006# 2.85e-20
C3556 XM2/a_n100_n263579# m1_1634_n2388# 7.61e-19
C3557 XM1/a_n158_n87478# XM3/a_n158_n35106# 1.14e-21
C3558 XM4/w_n358_n132787# XM3/a_n100_35245# 0.008249f
C3559 XM4/w_n358_n132787# XM4/a_n100_n111867# -0.004445f
C3560 XM3/a_n158_n82762# m1_1634_n2388# 6.1e-20
C3561 XM1/a_n100_60333# XM4/w_n358_n132787# 0.013481f
C3562 XM4/w_n358_n132787# XM2/a_100_n329382# 0.106052f
C3563 XM4/w_n358_n132787# XM1/a_100_n154970# 0.055165f
C3564 XM1/a_n158_n51578# XM2/a_n158_n205490# 9.28e-21
C3565 XM2/a_100_n202854# XM3/a_n100_1057# 0.005074f
C3566 XM1/a_100_71918# XM4/w_n358_n132787# 0.050159f
C3567 XM2/a_n158_n110594# XM3/a_n158_96466# 4.64e-21
C3568 XM1/a_n158_n40090# XM2/a_n158_n194946# 4.64e-21
C3569 XM2/a_100_n81598# XM3/a_n100_124341# 0.010147f
C3570 XM2/a_n158_n34150# XM4/w_n358_n132787# 0.101988f
C3571 XM1/a_n158_66174# XM2/a_n100_n89603# 7.26e-20
C3572 XM1/a_n100_124953# XM4/w_n358_n132787# 0.012279f
C3573 XM1/a_n158_60430# XM2/a_n100_n92239# 7.26e-20
C3574 XM1/a_n100_n169427# XM2/a_100_n324110# 8.75e-20
C3575 XM1/a_n100_n119167# XM2/a_100_n271390# 1.67e-20
C3576 XM2/a_n158_n152770# XM3/a_n158_53990# 4.64e-21
C3577 XM4/a_n100_57001# m1_1634_n2388# 0.072015f
C3578 XM2/a_100_n260846# XM3/a_n100_n56959# 0.004756f
C3579 XM1/a_n158_n182254# pcbias 0.011931f
C3580 XM4/w_n358_n132787# XM3/a_n100_n92183# 0.009186f
C3581 XM4/a_100_n77582# m1_1634_n2388# 6.1e-20
C3582 XM3/a_n100_9345# XM4/a_n100_9345# 0.009521f
C3583 XM3/a_n100_94297# XM4/a_n100_94297# 0.009521f
C3584 XM1/a_100_92022# XM2/a_n158_n63146# 0.081031f
C3585 XM1/a_n100_n172299# XM3/a_n158_n121094# 2.79e-20
C3586 XM2/a_n158_n194946# XM3/a_n158_11514# 4.64e-21
C3587 XM1/a_n100_66077# XM2/a_n158_n86870# 0.005074f
C3588 XM3/a_n100_73577# m1_1634_n2388# 0.072015f
C3589 XM3/a_n158_n122130# m1_1634_n2388# 6.1e-20
C3590 XM1/a_n100_n81831# XM2/a_100_n234486# 7.26e-20
C3591 XM4/w_n358_n132787# XM2/a_n158_n81598# 0.101988f
C3592 XM1/a_100_n183690# XM3/a_n100_n131551# 2.85e-20
C3593 XM1/a_100_n134866# XM2/a_n100_n287303# 0.002589f
C3594 XM1/a_100_129358# XM2/a_n158_n26242# 0.038969f
C3595 XM1/a_n100_n55983# XM2/a_n100_n208223# 0.002453f
C3596 XM3/a_n100_18669# m1_1634_n2388# 0.072015f
C3597 XM4/w_n358_n132787# XM2/a_n100_n268851# 0.025738f
C3598 XM1/a_100_89150# XM4/w_n358_n132787# 0.051635f
C3599 XM2/a_n100_n110691# XM4/a_100_93358# 1.29e-20
C3600 XM3/a_n158_114078# m1_1634_n2388# 6.1e-20
C3601 XM4/a_n100_n14483# m1_1634_n2388# 0.072015f
C3602 XM2/a_n158_n297750# XM3/a_n100_n92183# 1.45e-19
C3603 XM4/w_n358_n132787# XM3/a_n158_n27854# 0.038367f
C3604 XM4/w_n358_n132787# XM3/a_n158_60206# 0.032295f
C3605 XM1/a_n158_n119070# XM2/a_n100_n271487# 1.67e-20
C3606 XM4/a_n100_17633# m1_1634_n2388# 0.072015f
C3607 XM2/a_n158_13298# XM4/w_n358_n132787# 0.101988f
C3608 XM1/a_n100_2893# XM2/a_100_n152770# 7.26e-20
C3609 XM1/a_n100_57461# XM3/a_n100_107765# 0.001249f
C3610 XM1/a_n100_44537# XM2/a_100_n107958# 7.26e-20
C3611 XM4/w_n358_n132787# XM3/a_n100_n131551# 0.009186f
C3612 XM4/a_100_n116950# m1_1634_n2388# 6.1e-20
C3613 XM4/w_n358_n132787# XM1/a_n100_n140707# 0.013423f
C3614 XM1/a_n158_n65938# XM2/a_n158_n221306# 4.64e-21
C3615 XM2/a_n100_n137051# XM3/a_n158_67458# 0.005074f
C3616 XM2/a_n100_n292575# XM3/a_n158_n85870# 0.005074f
C3617 XM3/a_n100_21# m1_1634_n2388# 0.072015f
C3618 XM1/a_100_83406# XM2/a_n158_n71054# 0.116862f
C3619 XM4/w_n358_n132787# XM1/a_n100_145057# 0.012279f
C3620 XM3/a_n100_120197# XM4/a_n100_120197# 0.009521f
C3621 XM2/a_n100_n334751# XM3/a_n100_n127407# 0.004186f
C3622 XM1/a_n100_n163683# XM2/a_n158_n316202# 0.005074f
C3623 XM2/a_n100_n179227# XM3/a_n158_24982# 0.005074f
C3624 XM1/a_n158_n25730# XM3/a_n100_25921# 1.94e-20
C3625 XM1/a_100_n34346# m1_1634_n2388# 0.001456f
C3626 XM4/w_n358_n132787# XM4/a_n100_111909# -0.004445f
C3627 XM1/a_n158_24530# XM3/a_n100_76685# 1.94e-20
C3628 XM2/a_100_n136954# m1_1634_n2388# 0.017213f
C3629 XM1/a_n100_73257# XM3/a_n158_124438# 2.85e-20
C3630 XM4/w_n358_n132787# XM2/a_n158_n205490# 0.107093f
C3631 XM1/a_n100_n10031# XM2/a_n158_n165950# 0.004756f
C3632 XM2/a_n100_n18431# XM1/a_n158_135102# 7.26e-20
C3633 XM1/a_n100_50281# XM3/a_n100_100513# 2.08e-19
C3634 XM3/a_n158_98538# m1_1634_n2388# 6.1e-20
C3635 XM4/w_n358_n132787# XM3/a_n158_n67222# 0.038551f
C3636 XM4/a_n100_n53851# m1_1634_n2388# 0.072015f
C3637 XM1/a_100_n65938# XM2/a_100_n221306# 4.64e-21
C3638 XM1/a_100_21658# XM3/a_n100_72541# 2.85e-20
C3639 XM2/a_100_n326746# XM3/a_n158_n121094# 0.077916f
C3640 XM1/a_n158_n126250# XM3/a_n100_n75607# 4.81e-21
C3641 XM1/a_100_n68810# XM3/a_n100_n17591# 0.001743f
C3642 XM1/a_n158_76226# XM3/a_n100_127449# 2.89e-20
C3643 XM1/a_n100_173777# XM2/a_100_21206# 7.26e-20
C3644 XM4/w_n358_n132787# XM3/a_n158_112006# 0.038462f
C3645 XM3/a_n158_43630# m1_1634_n2388# 6.1e-20
C3646 XM2/a_n158_n237122# XM3/a_n158_n33034# 4.64e-21
C3647 XM1/a_n100_34485# XM2/a_100_n118502# 7.26e-20
C3648 XM1/a_100_14478# XM3/a_n100_66325# 2.85e-20
C3649 XM2/a_n158_n279298# XM3/a_n100_n74571# 9.05e-20
C3650 XM4/a_n100_8309# m1_1634_n2388# 0.072015f
C3651 XM1/a_n100_73257# XM4/w_n358_n132787# 0.0129f
C3652 XM1/a_n158_n53014# XM2/a_n100_n205587# 7.26e-20
C3653 XM1/a_n100_n18647# XM3/a_n158_32234# 2.85e-20
C3654 XM2/a_100_n97414# XM3/a_n158_106826# 0.023391f
C3655 XM1/a_n100_48845# XM3/a_n158_100610# 2.08e-20
C3656 XM1/a_100_31710# XM2/a_100_n121138# 4.64e-21
C3657 XM1/a_n158_74790# XM3/a_n100_125377# 1.94e-20
C3658 XM2/a_100_n234486# XM3/a_n158_n27854# 0.055327f
C3659 XM4/w_n358_n132787# XM4/a_n100_72541# -0.004445f
C3660 XM1/a_100_n113326# XM2/a_n100_n266215# 0.005074f
C3661 XM1/a_n100_n87575# XM3/a_n158_n35106# 4.65e-19
C3662 XM2/a_n100_n239855# XM4/a_100_n33034# 2.56e-20
C3663 XM1/a_100_n5626# XM3/a_n100_46641# 8.56e-19
C3664 XM3/a_n100_n34167# m1_1634_n2388# 0.072015f
C3665 XM1/a_n100_n37315# XM2/a_100_n189674# 7.26e-20
C3666 XM1/a_100_n18550# XM3/a_n100_32137# 2.85e-20
C3667 XM1/a_100_102074# XM2/a_n158_n52602# 0.116862f
C3668 XM1/a_100_28838# XM2/a_100_n123774# 4.64e-21
C3669 XM1/a_n158_n136302# XM3/a_n100_n84931# 3.89e-20
C3670 XM2/a_n100_n76423# m1_1634_n2388# 9.92e-19
C3671 XM4/w_n358_n132787# XM3/a_n158_n106590# 0.038462f
C3672 XM4/a_n100_n93219# m1_1634_n2388# 0.072015f
C3673 XM4/w_n358_n132787# XM2/a_100_n142226# 0.103342f
C3674 XM2/a_100_n260846# m1_1634_n2388# 0.024866f
C3675 XM1/a_n158_n104710# XM3/a_n100_n53851# 1.94e-20
C3676 XM1/a_n100_n123475# XM2/a_100_n279298# 7.26e-20
C3677 XM2/a_100_n113230# XM3/a_n100_91189# 0.005074f
C3678 XM4/w_n358_n132787# XM2/a_n158_n329382# 0.107093f
C3679 XM1/a_100_n103274# m1_1634_n2388# 2.44e-19
C3680 XM3/a_n100_103621# XM4/a_n100_103621# 0.009521f
C3681 XM2/a_n158_n202854# XM3/a_n100_1057# 7.26e-20
C3682 XM2/a_n100_n50063# XM4/w_n358_n132787# 0.012279f
C3683 XM2/a_100_n155406# XM3/a_n100_48713# 0.005074f
C3684 XM4/a_100_106826# m1_1634_n2388# 6.1e-20
C3685 XM3/a_n100_62181# XM4/a_n100_62181# 0.009521f
C3686 XM2/a_100_n308294# XM3/a_n158_n103482# 0.077916f
C3687 XM2/a_n100_n110691# XM3/a_n158_96466# 0.005074f
C3688 XM1/a_n100_7201# m1_1634_n2388# 6.74e-20
C3689 XM1/a_n158_n40090# XM2/a_n100_n195043# 4.59e-20
C3690 XM4/w_n358_n132787# XM4/a_n100_33173# -0.004445f
C3691 XM2/a_n158_n81598# XM3/a_n100_124341# 1.45e-19
C3692 XM3/a_n100_n73535# m1_1634_n2388# 0.072014f
C3693 XM1/a_n100_n169427# XM2/a_n158_n324110# 0.005482f
C3694 XM1/a_n100_n119167# XM2/a_n158_n271390# 8.32e-19
C3695 XM1/a_100_n24294# XM2/a_100_n179130# 4.64e-21
C3696 XM2/a_n100_n152867# XM3/a_n158_53990# 0.005074f
C3697 XM1/a_n100_n178043# m1_1634_n2388# 1.13e-19
C3698 XM2/a_n158_n260846# XM3/a_n100_n56959# 6.06e-20
C3699 XM1/a_n158_56122# XM2/a_n158_n97414# 4.64e-21
C3700 XM3/a_n100_n18627# XM4/a_n100_n18627# 0.009521f
C3701 XM1/a_100_130794# XM2/a_n158_n23606# 0.116862f
C3702 XM1/a_n158_n18550# XM2/a_n158_n173858# 4.64e-21
C3703 XM2/a_n100_n195043# XM3/a_n158_11514# 0.002512f
C3704 XM1/a_100_n123378# XM3/a_n100_n72499# 2.85e-20
C3705 XM1/a_n100_n81831# XM2/a_n158_n234486# 0.005074f
C3706 XM2/a_100_n216034# XM3/a_n158_n10242# 0.077916f
C3707 XM4/w_n358_n132787# XM2/a_n100_n81695# 0.024817f
C3708 XM1/a_n158_8734# XM2/a_n158_n144862# 4.64e-21
C3709 XM1/a_n100_n153631# XM2/a_100_n308294# 1.05e-19
C3710 XM2/a_n100_n200315# m1_1634_n2388# 7.61e-19
C3711 XM1/a_n100_n12903# m1_1634_n2388# 9.78e-20
C3712 XM4/w_n358_n132787# XM3/a_n100_53893# 0.009071f
C3713 XM4/a_100_n130418# m1_1634_n2388# 6.1e-20
C3714 XM2/a_100_n258210# XM3/a_n100_n51779# 0.005074f
C3715 XM4/w_n358_n132787# XM4/a_n100_n38311# -0.004445f
C3716 XM4/w_n358_n132787# XM2/a_100_n266118# 0.10657f
C3717 XM1/a_n158_n81734# XM2/a_n158_n237122# 4.64e-21
C3718 XM3/a_n158_n9206# m1_1634_n2388# 6.1e-20
C3719 XM1/a_n100_8637# XM4/w_n358_n132787# 0.011718f
C3720 XM3/a_n100_113981# m1_1634_n2388# 0.072015f
C3721 XM4/a_100_67458# m1_1634_n2388# 6.1e-20
C3722 XM1/a_100_n165022# XM3/a_n100_n113939# 2.85e-20
C3723 XM1/a_100_n136302# XM2/a_100_n289842# 4.64e-21
C3724 XM1/a_n158_148026# XM2/a_n158_n5154# 4.64e-21
C3725 XM2/a_100_n142226# XM3/a_n100_63217# 0.010147f
C3726 XM1/a_n100_27305# m1_1634_n2388# 7.08e-20
C3727 XM1/a_n100_n126347# XM3/a_n158_n75510# 2.85e-20
C3728 XM3/a_n100_n112903# m1_1634_n2388# 0.072015f
C3729 XM2/a_n100_n108055# XM4/a_100_98538# 2.53e-20
C3730 XM2/a_100_n184402# XM3/a_n100_20741# 0.010147f
C3731 XM1/a_n158_n65938# XM2/a_n100_n221403# 7.26e-20
C3732 XM1/a_n100_2893# XM2/a_n158_n152770# 0.005074f
C3733 XM1/a_100_122178# XM2/a_n158_n31514# 0.116862f
C3734 XM1/a_n100_81873# XM2/a_n158_n73690# 0.005074f
C3735 XM1/a_n100_44537# XM2/a_n158_n107958# 0.005074f
C3736 XM3/a_n100_n38311# XM4/a_n100_n38311# 0.009521f
C3737 XM1/a_n100_27305# XM3/a_n100_79793# 0.001145f
C3738 XM2/a_n100_n295211# XM4/a_100_n91050# 2.56e-20
C3739 XM4/a_n100_130557# m1_1634_n2388# 0.072015f
C3740 XM1/a_100_n119070# XM3/a_n100_n68355# 2.85e-20
C3741 XM4/w_n358_n132787# XM3/a_n100_n18627# 0.009026f
C3742 XM4/a_100_n4026# m1_1634_n2388# 6.1e-20
C3743 XM1/a_n100_120645# XM2/a_n100_n31611# 0.004186f
C3744 XM3/a_n100_92225# m1_1634_n2388# 0.072015f
C3745 XM2/a_100_n332018# XM3/a_n100_n127407# 0.005074f
C3746 XM1/a_100_24530# XM3/a_n100_75649# 9.2e-20
C3747 XM1/a_n100_n24391# XM3/a_n158_28090# 0.001368f
C3748 XM4/w_n358_n132787# XM4/a_n100_n77679# -0.004445f
C3749 XM1/a_100_n40090# XM2/a_100_n194946# 4.64e-21
C3750 XM4/w_n358_n132787# XM1/a_n100_n152195# 0.014098f
C3751 XM1/a_100_n126250# XM2/a_100_n281934# 4.64e-21
C3752 XM3/a_n158_n48574# m1_1634_n2388# 6.1e-20
C3753 XM1/a_n100_37357# XM4/w_n358_n132787# 0.01363f
C3754 XM4/a_100_28090# m1_1634_n2388# 6.1e-20
C3755 XM3/a_n100_37317# m1_1634_n2388# 0.072015f
C3756 XM4/w_n358_n132787# XM2/a_n100_n205587# 0.025738f
C3757 XM2/a_100_n197582# XM3/a_n100_6237# 4.8e-19
C3758 XM1/a_n100_n10031# XM2/a_n100_n166047# 4.97e-19
C3759 XM2/a_n100_n324207# m1_1634_n2388# 7.61e-19
C3760 XM1/a_100_n65938# XM2/a_n158_n221306# 0.061558f
C3761 XM2/a_n100_n181863# XM4/a_100_22910# 2.56e-20
C3762 XM1/a_n158_51814# XM3/a_n100_102585# 1.94e-20
C3763 XM1/a_n158_37454# XM2/a_n158_n115866# 4.64e-21
C3764 XM1/a_n158_n170766# XM3/a_n100_n119119# 1.94e-20
C3765 XM1/a_n158_n78862# XM3/a_n100_n26915# 1.94e-20
C3766 XM1/a_100_152334# XM4/w_n358_n132787# 0.049492f
C3767 XM4/w_n358_n132787# XM3/a_n158_78854# 0.032295f
C3768 XM2/a_100_n129046# XM3/a_n100_77721# 0.005074f
C3769 XM1/a_n158_n154970# XM2/a_n158_n310930# 4.64e-21
C3770 XM2/a_100_n239758# XM3/a_n100_n34167# 0.010147f
C3771 XM4/w_n358_n132787# XM3/a_n100_111909# 0.008953f
C3772 XM1/a_100_57558# XM3/a_n100_108801# 9.01e-20
C3773 XM1/a_n158_13042# XM3/a_n100_65289# 1.94e-20
C3774 XM2/a_n100_n237219# XM3/a_n158_n33034# 0.005074f
C3775 XM1/a_100_n78862# m1_1634_n2388# 1.22e-19
C3776 XM1/a_100_n68810# m1_1634_n2388# 5.46e-19
C3777 XM1/a_n158_50378# XM3/a_n100_101549# 3.31e-20
C3778 XM1/a_n100_34485# XM2/a_n158_n118502# 0.005074f
C3779 XM4/w_n358_n132787# XM3/a_n158_23946# 0.032295f
C3780 XM2/a_100_n171222# XM3/a_n100_35245# 0.005074f
C3781 XM2/a_n100_n279395# XM3/a_n100_n74571# 0.004501f
C3782 XM3/a_n100_n57995# XM4/a_n100_n57995# 0.009521f
C3783 XM1/a_100_n9934# XM4/w_n358_n132787# 0.054467f
C3784 XM1/a_100_107818# XM4/w_n358_n132787# 0.053546f
C3785 XM1/a_n100_n7159# XM3/a_n158_43630# 6.79e-19
C3786 XM4/a_n100_91189# m1_1634_n2388# 0.072014f
C3787 XM4/a_100_n43394# m1_1634_n2388# 6.1e-20
C3788 XM2/a_100_n97414# XM3/a_n100_106729# 0.005074f
C3789 XM2/a_n158_n97414# XM3/a_n158_106826# 4.64e-21
C3790 XM1/a_n100_48845# XM3/a_n100_100513# 3.77e-19
C3791 XM1/a_100_31710# XM2/a_n158_n121138# 0.043643f
C3792 XM4/w_n358_n132787# XM3/a_n100_n57995# 0.009065f
C3793 XM1/a_n100_18689# m1_1634_n2388# 1.3e-19
C3794 XM2/a_n158_n234486# XM3/a_n158_n27854# 4.64e-21
C3795 XM4/w_n358_n132787# XM4/a_n100_n117047# -0.004445f
C3796 XM1/a_n158_n7062# XM3/a_n100_43533# 1.94e-20
C3797 XM3/a_n158_n87942# m1_1634_n2388# 6.1e-20
C3798 XM1/a_n100_n37315# XM2/a_n158_n189674# 0.005074f
C3799 XM1/a_100_28838# XM2/a_n158_n123774# 0.020665f
C3800 XM1/a_100_n11370# XM3/a_n100_40425# 2.85e-20
C3801 XM3/a_n100_30065# XM4/a_n100_30065# 0.009521f
C3802 XM1/a_n100_n159375# XM3/a_n100_n107723# 5.85e-19
C3803 XM4/w_n358_n132787# XM2/a_n158_n142226# 0.107027f
C3804 XM2/a_n158_n260846# m1_1634_n2388# 2.36e-21
C3805 XM1/a_n100_n123475# XM2/a_n158_n279298# 0.005074f
C3806 XM1/a_n158_179618# XM2/a_n158_23842# 4.64e-21
C3807 XM2/a_n158_n113230# XM3/a_n100_91189# 7.26e-20
C3808 XM4/w_n358_n132787# XM2/a_n100_n329479# 0.024713f
C3809 XM1/a_100_n24294# m1_1634_n2388# 6.07e-19
C3810 XM3/a_n158_62278# m1_1634_n2388# 6.1e-20
C3811 XM1/a_n100_n150759# XM3/a_n100_n100471# 6.96e-19
C3812 XM3/a_n100_n77679# XM4/a_n100_n77679# 0.009521f
C3813 XM1/a_n100_133569# XM2/a_100_n20970# 1.45e-19
C3814 XM1/a_n100_123517# XM4/w_n358_n132787# 0.012279f
C3815 XM1/a_n100_20125# XM4/w_n358_n132787# 0.013401f
C3816 XM2/a_n158_n155406# XM3/a_n100_48713# 7.26e-20
C3817 XM4/a_n100_51821# m1_1634_n2388# 0.072015f
C3818 iout XM4/w_n358_n132787# 0.00293f
C3819 XM4/w_n358_n132787# XM3/a_n100_n97363# 0.009186f
C3820 XM4/a_100_n82762# m1_1634_n2388# 6.1e-20
C3821 XM2/a_100_n107958# XM3/a_n158_96466# 0.041306f
C3822 XM2/a_100_n221306# XM3/a_n100_n16555# 0.006531f
C3823 XM1/a_100_n50142# XM2/a_100_n205490# 4.64e-21
C3824 XM1/a_100_176746# XM4/w_n358_n132787# 0.053546f
C3825 XM2/a_100_n81598# XM3/a_n158_125474# 0.012486f
C3826 XM1/a_n100_41665# m1_1634_n2388# 1.41e-19
C3827 XM1/a_100_n106146# XM3/a_n100_n53851# 2.85e-20
C3828 XM1/a_100_n47270# XM4/w_n358_n132787# 0.054609f
C3829 XM1/a_n158_66174# XM2/a_n158_n86870# 4.64e-21
C3830 XM3/a_n158_n127310# m1_1634_n2388# 6.1e-20
C3831 XM1/a_100_n24294# XM2/a_n158_n179130# 0.113357f
C3832 XM1/a_n100_n169427# XM2/a_n100_n324207# 0.004872f
C3833 XM1/a_n100_n119167# XM2/a_n100_n271487# 0.003705f
C3834 XM2/a_100_n150134# XM3/a_n158_53990# 0.012096f
C3835 XM1/a_n158_n183690# iout_n 0.011231f
C3836 XM2/a_n100_n260943# XM3/a_n100_n56959# 4.97e-19
C3837 XM1/a_n158_56122# XM2/a_n100_n97511# 5.19e-20
C3838 XM1/a_n158_n18550# XM2/a_n100_n173955# 7.26e-20
C3839 XM4/w_n358_n132787# XM3/a_n158_n33034# 0.038462f
C3840 XM4/a_n100_n19663# m1_1634_n2388# 0.072015f
C3841 XM1/a_100_81970# XM2/a_n100_n73787# 0.005074f
C3842 XM4/w_n358_n132787# XM2/a_100_n78962# 0.103341f
C3843 XM1/a_n158_8734# XM2/a_n100_n144959# 2.99e-21
C3844 XM1/a_n100_n153631# XM2/a_n158_n308294# 0.005892f
C3845 XM2/a_100_n197582# m1_1634_n2388# 0.023368f
C3846 XM1/a_100_118# m1_1634_n2388# 0.002244f
C3847 XM1/a_n100_38793# XM3/a_n100_89117# 9.89e-19
C3848 XM2/a_n158_n258210# XM3/a_n100_n51779# 7.26e-20
C3849 XM1/a_n100_129261# XM2/a_100_n23606# 7.26e-20
C3850 XM1/a_n100_119209# XM2/a_n100_n36883# 0.004759f
C3851 XM1/a_n158_n106146# XM3/a_n100_n53851# 1.94e-20
C3852 XM1/a_100_44634# XM3/a_n158_96466# 0.00544f
C3853 XM3/a_n100_n97363# XM4/a_n100_n97363# 0.009521f
C3854 XM4/w_n358_n132787# XM2/a_n158_n266118# 0.107093f
C3855 XM1/a_n158_n81734# XM2/a_n100_n237219# 7.26e-20
C3856 XM1/a_100_123614# XM2/a_100_n28878# 4.64e-21
C3857 XM4/a_n100_12453# m1_1634_n2388# 0.072015f
C3858 XM2/a_n100_n2615# XM4/w_n358_n132787# 0.01231f
C3859 XM1/a_100_87714# XM2/a_n158_n65782# 0.106736f
C3860 XM4/a_100_n122130# m1_1634_n2388# 6.1e-20
C3861 XM1/a_100_n136302# XM2/a_n158_n289842# 0.11102f
C3862 XM2/a_n158_n142226# XM3/a_n100_63217# 1.45e-19
C3863 XM1/a_n100_n109115# XM4/w_n358_n132787# 0.013576f
C3864 XM2/a_100_n208126# XM3/a_n100_n3087# 0.010147f
C3865 XM4/w_n358_n132787# XM3/a_n100_5201# 0.009103f
C3866 XM2/a_n158_n184402# XM3/a_n100_20741# 1.45e-19
C3867 XM1/a_n158_n24294# XM2/a_n158_n179130# 4.64e-21
C3868 XM1/a_n100_37357# XM3/a_n158_88178# 2.85e-20
C3869 XM4/w_n358_n132787# XM4/a_n100_106729# -0.004445f
C3870 XM2/a_100_n136954# XM3/a_n158_68494# 0.077916f
C3871 XM1/a_n158_n53014# XM3/a_n100_n1015# 1.78e-20
C3872 XM1/a_n100_n100499# XM4/w_n358_n132787# 0.01363f
C3873 XM4/a_n100_n59031# m1_1634_n2388# 0.072015f
C3874 XM2/a_100_n202854# XM3/a_n158_2190# 0.077916f
C3875 XM1/a_n158_n32910# XM3/a_n100_17633# 1.94e-20
C3876 XM1/a_100_n19986# XM3/a_n100_31101# 2.85e-20
C3877 XM2/a_n158_n332018# XM3/a_n100_n127407# 7.26e-20
C3878 XM4/w_n358_n132787# XM3/a_n158_n72402# 0.038462f
C3879 XM2/a_100_n179130# XM3/a_n158_26018# 0.077916f
C3880 XM1/a_n100_n172299# XM4/w_n358_n132787# 0.013614f
C3881 XM1/a_100_n40090# XM2/a_n158_n194946# 0.111409f
C3882 XM4/w_n358_n132787# XM3/a_n100_72541# 0.009135f
C3883 XM2/a_n100_n137051# m1_1634_n2388# 9.65e-19
C3884 XM3/a_n100_n117047# XM4/a_n100_n117047# 0.009521f
C3885 XM2/a_100_n287206# XM3/a_n158_n80690# 0.066621f
C3886 XM1/a_100_n126250# XM2/a_n158_n281934# 0.030791f
C3887 XM2/a_n100_n292575# XM4/a_100_n85870# 2.56e-20
C3888 XM1/a_100_176746# XM2/a_n100_21109# 0.005074f
C3889 XM2/a_100_n329382# XM3/a_n100_n122227# 0.003292f
C3890 XM4/w_n358_n132787# XM2/a_100_n202854# 0.10657f
C3891 XM2/a_n158_n197582# XM3/a_n100_6237# 1.37e-20
C3892 XM1/a_n100_n10031# XM2/a_100_n163314# 7.26e-20
C3893 XM2/a_n158_26478# XM1/a_100_181054# 0.116862f
C3894 XM2/a_100_n321474# m1_1634_n2388# 0.017213f
C3895 XM1/a_n100_n140707# XM2/a_100_n295114# 1.45e-19
C3896 XM1/a_100_n65938# XM2/a_n100_n221403# 0.005074f
C3897 XM4/w_n358_n132787# XM3/a_n100_17633# 0.009559f
C3898 XM1/a_100_149462# XM2/a_n158_n5154# 0.116862f
C3899 XM1/a_n100_79001# XM4/w_n358_n132787# 0.013474f
C3900 XM1/a_100_74790# XM3/a_n100_126413# 2.85e-20
C3901 XM1/a_n100_56025# XM3/a_n158_107862# 2.85e-20
C3902 XM1/a_n158_37454# XM2/a_n100_n115963# 7.26e-20
C3903 XM1/a_100_n123378# XM4/w_n358_n132787# 0.054609f
C3904 XM1/a_n100_n18647# XM2/a_100_n173858# 7.26e-20
C3905 XM1/a_n100_n8595# XM3/a_n158_43630# 7.19e-19
C3906 XM2/a_n158_n129046# XM3/a_n100_77721# 7.26e-20
C3907 XM1/a_100_13042# XM3/a_n100_64253# 8.1e-19
C3908 XM1/a_n158_n154970# XM2/a_n100_n311027# 7.26e-20
C3909 XM2/a_n158_n239758# XM3/a_n100_n34167# 1.45e-19
C3910 XM1/a_n158_n51578# XM3/a_n100_n1015# 1.94e-20
C3911 XM4/w_n358_n132787# XM4/a_n100_67361# -0.004445f
C3912 XM1/a_n158_n97530# XM3/a_n100_n46599# 7.21e-21
C3913 XM2/a_n158_n171222# XM3/a_n100_35245# 7.26e-20
C3914 XM1/a_n158_n144918# XM2/a_n158_n300386# 4.64e-21
C3915 XM3/a_n100_n39347# m1_1634_n2388# 0.072015f
C3916 XM2/a_n100_n179227# XM4/a_100_28090# 2.03e-20
C3917 XM1/a_n100_172341# XM2/a_n158_18570# 0.010147f
C3918 XM3/a_n100_82901# XM4/a_n100_82901# 0.009521f
C3919 XM2/a_100_n123774# XM3/a_n158_82998# 0.041696f
C3920 XM1/a_100_15914# XM3/a_n158_67458# 0.00544f
C3921 XM2/a_n158_n97414# XM3/a_n100_106729# 7.26e-20
C3922 XM2/a_n100_n97511# XM3/a_n158_106826# 0.005074f
C3923 XM1/a_100_31710# XM2/a_n100_n121235# 0.005074f
C3924 XM4/w_n358_n132787# XM3/a_n158_n111770# 0.038462f
C3925 XM4/a_n100_n98399# m1_1634_n2388# 0.072015f
C3926 XM2/a_n100_n234583# XM3/a_n158_n27854# 0.005074f
C3927 XM1/a_100_n88914# XM3/a_n158_n38214# 0.002797f
C3928 XM2/a_100_n165950# XM3/a_n158_40522# 0.070905f
C3929 XM2/a_n100_n276759# XM3/a_n100_n69391# 0.001586f
C3930 XM1/a_100_28838# XM2/a_n100_n123871# 0.005074f
C3931 XM1/a_100_n41526# XM2/a_n100_n197679# 0.002941f
C3932 XM1/a_100_24530# XM2/a_100_n129046# 4.64e-21
C3933 XM3/a_n100_55965# m1_1634_n2388# 0.072015f
C3934 XM4/w_n358_n132787# XM4/a_n100_n4123# -0.004445f
C3935 XM4/w_n358_n132787# XM2/a_n100_n142323# 0.025677f
C3936 XM2/a_n100_n260943# m1_1634_n2388# 8.39e-19
C3937 XM4/a_100_101646# m1_1634_n2388# 6.1e-20
C3938 XM3/a_n158_1154# m1_1634_n2388# 6.1e-20
C3939 XM1/a_n100_142185# XM2/a_n158_n10426# 0.005074f
C3940 XM4/w_n358_n132787# XM3/a_n158_97502# 0.032295f
C3941 XM4/w_n358_n132787# XM2/a_100_n326746# 0.103342f
C3942 XM2/a_100_n268754# XM3/a_n158_n63078# 0.077916f
C3943 XM4/w_n358_n132787# XM4/a_n100_27993# -0.004445f
C3944 XM2/a_100_n310930# XM3/a_n100_n104615# 0.005074f
C3945 XM3/a_n100_n78715# m1_1634_n2388# 0.072015f
C3946 XM4/w_n358_n132787# XM3/a_n158_42594# 0.032295f
C3947 XM2/a_n158_n107958# XM3/a_n158_96466# 4.64e-21
C3948 XM2/a_n158_n221306# XM3/a_n100_n16555# 1.12e-19
C3949 XM1/a_100_n50142# XM2/a_n158_n205490# 0.063506f
C3950 XM2/a_n158_n81598# XM3/a_n158_125474# 4.64e-21
C3951 XM2/a_100_n81598# XM3/a_n100_125377# 0.005074f
C3952 XM1/a_100_n124814# XM3/a_n100_n72499# 2.58e-20
C3953 XM1/a_100_n120506# XM4/w_n358_n132787# 0.050035f
C3954 XM1/a_n158_n113326# XM3/a_n100_n61103# 1.94e-20
C3955 XM1/a_n158_66174# XM2/a_n100_n86967# 7.26e-20
C3956 XM1/a_100_n24294# XM2/a_n100_n179227# 7.31e-19
C3957 XM2/a_n158_n150134# XM3/a_n158_53990# 4.64e-21
C3958 XM1/a_n100_94797# XM2/a_100_n57874# 7.26e-20
C3959 XM4/w_n358_n132787# XM4/a_n100_n43491# -0.004445f
C3960 XM3/a_n158_n14386# m1_1634_n2388# 6.1e-20
C3961 XM1/a_n158_51814# XM2/a_n158_n102686# 9.28e-21
C3962 XM4/a_100_62278# m1_1634_n2388# 6.1e-20
C3963 XM4/w_n358_n132787# XM2/a_n158_n78962# 0.105768f
C3964 XM1/a_n100_n153631# XM2/a_n100_n308391# 0.003018f
C3965 XM1/a_n100_34485# m1_1634_n2388# 1.02e-19
C3966 XM1/a_n100_n31571# XM4/w_n358_n132787# 0.013513f
C3967 XM1/a_n158_50378# XM2/a_n158_n105322# 4.64e-21
C3968 XM3/a_n100_n118083# m1_1634_n2388# 0.072015f
C3969 XM4/w_n358_n132787# XM2/a_n100_n266215# 0.025738f
C3970 XM3/a_n158_80926# m1_1634_n2388# 6.1e-20
C3971 XM1/a_100_n143482# XM3/a_n100_n93219# 1.76e-20
C3972 XM4/w_n358_n132787# XM3/a_n100_n1015# 0.009008f
C3973 XM3/a_n158_115114# m1_1634_n2388# 6.1e-20
C3974 XM1/a_n100_40229# XM3/a_n158_91286# 0.001634f
C3975 XM1/a_100_n136302# XM2/a_n100_n289939# 0.002512f
C3976 XM1/a_100_81970# XM4/w_n358_n132787# 0.053546f
C3977 XM3/a_n158_26018# m1_1634_n2388# 6.1e-20
C3978 XM4/a_n100_125377# m1_1634_n2388# 0.072015f
C3979 XM2/a_100_n250302# XM3/a_n158_n45466# 0.077916f
C3980 XM4/w_n358_n132787# XM3/a_n100_n23807# 0.009186f
C3981 XM4/a_100_n9206# m1_1634_n2388# 6.1e-20
C3982 XM2/a_n158_n208126# XM3/a_n100_n3087# 1.45e-19
C3983 XM1/a_n158_44634# XM2/a_n158_n110594# 4.64e-21
C3984 XM1/a_n158_n24294# XM2/a_n100_n179227# 2.69e-20
C3985 XM2/a_100_n292478# XM3/a_n100_n87003# 0.010147f
C3986 XM1/a_n158_n65938# XM2/a_n158_n218670# 4.64e-21
C3987 XM1/a_n100_2893# XM2/a_100_n150134# 7.26e-20
C3988 XM1/a_n158_116434# XM2/a_n100_n36883# 7.26e-20
C3989 XM4/w_n358_n132787# XM4/a_n100_n82859# -0.004445f
C3990 XM2/a_n100_n289939# XM3/a_n158_n85870# 0.004513f
C3991 XM3/a_n158_n53754# m1_1634_n2388# 6.1e-20
C3992 XM1/a_n100_83309# XM2/a_100_n71054# 1.45e-19
C3993 XM4/a_100_22910# m1_1634_n2388# 6.1e-20
C3994 XM1/a_100_34582# XM3/a_n100_84973# 2.85e-20
C3995 XM2/a_n100_n332115# XM3/a_n100_n127407# 7.77e-20
C3996 XM1/a_n158_n147790# XM3/a_n100_n97363# 1.94e-20
C3997 XM2/a_n158_26478# XM1/a_n100_180957# 0.010147f
C3998 XM1/a_100_n153534# XM3/a_n100_n101507# 2.85e-20
C3999 XM1/a_n158_n5626# XM2/a_n158_n160678# 4.64e-21
C4000 XM1/a_100_n40090# XM2/a_n100_n195043# 0.00216f
C4001 XM2/a_100_n134318# m1_1634_n2388# 0.019665f
C4002 XM2/a_n158_n287206# XM3/a_n158_n80690# 4.64e-21
C4003 XM1/a_100_n126250# XM2/a_n100_n282031# 0.005074f
C4004 XM1/a_n100_73257# XM3/a_n158_125474# 0.001477f
C4005 XM2/a_n158_n329382# XM3/a_n100_n122227# 3.76e-20
C4006 XM4/a_100_2190# m1_1634_n2388# 6.1e-20
C4007 XM4/w_n358_n132787# XM2/a_n158_n202854# 0.107093f
C4008 XM2/a_n100_n197679# XM3/a_n100_6237# 0.004047f
C4009 XM1/a_n100_n10031# XM2/a_n158_n163314# 0.005074f
C4010 XM2/a_n158_n13062# XM1/a_n100_139313# 0.005074f
C4011 XM1/a_n100_50281# XM3/a_n100_101549# 3.77e-19
C4012 XM1/a_n100_n140707# XM2/a_n158_n295114# 0.010147f
C4013 XM1/a_100_n65938# XM2/a_100_n218670# 4.64e-21
C4014 XM3/a_n100_50785# XM4/a_n100_50785# 0.009521f
C4015 XM1/a_n100_21561# XM3/a_n158_72638# 2.85e-20
C4016 XM1/a_n100_110593# XM2/a_n158_n44694# 0.005074f
C4017 XM1/a_n100_n18647# XM2/a_n158_n173858# 0.005074f
C4018 XM1/a_n158_76226# XM3/a_n100_128485# 1.94e-20
C4019 XM4/a_n100_86009# m1_1634_n2388# 0.072015f
C4020 XM4/w_n358_n132787# XM3/a_n100_n63175# 0.009093f
C4021 XM4/a_100_n48574# m1_1634_n2388# 6.1e-20
C4022 XM1/a_n100_142185# XM4/w_n358_n132787# 0.012279f
C4023 XM4/w_n358_n132787# XM3/a_n158_113042# 0.032295f
C4024 XM1/a_100_57558# XM3/a_n158_109934# 3.95e-20
C4025 XM1/a_n158_n167894# XM3/a_n100_n116011# 1.94e-20
C4026 XM1/a_100_n144918# m1_1634_n2388# 5.46e-19
C4027 XM4/w_n358_n132787# XM4/a_n100_n122227# -0.004445f
C4028 XM1/a_n158_18786# XM3/a_n100_70469# 1.68e-20
C4029 XM1/a_n100_14381# XM3/a_n158_66422# 2.85e-20
C4030 XM1/a_n100_5765# XM3/a_n100_57001# 7.93e-19
C4031 XM3/a_n158_n93122# m1_1634_n2388# 6.1e-20
C4032 XM1/a_n158_n144918# XM2/a_n100_n300483# 7.26e-20
C4033 XM1/a_n100_n70343# XM2/a_100_n223942# 1.44e-19
C4034 XM1/a_100_n70246# XM2/a_n158_n223942# 0.116862f
C4035 XM2/a_100_n73690# XM3/a_n158_130654# 0.033517f
C4036 XM2/a_n158_n123774# XM3/a_n158_82998# 4.64e-21
C4037 XM1/a_n100_n113423# m1_1634_n2388# 1.05e-19
C4038 XM2/a_n158_n7790# XM1/a_n100_145057# 0.005074f
C4039 XM2/a_100_n97414# XM3/a_n158_107862# 0.077916f
C4040 XM1/a_n158_74790# XM3/a_n100_126413# 1.94e-20
C4041 XM1/a_100_70482# XM4/w_n358_n132787# 0.048442f
C4042 XM1/a_100_n114762# XM3/a_n100_n63175# 2.85e-20
C4043 XM1/a_100_n97530# XM3/a_n100_n46599# 0.001364f
C4044 XM2/a_n100_n237219# XM4/a_100_n33034# 2.56e-20
C4045 XM1/a_n100_n77523# XM3/a_n158_n26818# 2.85e-20
C4046 XM2/a_n158_n165950# XM3/a_n158_40522# 4.64e-21
C4047 XM1/a_n100_n5723# XM3/a_n158_46738# 2.85e-20
C4048 XM2/a_100_n274026# XM3/a_n100_n69391# 0.005074f
C4049 XM1/a_n158_n31474# XM3/a_n100_20741# 1.94e-20
C4050 XM1/a_n100_n18647# XM4/w_n358_n132787# 0.01363f
C4051 XM4/w_n358_n132787# XM3/a_n100_91189# 0.009186f
C4052 XM1/a_n100_n93319# m1_1634_n2388# 1.3e-19
C4053 XM1/a_100_n41526# XM2/a_100_n194946# 4.64e-21
C4054 XM1/a_100_97766# XM2/a_100_n57874# 4.64e-21
C4055 XM1/a_100_24530# XM2/a_n158_n129046# 0.114525f
C4056 XM2/a_n100_n313663# XM3/a_n100_n109795# 0.004948f
C4057 XM4/w_n358_n132787# XM2/a_100_n139590# 0.105983f
C4058 XM2/a_100_n258210# m1_1634_n2388# 0.017213f
C4059 XM4/w_n358_n132787# XM3/a_n100_36281# 0.009186f
C4060 XM4/a_n100_46641# m1_1634_n2388# 0.072015f
C4061 XM4/a_100_n87942# m1_1634_n2388# 6.1e-20
C4062 XM1/a_n100_n123475# XM2/a_100_n276662# 7.26e-20
C4063 XM1/a_100_156642# XM2/a_n158_2754# 0.116862f
C4064 XM4/w_n358_n132787# XM1/a_100_n169330# 0.048442f
C4065 XM4/w_n358_n132787# XM3/a_n100_n102543# 0.008963f
C4066 XM2/a_n100_n123871# XM4/a_100_80926# 2.56e-20
C4067 XM4/w_n358_n132787# XM2/a_n158_n326746# 0.107093f
C4068 XM3/a_n158_n132490# m1_1634_n2388# 3.05e-20
C4069 XM2/a_n158_n310930# XM3/a_n100_n104615# 7.26e-20
C4070 XM1/a_n158_21658# XM2/a_n158_n134318# 4.64e-21
C4071 XM2/a_n100_n108055# XM3/a_n158_96466# 0.005074f
C4072 XM2/a_n100_n221403# XM3/a_n100_n16555# 0.002257f
C4073 XM1/a_100_n50142# XM2/a_n100_n205587# 0.005074f
C4074 XM2/a_n158_n81598# XM3/a_n100_125377# 7.26e-20
C4075 XM2/a_n100_n81695# XM3/a_n158_125474# 0.005074f
C4076 XM2/a_100_n197582# XM3/a_n158_7370# 0.077916f
C4077 XM1/a_n100_n28699# XM4/w_n358_n132787# 0.013484f
C4078 XM2/a_n158_n31514# XM4/w_n358_n132787# 0.103459f
C4079 XM1/a_n100_n142143# XM3/a_n158_n91050# 2.85e-20
C4080 XM4/w_n358_n132787# XM3/a_n158_n38214# 0.038943f
C4081 XM4/a_n100_n24843# m1_1634_n2388# 0.072015f
C4082 XM1/a_n158_n133430# XM2/a_n158_n287206# 9.28e-21
C4083 XM2/a_n100_n150231# XM3/a_n158_53990# 0.005074f
C4084 XM1/a_n100_50281# XM2/a_100_n105322# 7.26e-20
C4085 XM1/a_n158_15914# XM2/a_n158_n139590# 4.64e-21
C4086 XM1/a_n100_n34443# XM2/a_100_n189674# 7.26e-20
C4087 XM1/a_n158_n18550# XM2/a_n158_n171222# 4.64e-21
C4088 XM1/a_100_92022# XM2/a_n158_n60510# 0.012875f
C4089 XM3/a_n100_74613# m1_1634_n2388# 0.072015f
C4090 XM1/a_n100_n51675# XM3/a_n100_21# 1.3e-20
C4091 XM1/a_100_129358# XM2/a_n158_n23606# 0.054937f
C4092 XM4/w_n358_n132787# XM2/a_n100_n79059# 0.025318f
C4093 XM4/a_100_n127310# m1_1634_n2388# 6.1e-20
C4094 XM2/a_n100_n197679# m1_1634_n2388# 0.002699f
C4095 XM1/a_100_n157842# XM3/a_n100_n105651# 2.85e-20
C4096 XM3/a_n100_19705# m1_1634_n2388# 0.072015f
C4097 XM1/a_100_126486# XM2/a_n158_n28878# 0.061948f
C4098 XM1/a_n158_50378# XM2/a_n100_n105419# 7.26e-20
C4099 XM4/w_n358_n132787# XM2/a_100_n263482# 0.103341f
C4100 XM1/a_n158_n81734# XM2/a_n158_n234486# 4.64e-21
C4101 XM4/w_n358_n132787# XM1/a_100_140846# 0.048442f
C4102 XM3/a_n100_115017# m1_1634_n2388# 0.072015f
C4103 XM1/a_100_n57322# XM3/a_n100_n6195# 8.1e-20
C4104 XM4/w_n358_n132787# XM4/a_n100_101549# -0.004445f
C4105 XM3/a_n100_n5159# m1_1634_n2388# 0.072015f
C4106 XM4/w_n358_n132787# XM3/a_n158_61242# 0.032295f
C4107 XM1/a_100_119306# XM4/w_n358_n132787# 0.052075f
C4108 XM1/a_100_8734# XM4/w_n358_n132787# 0.048537f
C4109 XM1/a_n158_7298# XM2/a_n158_n147498# 9.28e-21
C4110 XM1/a_100_n77426# XM4/w_n358_n132787# 0.048442f
C4111 XM4/w_n358_n132787# XM3/a_n158_n77582# 0.038462f
C4112 XM4/a_n100_n64211# m1_1634_n2388# 0.072014f
C4113 XM1/a_n158_44634# XM2/a_n100_n110691# 7.26e-20
C4114 XM2/a_n158_15934# XM4/w_n358_n132787# 0.102727f
C4115 XM2/a_n158_n292478# XM3/a_n100_n87003# 1.45e-19
C4116 XM1/a_n158_n65938# XM2/a_n100_n218767# 7.26e-20
C4117 XM1/a_n100_2893# XM2/a_n158_n150134# 0.005074f
C4118 XM1/a_100_n117634# XM3/a_n100_n65247# 4.62e-21
C4119 XM1/a_100_n78862# XM3/a_n100_n27951# 4.32e-20
C4120 XM3/a_n100_18669# XM4/a_n100_18669# 0.009521f
C4121 XM1/a_n100_n30135# m1_1634_n2388# 1.3e-19
C4122 XM1/a_n158_28838# XM3/a_n100_79793# 1.94e-20
C4123 XM1/a_n158_n153534# XM3/a_n100_n102543# 1.94e-20
C4124 XM1/a_n158_n5626# XM2/a_n100_n160775# 7.26e-20
C4125 XM1/a_n158_n180818# XM3/a_n100_n130515# 1.94e-20
C4126 XM1/a_100_n173638# XM4/w_n358_n132787# 0.054711f
C4127 XM1/a_100_n149226# XM3/a_n100_n97363# 2.85e-20
C4128 XM1/a_100_n124814# XM4/w_n358_n132787# 0.048442f
C4129 XM2/a_n158_n134318# m1_1634_n2388# 5.91e-22
C4130 XM1/a_100_n172202# XM2/a_n158_n326746# 0.116862f
C4131 XM1/a_n100_n143579# XM3/a_n100_n91147# 4.16e-19
C4132 XM2/a_n100_n287303# XM3/a_n158_n80690# 0.005074f
C4133 XM1/a_100_n126250# XM2/a_100_n279298# 4.64e-21
C4134 XM2/a_n100_n329479# XM3/a_n100_n122227# 0.001959f
C4135 XM4/w_n358_n132787# XM2/a_n100_n202951# 0.025738f
C4136 XM3/a_n158_99574# m1_1634_n2388# 6.1e-20
C4137 XM4/w_n358_n132787# XM4/a_n100_62181# -0.004445f
C4138 XM2/a_n100_n321571# m1_1634_n2388# 7.61e-19
C4139 XM1/a_100_n94658# XM3/a_n100_n42455# 2.85e-20
C4140 XM1/a_100_n65938# XM2/a_n158_n218670# 0.032348f
C4141 XM1/a_100_21658# XM3/a_n100_73577# 2.85e-20
C4142 XM1/a_n158_n159278# XM2/a_n158_n313566# 9.28e-21
C4143 XM3/a_n100_n44527# m1_1634_n2388# 0.072015f
C4144 XM1/a_n158_51814# XM3/a_n100_103621# 1.94e-20
C4145 XM1/a_n100_31613# XM4/w_n358_n132787# 0.013551f
C4146 XM2/a_100_n126410# XM3/a_n100_77721# 0.005074f
C4147 XM1/a_n158_n154970# XM2/a_n158_n308294# 4.64e-21
C4148 XM4/a_n100_n103579# m1_1634_n2388# 0.072015f
C4149 XM3/a_n158_44666# m1_1634_n2388# 6.1e-20
C4150 XM4/w_n358_n132787# XM3/a_n100_112945# 0.009036f
C4151 XM1/a_100_57558# XM3/a_n100_109837# 8.96e-19
C4152 XM1/a_100_n170766# XM3/a_n158_n120058# 0.00544f
C4153 XM4/w_n358_n132787# XM3/a_n158_n116950# 0.039233f
C4154 XM3/a_n100_n4123# XM4/a_n100_n4123# 0.009521f
C4155 XM3/a_n100_127449# XM4/a_n100_127449# 0.009521f
C4156 XM1/a_100_53250# m1_1634_n2388# 0.004003f
C4157 XM1/a_100_n169330# XM3/a_n100_n117047# 2.85e-20
C4158 XM1/a_n158_50378# XM3/a_n100_102585# 1.94e-20
C4159 XM2/a_n100_n284667# XM4/a_n100_n80787# 2.06e-20
C4160 XM2/a_100_n168586# XM3/a_n100_35245# 0.001535f
C4161 XM2/a_100_n321474# XM3/a_n158_n115914# 0.077916f
C4162 XM1/a_n100_n70343# XM2/a_n158_n223942# 0.010128f
C4163 XM1/a_n158_176746# XM2/a_n100_21109# 7.26e-20
C4164 XM2/a_100_n73690# XM3/a_n100_130557# 0.005074f
C4165 XM1/a_n100_61769# m1_1634_n2388# 8.08e-20
C4166 XM2/a_n100_n123871# XM3/a_n158_82998# 0.005074f
C4167 XM1/a_n100_n101935# m1_1634_n2388# 7.01e-20
C4168 XM1/a_n100_n18647# XM3/a_n158_33270# 2.85e-20
C4169 XM2/a_100_n97414# XM3/a_n100_107765# 0.010147f
C4170 XM4/w_n358_n132787# XM4/a_n100_n9303# -0.004445f
C4171 XM1/a_100_n1318# XM3/a_n100_49749# 2.85e-20
C4172 XM1/a_n100_n165119# XM3/a_n100_n113939# 8.27e-19
C4173 XM2/a_n100_n166047# XM3/a_n158_40522# 0.003566f
C4174 XM4/a_100_96466# m1_1634_n2388# 6.1e-20
C4175 XM2/a_n158_n274026# XM3/a_n100_n69391# 7.26e-20
C4176 XM1/a_100_n18550# XM3/a_n100_33173# 2.85e-20
C4177 XM1/a_n100_168033# XM2/a_n100_13201# 0.003522f
C4178 XM1/a_100_n41526# XM2/a_n158_n194946# 0.099336f
C4179 XM4/w_n358_n132787# XM4/a_n100_22813# -0.004445f
C4180 XM1/a_100_24530# XM2/a_n100_n129143# 4.89e-19
C4181 XM1/a_n100_n113423# XM3/a_n100_n62139# 1.69e-19
C4182 XM1/a_n158_n94658# XM3/a_n100_n42455# 1.94e-20
C4183 XM1/a_n158_n87478# XM3/a_n100_n36239# 3.89e-20
C4184 XM3/a_n100_n83895# m1_1634_n2388# 0.072015f
C4185 XM2/a_100_n229214# XM3/a_n158_n22674# 0.064285f
C4186 XM4/w_n358_n132787# XM3/a_n158_6334# 0.036834f
C4187 XM1/a_n158_103510# XM2/a_n100_n50063# 7.26e-20
C4188 XM4/w_n358_n132787# XM2/a_n158_n139590# 0.107093f
C4189 XM2/a_n100_n234583# XM4/a_100_n27854# 2.56e-20
C4190 XM1/a_n100_n123475# XM2/a_n158_n276662# 0.005074f
C4191 XM2/a_100_n271390# XM3/a_n100_n64211# 0.001183f
C4192 XM3/a_n100_n23807# XM4/a_n100_n23807# 0.009521f
C4193 XM1/a_n100_70385# XM4/w_n358_n132787# 0.013405f
C4194 XM2/a_100_n113230# XM3/a_n100_92225# 0.010147f
C4195 XM4/w_n358_n132787# XM2/a_n100_n326843# 0.025738f
C4196 XM1/a_100_27402# XM2/a_n158_n126410# 0.116862f
C4197 XM4/w_n358_n132787# XM4/a_n100_2093# -0.004445f
C4198 XM2/a_n100_n47427# XM4/w_n358_n132787# 0.011611f
C4199 XM2/a_n100_n311027# XM3/a_n100_n104615# 0.005614f
C4200 XM1/a_n158_21658# XM2/a_n100_n134415# 7.26e-20
C4201 XM2/a_100_n155406# XM3/a_n100_49749# 0.010147f
C4202 XM1/a_n100_80437# m1_1634_n2388# 2.94e-20
C4203 XM1/a_n100_97669# XM2/a_100_n57874# 7.26e-20
C4204 XM1/a_100_60430# XM2/a_100_n94778# 4.64e-21
C4205 XM4/w_n358_n132787# XM4/a_n100_n48671# -0.004445f
C4206 XM3/a_n158_n19566# m1_1634_n2388# 6.1e-20
C4207 XM1/a_n158_150898# XM2/a_n100_n5251# 3.76e-20
C4208 XM2/a_n100_n121235# XM4/a_100_86106# 1.4e-20
C4209 XM1/a_100_n50142# XM2/a_100_n202854# 4.64e-21
C4210 XM2/a_100_n78962# XM3/a_n158_125474# 0.042475f
C4211 XM1/a_n100_15817# XM4/w_n358_n132787# 0.013586f
C4212 XM4/a_100_57098# m1_1634_n2388# 6.1e-20
C4213 XM1/a_n100_152237# XM2/a_100_n2518# 7.26e-20
C4214 XM1/a_100_56122# XM2/a_100_n97414# 4.64e-21
C4215 XM2/a_100_n303022# XM3/a_n158_n98302# 0.070126f
C4216 XM1/a_100_148026# XM4/w_n358_n132787# 0.053546f
C4217 XM1/a_n100_50281# XM2/a_n158_n105322# 0.005074f
C4218 XM1/a_n158_15914# XM2/a_n100_n139687# 7.26e-20
C4219 XM1/a_n100_n109115# XM3/a_n158_n57898# 2.43e-20
C4220 XM3/a_n100_110873# XM4/a_n100_110873# 0.009521f
C4221 XM3/a_n100_n123263# m1_1634_n2388# 0.072015f
C4222 XM2/a_n100_n218767# XM3/a_n100_n11375# 6.21e-20
C4223 XM1/a_n100_n34443# XM2/a_n158_n189674# 0.005074f
C4224 XM1/a_n158_n18550# XM2/a_n100_n171319# 7.26e-20
C4225 XM1/a_n100_n74651# m1_1634_n2388# 1.3e-19
C4226 XM4/w_n358_n132787# XM2/a_100_n76326# 0.104629f
C4227 XM3/a_n100_n43491# XM4/a_n100_n43491# 0.009521f
C4228 XM2/a_100_n194946# m1_1634_n2388# 0.017213f
C4229 XM4/w_n358_n132787# XM3/a_n100_54929# 0.009186f
C4230 XM4/a_n100_120197# m1_1634_n2388# 0.072015f
C4231 XM1/a_100_40326# XM3/a_n100_91189# 2.85e-20
C4232 XM4/w_n358_n132787# XM2/a_n158_n263482# 0.107093f
C4233 XM1/a_n158_n81734# XM2/a_n100_n234583# 7.26e-20
C4234 XM4/w_n358_n132787# XM3/a_n100_n28987# 0.009186f
C4235 XM4/a_100_n14386# m1_1634_n2388# 6.1e-20
C4236 XM1/a_n158_n166458# XM3/a_n100_n116011# 1.94e-20
C4237 XM1/a_n158_n163586# XM3/a_n100_n111867# 1.94e-20
C4238 XM2/a_100_n210762# XM3/a_n158_n5062# 0.077916f
C4239 XM1/a_n100_48845# XM2/a_100_n105322# 1.45e-19
C4240 XM4/w_n358_n132787# XM4/a_n100_n88039# -0.004445f
C4241 XM3/a_n100_71505# XM4/a_n100_71505# 0.009521f
C4242 XM2/a_100_n142226# XM3/a_n100_64253# 0.005074f
C4243 XM3/a_n158_n58934# m1_1634_n2388# 6.1e-20
C4244 XM2/a_100_n252938# XM3/a_n100_n46599# 0.005074f
C4245 XM1/a_100_84842# XM2/a_100_n71054# 4.64e-21
C4246 XM1/a_100_n140610# XM3/a_n100_n90111# 2.85e-20
C4247 XM4/a_100_17730# m1_1634_n2388# 6.1e-20
C4248 XM1/a_100_n179382# XM2/a_100_n334654# 4.64e-21
C4249 XM2/a_100_n184402# XM3/a_n100_21777# 0.010147f
C4250 XM1/a_n100_81873# XM2/a_n158_n71054# 0.005074f
C4251 XM1/a_n100_57461# XM3/a_n158_109934# 9.08e-19
C4252 XM1/a_n100_n119167# XM3/a_n158_n67222# 0.001414f
C4253 XM1/a_n100_n97627# XM3/a_n158_n46502# 2.85e-20
C4254 XM1/a_n158_n61630# XM3/a_n100_n9303# 1.46e-20
C4255 XM2/a_n100_n102783# XM4/a_100_103718# 1.05e-21
C4256 XM2/a_n158_n15698# XM1/a_100_137974# 0.116862f
C4257 XM2/a_n158_n18334# XM1/a_n100_136441# 0.005074f
C4258 XM2/a_n158_n20970# XM1/a_n100_135005# 0.001535f
C4259 XM3/a_n100_93261# m1_1634_n2388# 0.072015f
C4260 XM3/a_n100_n63175# XM4/a_n100_n63175# 0.009521f
C4261 XM1/a_100_112126# XM4/w_n358_n132787# 0.048442f
C4262 XM1/a_100_24530# XM3/a_n100_76685# 2.85e-20
C4263 XM1/a_n100_n22955# m1_1634_n2388# 8.88e-20
C4264 XM1/a_n100_41665# XM2/a_100_n113230# 7.26e-20
C4265 XM1/a_100_n111890# XM4/w_n358_n132787# 0.048442f
C4266 XM4/a_n100_80829# m1_1634_n2388# 0.072015f
C4267 XM2/a_n100_n134415# m1_1634_n2388# 0.002277f
C4268 XM1/a_n100_20125# XM3/a_n158_70566# 1.29e-20
C4269 XM1/a_100_n126250# XM2/a_n158_n279298# 0.063116f
C4270 XM4/w_n358_n132787# XM3/a_n100_n68355# 0.009186f
C4271 XM4/a_100_n53754# m1_1634_n2388# 6.1e-20
C4272 XM3/a_n100_38353# m1_1634_n2388# 0.072015f
C4273 XM2/a_n100_n289939# XM4/a_100_n85870# 1.82e-20
C4274 XM2/a_100_n326746# XM3/a_n100_n122227# 0.005074f
C4275 XM1/a_100_n127686# XM4/w_n358_n132787# 0.048442f
C4276 XM4/w_n358_n132787# XM2/a_100_n200218# 0.103341f
C4277 XM1/a_n158_56122# XM3/a_n100_106729# 1.94e-20
C4278 XM1/a_n100_50281# XM3/a_n158_102682# 2.85e-20
C4279 XM4/w_n358_n132787# XM4/a_n100_n127407# -0.004445f
C4280 XM2/a_100_n318838# m1_1634_n2388# 0.023432f
C4281 XM1/a_100_n65938# XM2/a_n100_n218767# 0.005074f
C4282 XM1/a_n100_n40187# XM2/a_100_n194946# 7.26e-20
C4283 XM3/a_n158_n98302# m1_1634_n2388# 6.1e-20
C4284 XM1/a_n100_n18647# XM2/a_100_n171222# 7.26e-20
C4285 sw_b sw_bn 0.034913f
C4286 XM1/a_n100_68949# XM3/a_n100_120197# 6.37e-19
C4287 XM4/w_n358_n132787# XM3/a_n158_79890# 0.032295f
C4288 XM2/a_n158_n126410# XM3/a_n100_77721# 7.26e-20
C4289 XM1/a_n100_17253# XM3/a_n100_68397# 2.98e-19
C4290 XM1/a_n158_n154970# XM2/a_n100_n308391# 7.26e-20
C4291 XM4/a_100_8406# m1_1634_n2388# 6.1e-20
C4292 XM1/a_n100_n90447# XM4/w_n358_n132787# 0.01363f
C4293 XM2/a_n100_n200315# XM4/a_100_6334# 2.56e-20
C4294 XM4/w_n358_n132787# XM3/a_n158_24982# 0.038676f
C4295 XM2/a_n158_n168586# XM3/a_n100_35245# 2.27e-20
C4296 XM1/a_n158_n144918# XM2/a_n158_n297750# 4.64e-21
C4297 XM1/a_n100_n70343# XM2/a_n100_n224039# 1.55e-20
C4298 XM4/w_n358_n132787# XM3/a_n158_n4026# 0.03903f
C4299 XM2/a_n100_n176591# XM4/a_100_28090# 2.56e-20
C4300 XM1/a_n158_173874# XM2/a_n100_18473# 7.26e-20
C4301 XM1/a_100_n182254# XM2/a_100_n337290# 4.64e-21
C4302 XM1/a_n100_n7159# XM3/a_n158_44666# 2.85e-20
C4303 XM2/a_100_n121138# XM3/a_n158_82998# 0.013265f
C4304 XM1/a_n158_11606# XM3/a_n100_62181# 1.94e-20
C4305 XM1/a_100_n87478# XM3/a_n158_n35106# 0.00106f
C4306 XM2/a_100_n234486# XM3/a_n100_n28987# 0.010147f
C4307 XM2/a_n158_n97414# XM3/a_n100_107765# 1.45e-19
C4308 XM3/a_n100_n82859# XM4/a_n100_n82859# 0.009521f
C4309 XM2/a_n100_n231947# XM3/a_n158_n27854# 0.004998f
C4310 XM2/a_n100_21# XM4/w_n358_n132787# 0.013902f
C4311 XM1/a_n100_28741# XM4/w_n358_n132787# 0.01363f
C4312 XM4/a_n100_41461# m1_1634_n2388# 0.072015f
C4313 XM1/a_n158_n7062# XM3/a_n100_44569# 1.94e-20
C4314 XM4/w_n358_n132787# XM3/a_n100_n107723# 0.009042f
C4315 XM4/a_100_n93122# m1_1634_n2388# 6.1e-20
C4316 XM2/a_n100_n274123# XM3/a_n100_n69391# 9.71e-19
C4317 XM1/a_n158_158078# XM2/a_n158_2754# 4.64e-21
C4318 XM1/a_n100_43101# m1_1634_n2388# 6.74e-20
C4319 XM1/a_n100_n111987# XM4/w_n358_n132787# 0.01363f
C4320 XM1/a_100_n41526# XM2/a_n100_n195043# 0.005074f
C4321 XM1/a_n158_n165022# XM3/a_n100_n112903# 1.94e-20
C4322 XM2/a_n158_n229214# XM3/a_n158_n22674# 4.64e-21
C4323 XM4/w_n358_n132787# XM2/a_n100_n139687# 0.024619f
C4324 XM2/a_n100_n258307# m1_1634_n2388# 7.61e-19
C4325 XM2/a_n158_n271390# XM3/a_n100_n64211# 1.97e-20
C4326 XM1/a_n158_179618# XM2/a_n158_26478# 4.64e-21
C4327 XM2/a_n158_n113230# XM3/a_n100_92225# 1.45e-19
C4328 XM4/w_n358_n132787# XM2/a_100_n324110# 0.10657f
C4329 XM3/a_n158_63314# m1_1634_n2388# 6.1e-20
C4330 XM4/w_n358_n132787# XM3/a_n158_n43394# 0.038462f
C4331 XM4/a_n100_n30023# m1_1634_n2388# 0.072015f
C4332 XM1/a_n100_n66035# XM2/a_100_n221306# 7.26e-20
C4333 XM2/a_n158_n155406# XM3/a_n100_49749# 1.45e-19
C4334 XM1/a_n100_n77523# m1_1634_n2388# 9.41e-20
C4335 XM1/a_100_n73118# XM2/a_n100_n229311# 2.49e-20
C4336 XM1/a_100_60430# XM2/a_n158_n94778# 0.077137f
C4337 XM1/a_n100_n134963# XM4/w_n358_n132787# 0.012803f
C4338 XM1/a_n100_n66035# XM3/a_n158_n15422# 2.85e-20
C4339 XM2/a_100_n78962# XM3/a_n100_125377# 0.005074f
C4340 XM2/a_n158_n78962# XM3/a_n158_125474# 4.64e-21
C4341 XM2/a_100_n107958# XM3/a_n158_97502# 0.077916f
C4342 XM3/a_n100_n102543# XM4/a_n100_n102543# 0.009521f
C4343 XM1/a_100_n50142# XM2/a_n158_n202854# 0.030401f
C4344 XM1/a_100_94894# XM2/a_n158_n60510# 0.058053f
C4345 XM1/a_100_155206# XM2/a_n100_21# 0.005074f
C4346 XM1/a_n100_132133# XM2/a_n158_n23606# 0.005074f
C4347 XM1/a_100_56122# XM2/a_n158_n97414# 0.110631f
C4348 XM2/a_100_n150134# XM3/a_n158_55026# 0.077916f
C4349 XM2/a_n158_n303022# XM3/a_n158_n98302# 4.64e-21
C4350 XM1/a_100_n42962# XM4/w_n358_n132787# 0.048442f
C4351 XM1/a_100_n24294# XM3/a_n100_25921# 3.44e-21
C4352 XM2/a_100_n216034# XM3/a_n100_n11375# 0.005074f
C4353 XM1/a_n158_n51578# XM3/a_n100_21# 1.94e-20
C4354 XM2/a_100_n192310# XM3/a_n158_12550# 0.077916f
C4355 XM3/a_n100_39389# XM4/a_n100_39389# 0.009521f
C4356 XM1/a_100_81970# XM2/a_n100_n71151# 0.005074f
C4357 XM4/w_n358_n132787# XM2/a_n158_n76326# 0.107093f
C4358 XM4/w_n358_n132787# XM4/a_n100_96369# -0.004445f
C4359 XM1/a_100_n144918# XM2/a_100_n300386# 4.64e-21
C4360 XM3/a_n100_n10339# m1_1634_n2388# 0.072015f
C4361 XM1/a_100_n21422# XM3/a_n100_29029# 2.85e-20
C4362 XM2/a_n100_n255671# XM3/a_n100_n51779# 0.004434f
C4363 XM1/a_n158_50378# XM2/a_n158_n102686# 4.64e-21
C4364 XM1/a_n100_11509# XM4/w_n358_n132787# 0.01363f
C4365 XM4/w_n358_n132787# XM3/a_n158_n82762# 0.038635f
C4366 XM4/a_n100_n69391# m1_1634_n2388# 0.072015f
C4367 XM4/w_n358_n132787# XM2/a_n100_n263579# 0.025738f
C4368 XM1/a_100_116434# XM2/a_n100_n39519# 0.005074f
C4369 XM3/a_n158_116150# m1_1634_n2388# 6.1e-20
C4370 XM1/a_n100_48845# XM2/a_n158_n105322# 0.010147f
C4371 XM1/a_n100_n116295# XM3/a_n158_n65150# 2.85e-20
C4372 XM1/a_n100_n107679# XM3/a_n158_n55826# 2.85e-20
C4373 XM1/a_100_41762# XM3/a_n158_93358# 0.003891f
C4374 XM2/a_n158_n142226# XM3/a_n100_64253# 7.26e-20
C4375 XM3/a_n100_n122227# XM4/a_n100_n122227# 0.009521f
C4376 XM2/a_n158_n252938# XM3/a_n100_n46599# 7.26e-20
C4377 XM1/a_n100_31613# XM3/a_n100_81865# 4.24e-19
C4378 XM1/a_100_n179382# XM2/a_n158_n334654# 0.070905f
C4379 XM2/a_100_n208126# XM3/a_n100_n2051# 0.010147f
C4380 XM1/a_n158_44634# XM2/a_n158_n107958# 4.64e-21
C4381 XM2/a_n158_n184402# XM3/a_n100_21777# 1.45e-19
C4382 XM1/a_n100_37357# XM3/a_n158_89214# 2.85e-20
C4383 XM1/a_n158_n24294# XM3/a_n100_25921# 1.8e-21
C4384 XM4/a_100_130654# m1_1634_n2388# 6.1e-20
C4385 XM1/a_n100_77565# XM3/a_n158_128582# 2.85e-20
C4386 XM2/a_100_n136954# XM3/a_n158_69530# 0.069737f
C4387 XM1/a_100_n1318# XM2/a_n158_n155406# 0.116862f
C4388 XM1/a_n158_n32910# XM3/a_n100_18669# 1.94e-20
C4389 XM1/a_100_n19986# XM3/a_n100_32137# 2.85e-20
C4390 XM4/w_n358_n132787# XM4/a_n100_57001# -0.004445f
C4391 XM3/a_n100_n49707# m1_1634_n2388# 0.072015f
C4392 XM2/a_100_n179130# XM3/a_n158_27054# 0.077916f
C4393 XM1/a_n158_n5626# XM2/a_n158_n158042# 4.64e-21
C4394 XM1/a_100_113562# XM2/a_n100_n42155# 0.005074f
C4395 XM1/a_n100_41665# XM2/a_n158_n113230# 0.005074f
C4396 XM4/w_n358_n132787# XM3/a_n100_73577# 0.009186f
C4397 XM2/a_100_n131682# m1_1634_n2388# 0.017698f
C4398 XM4/w_n358_n132787# XM3/a_n158_n122130# 0.037109f
C4399 XM4/a_n100_n108759# m1_1634_n2388# 0.072015f
C4400 XM1/a_100_n126250# XM2/a_n100_n279395# 0.005074f
C4401 XM1/a_100_176746# XM2/a_n100_23745# 0.005074f
C4402 XM2/a_n158_n326746# XM3/a_n100_n122227# 7.26e-20
C4403 XM1/a_100_n129122# XM2/a_100_n284570# 4.64e-21
C4404 XM4/w_n358_n132787# XM2/a_n158_n200218# 0.107093f
C4405 XM1/a_n100_n180915# XM3/a_n158_n128346# 8.15e-21
C4406 XM2/a_n158_n318838# m1_1634_n2388# 2.36e-21
C4407 XM1/a_100_n74554# XM3/a_n100_n22771# 2.85e-20
C4408 XM1/a_n100_n40187# XM2/a_n158_n194946# 0.005074f
C4409 XM4/w_n358_n132787# XM3/a_n100_18669# 0.009068f
C4410 XM1/a_n158_n182254# sw_b 0.003166f
C4411 XM1/a_n100_n18647# XM2/a_n158_n171222# 0.005074f
C4412 XM1/a_100_13042# XM3/a_n100_65289# 2.85e-20
C4413 XM2/a_100_n281934# XM3/a_n158_n75510# 0.075579f
C4414 XM1/a_n100_n41623# m1_1634_n2388# 9.21e-20
C4415 XM1/a_100_173874# XM2/a_n158_18570# 0.06779f
C4416 XM4/w_n358_n132787# XM3/a_n158_114078# 0.032295f
C4417 XM2/a_n100_n287303# XM4/a_100_n80690# 2.56e-20
C4418 XM4/w_n358_n132787# XM4/a_n100_n14483# -0.004445f
C4419 XM2/a_100_n324110# XM3/a_n100_n117047# 0.005074f
C4420 XM2/a_n100_n168683# XM3/a_n100_35245# 0.003206f
C4421 XM4/a_100_91286# m1_1634_n2388# 6.1e-20
C4422 XM1/a_n158_n144918# XM2/a_n100_n297847# 7.26e-20
C4423 XM1/a_n158_34582# XM2/a_n158_n121138# 4.64e-21
C4424 XM1/a_100_n182254# XM2/a_n158_n337290# 0.093884f
C4425 XM2/a_100_n73690# XM3/a_n158_131690# 0.077916f
C4426 XM2/a_100_n97414# XM3/a_n158_108898# 0.077916f
C4427 XM2/a_n158_n121138# XM3/a_n158_82998# 4.64e-21
C4428 XM1/a_100_18786# m1_1634_n2388# 0.002304f
C4429 XM2/a_n158_n234486# XM3/a_n100_n28987# 1.45e-19
C4430 XM4/w_n358_n132787# XM4/a_n100_17633# -0.004445f
C4431 XM3/a_n100_n89075# m1_1634_n2388# 0.072015f
C4432 XM4/w_n358_n132787# XM3/a_n100_21# 0.009023f
C4433 XM2/a_n100_n173955# XM4/a_100_33270# 2.56e-20
C4434 XM3/a_n100_57001# m1_1634_n2388# 0.072015f
C4435 XM1/a_100_n60194# XM2/a_100_n216034# 4.64e-21
C4436 XM1/a_100_n34346# XM4/w_n358_n132787# 0.05497f
C4437 XM1/a_n100_64641# XM3/a_n158_115114# 2.23e-20
C4438 XM1/a_100_n156406# XM3/a_n100_n104615# 2.85e-20
C4439 XM2/a_n100_n229311# XM3/a_n158_n22674# 0.005074f
C4440 XM4/w_n358_n132787# XM2/a_100_n136954# 0.103341f
C4441 XM2/a_100_n255574# m1_1634_n2388# 0.022118f
C4442 XM1/a_n100_n143579# m1_1634_n2388# 8.14e-20
C4443 XM2/a_n100_n271487# XM3/a_n100_n64211# 0.003456f
C4444 XM4/w_n358_n132787# XM4/a_n100_n53851# -0.004445f
C4445 XM3/a_n158_n24746# m1_1634_n2388# 6.1e-20
C4446 XM4/w_n358_n132787# XM3/a_n158_98538# 0.034231f
C4447 XM4/w_n358_n132787# XM2/a_n158_n324110# 0.102439f
C4448 XM1/a_n100_n133527# m1_1634_n2388# 1.3e-19
C4449 XM1/a_n100_n71779# XM2/a_100_n226578# 7.26e-20
C4450 XM3/a_n100_5201# XM4/a_n100_5201# 0.009521f
C4451 XM4/a_100_51918# m1_1634_n2388# 6.1e-20
C4452 XM1/a_n158_n183690# XM3/a_n100_n131551# 1.94e-20
C4453 XM1/a_n100_n66035# XM2/a_n158_n221306# 0.005074f
C4454 XM1/a_n158_21658# XM2/a_n158_n131682# 4.64e-21
C4455 XM4/w_n358_n132787# XM3/a_n158_43630# 0.039314f
C4456 XM1/a_100_n73118# XM2/a_100_n226578# 4.64e-21
C4457 XM1/a_100_60430# XM2/a_n100_n94875# 0.005074f
C4458 XM3/a_n100_92225# XM4/a_n100_92225# 0.009521f
C4459 XM1/a_n100_n178043# XM3/a_n158_n126274# 2.2e-20
C4460 XM2/a_n158_n78962# XM3/a_n100_125377# 7.26e-20
C4461 XM2/a_n100_n79059# XM3/a_n158_125474# 0.005074f
C4462 XM3/a_n100_n128443# m1_1634_n2388# 0.072015f
C4463 XM2/a_100_n263482# XM3/a_n158_n57898# 0.077916f
C4464 XM1/a_100_n50142# XM2/a_n100_n202951# 0.005074f
C4465 XM4/w_n358_n132787# XM4/a_n100_8309# -0.004445f
C4466 XM1/a_n100_n15775# m1_1634_n2388# 1.3e-19
C4467 XM2/a_100_n305658# XM3/a_n100_n99435# 0.009343f
C4468 XM1/a_100_56122# XM2/a_n100_n97511# 0.002863f
C4469 XM1/a_n100_n170863# XM3/a_n158_n120058# 2.85e-20
C4470 XM1/a_n158_n152098# XM2/a_n158_n305658# 4.64e-21
C4471 XM1/a_100_168130# XM2/a_n158_13298# 0.113746f
C4472 XM2/a_n100_n303119# XM3/a_n158_n98302# 0.004269f
C4473 XM1/a_n100_50281# XM2/a_100_n102686# 7.26e-20
C4474 XM1/a_n158_15914# XM2/a_n158_n136954# 4.64e-21
C4475 XM1/a_100_n173638# XM3/a_n100_n122227# 5.56e-19
C4476 XM1/a_100_n90350# XM4/w_n358_n132787# 0.048442f
C4477 XM4/a_n100_115017# m1_1634_n2388# 0.072015f
C4478 XM4/w_n358_n132787# XM3/a_n100_n34167# 0.009186f
C4479 XM4/a_100_n19566# m1_1634_n2388# 6.1e-20
C4480 XM1/a_100_n67374# XM2/a_n158_n221306# 0.116862f
C4481 XM2/a_n158_n216034# XM3/a_n100_n11375# 7.26e-20
C4482 XM1/a_n100_n53111# XM3/a_n158_n918# 2.85e-20
C4483 XM1/a_n100_n34443# XM2/a_100_n187038# 7.26e-20
C4484 XM4/w_n358_n132787# XM2/a_n100_n76423# 0.025015f
C4485 XM1/a_100_n144918# XM2/a_n158_n300386# 0.051822f
C4486 XM4/w_n358_n132787# XM4/a_n100_n93219# -0.004445f
C4487 XM1/a_n100_n132091# XM2/a_100_n287206# 7.26e-20
C4488 XM3/a_n158_n64114# m1_1634_n2388# 6.1e-20
C4489 XM1/a_100_n63066# XM2/a_100_n218670# 4.64e-21
C4490 XM2/a_n100_n195043# m1_1634_n2388# 0.002198f
C4491 XM1/a_100_166694# XM2/a_100_13298# 4.64e-21
C4492 XM1/a_n100_n35879# XM3/a_n100_16597# 9.89e-19
C4493 XM1/a_n158_50378# XM2/a_n100_n102783# 7.26e-20
C4494 XM4/a_100_12550# m1_1634_n2388# 6.1e-20
C4495 XM4/w_n358_n132787# XM2/a_100_n260846# 0.106421f
C4496 XM2/a_100_n213398# XM3/a_n100_n6195# 1.17e-21
C4497 XM3/a_n158_81962# m1_1634_n2388# 6.1e-20
C4498 XM3/a_n100_116053# m1_1634_n2388# 0.072015f
C4499 XM1/a_n158_46070# XM3/a_n100_96369# 1.86e-20
C4500 XM1/a_n100_40229# XM3/a_n158_92322# 2.85e-20
C4501 XM1/a_100_n103274# XM4/w_n358_n132787# 0.052497f
C4502 XM1/a_n100_n162247# XM3/a_n158_n109698# 1.4e-20
C4503 XM1/a_n100_n93319# XM3/a_n158_n42358# 2.85e-20
C4504 XM1/a_100_n90350# XM3/a_n100_n38311# 2.85e-20
C4505 XM1/a_100_n63066# XM3/a_n100_n11375# 0.001635f
C4506 XM2/a_n100_n253035# XM3/a_n100_n46599# 0.003389f
C4507 XM3/a_n158_27054# m1_1634_n2388# 6.1e-20
C4508 XM1/a_100_n179382# XM2/a_n100_n334751# 0.005074f
C4509 XM1/a_n100_n55983# XM3/a_n158_n4026# 0.001287f
C4510 XM2/a_n158_n208126# XM3/a_n100_n2051# 1.45e-19
C4511 XM1/a_n158_44634# XM2/a_n100_n108055# 7.26e-20
C4512 XM1/a_n100_117773# XM4/w_n358_n132787# 0.012279f
C4513 XM1/a_n100_7201# XM4/w_n358_n132787# 0.011991f
C4514 XM2/a_n158_23842# XM1/a_100_178182# 0.116862f
C4515 XM4/a_n100_75649# m1_1634_n2388# 0.072015f
C4516 XM2/a_n158_n136954# XM3/a_n158_69530# 4.64e-21
C4517 XM4/w_n358_n132787# XM3/a_n100_n73535# 0.009186f
C4518 XM4/a_100_n58934# m1_1634_n2388# 6.1e-20
C4519 XM1/a_100_n5626# XM2/a_100_n160678# 4.64e-21
C4520 XM2/a_n158_26478# XM1/a_n100_182393# 0.004836f
C4521 XM2/a_n100_26381# XM1/a_n158_182490# 6.36e-20
C4522 XM2/a_100_29114# XM1/a_100_182490# 4.64e-21
C4523 XM1/a_100_34582# XM3/a_n100_86009# 2.97e-19
C4524 XM1/a_n100_24433# m1_1634_n2388# 5.93e-19
C4525 XM1/a_n100_n178043# XM4/w_n358_n132787# 0.013551f
C4526 XM2/a_100_n245030# XM3/a_n158_n40286# 0.072463f
C4527 XM1/a_100_n84606# XM3/a_n158_n33034# 0.00544f
C4528 XM1/a_n158_n5626# XM2/a_n100_n158139# 7.26e-20
C4529 XM3/a_n158_n103482# m1_1634_n2388# 6.1e-20
C4530 XM2/a_100_n287206# XM3/a_n100_n81823# 0.010147f
C4531 XM3/a_n100_8309# m1_1634_n2388# 0.072015f
C4532 XM2/a_n158_n131682# m1_1634_n2388# 2.36e-21
C4533 XM1/a_100_n129122# XM2/a_n158_n284570# 0.053769f
C4534 XM4/w_n358_n132787# XM2/a_n100_n200315# 0.025738f
C4535 XM1/a_n100_n12903# XM4/w_n358_n132787# 0.0135f
C4536 XM2/a_n100_n318935# m1_1634_n2388# 9.56e-19
C4537 XM1/a_n158_n90350# XM3/a_n100_n38311# 1.94e-20
C4538 XM1/a_n100_n40187# XM2/a_n100_n195043# 0.00131f
C4539 XM1/a_n158_n8498# XM3/a_n158_43630# 1.14e-21
C4540 XM1/a_100_27402# XM3/a_n100_77721# 2.85e-20
C4541 XM1/a_n100_21561# XM3/a_n158_73674# 2.85e-20
C4542 XM4/w_n358_n132787# XM3/a_n158_n9206# 0.038462f
C4543 XM1/a_n100_110593# XM2/a_n158_n42058# 0.005074f
C4544 XM1/a_n100_68949# XM3/a_n158_121330# 2.85e-20
C4545 XM2/a_n158_n281934# XM3/a_n158_n75510# 4.64e-21
C4546 XM1/a_n100_n63163# XM3/a_n158_n11278# 2.85e-20
C4547 XM1/a_n100_n43059# m1_1634_n2388# 8.14e-20
C4548 XM1/a_n100_n22955# XM2/a_100_n176494# 9.95e-20
C4549 XM4/w_n358_n132787# XM3/a_n100_113981# 0.009186f
C4550 XM1/a_n100_18689# XM3/a_n158_69530# 2.85e-20
C4551 XM2/a_n158_n324110# XM3/a_n100_n117047# 7.26e-20
C4552 XM1/a_n100_n153631# m1_1634_n2388# 9.15e-20
C4553 XM1/a_n100_27305# XM4/w_n358_n132787# 0.01335f
C4554 XM4/a_n100_36281# m1_1634_n2388# 0.072015f
C4555 XM4/w_n358_n132787# XM3/a_n100_n112903# 0.009186f
C4556 XM4/a_100_n98302# m1_1634_n2388# 6.1e-20
C4557 XM1/a_n158_34582# XM2/a_n100_n121235# 7.26e-20
C4558 XM2/a_n100_n121235# XM3/a_n158_82998# 0.005074f
C4559 XM1/a_100_n182254# XM2/a_n100_n337387# 0.005074f
C4560 XM2/a_100_n73690# XM3/a_n100_131593# 0.010147f
C4561 XM2/a_100_n97414# XM3/a_n100_108801# 0.009971f
C4562 XM1/a_n100_n179479# XM3/a_n158_n128346# 2.85e-20
C4563 XM1/a_100_n126250# XM3/a_n158_n75510# 9.08e-19
C4564 XM1/a_n158_n98966# XM2/a_n158_n252938# 9.28e-21
C4565 XM4/w_n358_n132787# XM4/a_n100_130557# -0.004445f
C4566 XM1/a_100_n31474# XM3/a_n100_19705# 5.17e-20
C4567 XM4/w_n358_n132787# XM3/a_n100_92225# 0.009186f
C4568 XM1/a_100_97766# XM2/a_100_n55238# 4.64e-21
C4569 XM1/a_n158_n179382# XM3/a_n100_n128443# 1.84e-20
C4570 XM1/a_100_n121942# XM4/w_n358_n132787# 0.048442f
C4571 XM1/a_100_n60194# XM2/a_n158_n216034# 0.015602f
C4572 XM1/a_n100_64641# XM3/a_n100_115017# 3.12e-19
C4573 XM1/a_n158_n156406# XM3/a_n100_n105651# 1.94e-20
C4574 XM4/w_n358_n132787# XM3/a_n158_n48574# 0.038462f
C4575 XM4/a_n100_n35203# m1_1634_n2388# 0.072015f
C4576 XM4/w_n358_n132787# XM2/a_n158_n136954# 0.107093f
C4577 XM2/a_n158_n255574# m1_1634_n2388# 2.36e-21
C4578 XM2/a_n100_n231947# XM4/a_100_n27854# 2.45e-20
C4579 XM4/w_n358_n132787# XM3/a_n100_37317# 0.009055f
C4580 XM3/a_n100_60109# XM4/a_n100_60109# 0.009521f
C4581 XM2/a_100_n268754# XM3/a_n100_n64211# 0.005074f
C4582 XM4/w_n358_n132787# XM2/a_n100_n324207# 0.025375f
C4583 XM1/a_100_21658# XM2/a_100_n134318# 4.64e-21
C4584 XM1/a_n100_n91883# XM2/a_100_n247666# 7.26e-20
C4585 XM1/a_n100_n80395# m1_1634_n2388# 8.14e-20
C4586 XM1/a_n100_n71779# XM2/a_n158_n226578# 0.005074f
C4587 XM1/a_n158_21658# XM2/a_n100_n131779# 7.26e-20
C4588 XM1/a_100_n162150# XM2/a_n158_n316202# 0.116862f
C4589 XM1/a_100_67610# XM4/w_n358_n132787# 0.048442f
C4590 XM1/a_100_n78862# XM4/w_n358_n132787# 0.054613f
C4591 XM1/a_100_n73118# XM2/a_n158_n226578# 0.103231f
C4592 XM1/a_100_60430# XM2/a_100_n92142# 4.64e-21
C4593 XM1/a_100_n68810# XM4/w_n358_n132787# 0.054848f
C4594 XM2/a_100_n78962# XM3/a_n158_126510# 0.077916f
C4595 XM2/a_n100_n118599# XM4/a_100_86106# 2.56e-20
C4596 XM2/a_n158_n28878# XM4/w_n358_n132787# 0.107093f
C4597 XM4/w_n358_n132787# XM4/a_n100_91189# -0.004445f
C4598 XM1/a_n100_n176607# XM2/a_100_n332018# 7.26e-20
C4599 XM2/a_n158_n305658# XM3/a_n100_n99435# 1.36e-19
C4600 XM1/a_n158_n152098# XM2/a_n100_n305755# 3.29e-20
C4601 XM3/a_n100_n15519# m1_1634_n2388# 0.072015f
C4602 XM1/a_100_n45834# XM3/a_n100_5201# 2.85e-20
C4603 XM1/a_100_120742# XM4/w_n358_n132787# 0.049913f
C4604 XM1/a_n100_50281# XM2/a_n158_n102686# 0.005074f
C4605 XM1/a_n100_18689# XM4/w_n358_n132787# 0.01363f
C4606 XM1/a_n158_15914# XM2/a_n100_n137051# 7.26e-20
C4607 XM1/a_n158_n172202# XM3/a_n100_n120155# 1.94e-20
C4608 XM4/w_n358_n132787# XM3/a_n158_n87942# 0.038462f
C4609 XM4/a_n100_n74571# m1_1634_n2388# 0.072015f
C4610 XM2/a_n100_n216131# XM3/a_n100_n11375# 0.002506f
C4611 XM1/a_n100_n34443# XM2/a_n158_n187038# 0.005074f
C4612 XM3/a_n100_75649# m1_1634_n2388# 0.072015f
C4613 XM1/a_100_n144918# XM2/a_n100_n300483# 0.005074f
C4614 XM1/a_n100_n132091# XM2/a_n158_n287206# 0.005074f
C4615 XM1/a_n158_n91786# XM3/a_n100_n40383# 3.61e-20
C4616 XM1/a_100_n71682# XM3/a_n158_n19566# 0.001891f
C4617 XM1/a_100_n63066# XM2/a_n158_n218670# 0.03858f
C4618 XM2/a_100_n192310# m1_1634_n2388# 0.019664f
C4619 XM2/a_n100_n300483# XM3/a_n158_n93122# 0.002238f
C4620 XM3/a_n100_20741# m1_1634_n2388# 0.072015f
C4621 XM1/a_100_126486# XM2/a_n158_n26242# 0.031959f
C4622 XM4/w_n358_n132787# XM2/a_n158_n260846# 0.103717f
C4623 XM1/a_n158_122178# XM2/a_n158_n31514# 9.28e-21
C4624 XM1/a_n158_81970# XM2/a_n158_n73690# 4.64e-21
C4625 XM1/a_100_n142046# XM3/a_n100_n90111# 2.85e-20
C4626 XM2/a_n158_2754# XM4/w_n358_n132787# 0.107093f
C4627 XM4/w_n358_n132787# XM1/a_n100_139313# 0.012279f
C4628 XM1/a_100_n24294# XM4/w_n358_n132787# 0.04959f
C4629 XM1/a_n100_n99063# XM3/a_n158_n46502# 1.05e-20
C4630 XM4/a_100_125474# m1_1634_n2388# 6.1e-20
C4631 XM2/a_100_n139590# XM3/a_n100_64253# 0.002589f
C4632 XM4/w_n358_n132787# XM3/a_n158_62278# 0.038479f
C4633 XM1/a_100_n179382# XM2/a_100_n332018# 4.64e-21
C4634 XM1/a_100_n97530# m1_1634_n2388# 0.001092f
C4635 XM1/a_n100_n68907# XM3/a_n100_n18627# 6.81e-19
C4636 XM4/w_n358_n132787# XM4/a_n100_51821# -0.004445f
C4637 XM3/a_n100_n54887# m1_1634_n2388# 0.072015f
C4638 XM2/a_n158_18570# XM4/w_n358_n132787# 0.107093f
C4639 XM2/a_100_n334654# XM3/a_n158_n128346# 0.077916f
C4640 XM1/a_n100_41665# XM4/w_n358_n132787# 0.012605f
C4641 XM2/a_n100_n137051# XM3/a_n158_69530# 0.004619f
C4642 XM1/a_100_148026# XM2/a_n158_n7790# 0.017938f
C4643 XM4/w_n358_n132787# XM3/a_n158_n127310# 0.034105f
C4644 XM4/a_n100_n113939# m1_1634_n2388# 0.072015f
C4645 XM3/a_n100_n9303# XM4/a_n100_n9303# 0.009521f
C4646 XM1/a_100_n5626# XM2/a_n158_n160678# 0.092326f
C4647 XM1/a_100_n153534# XM4/w_n358_n132787# 0.048442f
C4648 XM2/a_n158_n245030# XM3/a_n158_n40286# 4.64e-21
C4649 sw_b XM2/a_n158_n337290# 0.003001f
C4650 XM2/a_n100_n10523# XM1/a_n158_145154# 7.26e-20
C4651 XM2/a_n158_n10426# XM1/a_100_145154# 0.040917f
C4652 XM2/a_100_n10426# XM1/a_n100_143621# 1.45e-19
C4653 XM1/a_n158_28838# XM3/a_n100_80829# 7.81e-21
C4654 XM2/a_n158_n287206# XM3/a_n100_n81823# 1.45e-19
C4655 XM1/a_100_n78862# XM2/a_100_n234486# 4.64e-21
C4656 XM1/a_n158_152334# XM2/a_n158_n2518# 4.64e-21
C4657 XM1/a_n100_41665# XM2/a_100_n110594# 4.26e-20
C4658 XM2/a_n100_n131779# m1_1634_n2388# 0.001257f
C4659 XM4/w_n358_n132787# XM4/a_n100_n19663# -0.004445f
C4660 XM1/a_100_n129122# XM2/a_n100_n284667# 0.005074f
C4661 XM4/w_n358_n132787# XM2/a_100_n197582# 0.105777f
C4662 XM1/a_100_118# XM4/w_n358_n132787# 0.054961f
C4663 XM1/a_100_155206# XM2/a_n158_2754# 0.005086f
C4664 XM2/a_n100_n15795# XM1/a_n100_137877# 6.96e-19
C4665 XM1/a_n158_110690# XM2/a_n158_n44694# 4.64e-21
C4666 XM1/a_n158_56122# XM3/a_n100_107765# 1.94e-20
C4667 XM1/a_n158_n183690# iout 0.010558f
C4668 XM2/a_100_n316202# m1_1634_n2388# 0.017213f
C4669 XM4/a_100_86106# m1_1634_n2388# 6.1e-20
C4670 XM1/a_100_n53014# XM3/a_n100_n2051# 2.85e-20
C4671 XM2/a_100_n126410# XM3/a_n100_78757# 0.010147f
C4672 XM1/a_n100_n129219# XM3/a_n158_n78618# 2.85e-20
C4673 XM2/a_n100_n282031# XM3/a_n158_n75510# 4.89e-19
C4674 XM1/a_n158_n84606# XM3/a_n100_n34167# 1.94e-20
C4675 XM4/w_n358_n132787# XM4/a_n100_12453# -0.004445f
C4676 XM1/a_n100_n22955# XM2/a_n158_n176494# 0.005805f
C4677 XM3/a_n158_45702# m1_1634_n2388# 6.1e-20
C4678 XM1/a_100_110690# XM2/a_n100_n44791# 0.005074f
C4679 XM3/a_n100_n94255# m1_1634_n2388# 0.072015f
C4680 XM1/a_n158_n119070# XM3/a_n100_n68355# 1.94e-20
C4681 XM1/a_100_n41526# XM3/a_n158_9442# 0.003891f
C4682 XM2/a_n100_n197679# XM4/a_100_6334# 3.43e-21
C4683 XM2/a_100_n168586# XM3/a_n100_36281# 0.010147f
C4684 XM1/a_100_150898# XM2/a_n100_n5251# 0.003292f
C4685 XM1/a_100_n182254# XM2/a_100_n334654# 4.64e-21
C4686 XM3/a_n100_n28987# XM4/a_n100_n28987# 0.009521f
C4687 XM1/a_n158_176746# XM2/a_n100_23745# 7.26e-20
C4688 XM2/a_n158_n97414# XM3/a_n100_108801# 1.38e-19
C4689 XM3/a_n100_27993# XM4/a_n100_27993# 0.009521f
C4690 XM1/a_100_n1318# XM3/a_n100_50785# 2.85e-20
C4691 XM1/a_100_n14242# XM4/w_n358_n132787# 0.048442f
C4692 XM2/a_100_n316202# XM3/a_n158_n110734# 0.077916f
C4693 XM4/w_n358_n132787# XM4/a_n100_n59031# -0.004445f
C4694 XM3/a_n158_n29926# m1_1634_n2388# 6.1e-20
C4695 XM1/a_100_n77426# XM2/a_n158_n231850# 0.116862f
C4696 XM1/a_n158_n157842# XM3/a_n100_n106687# 2.99e-20
C4697 XM1/a_100_n60194# XM2/a_n100_n216131# 0.005074f
C4698 XM4/a_100_46738# m1_1634_n2388# 6.1e-20
C4699 XM4/w_n358_n132787# XM2/a_n100_n137051# 0.025473f
C4700 XM1/a_100_160950# XM2/a_n100_5293# 0.005074f
C4701 XM1/a_n158_96330# XM2/a_n158_n57874# 9.28e-21
C4702 XM2/a_n100_n255671# m1_1634_n2388# 0.001922f
C4703 XM2/a_n158_n268754# XM3/a_n100_n64211# 7.26e-20
C4704 XM1/a_100_n101838# XM4/w_n358_n132787# 0.048442f
C4705 XM1/a_n100_91925# XM2/a_n158_n63146# 0.005074f
C4706 XM2/a_100_n113230# XM3/a_n100_93261# 0.005074f
C4707 XM1/a_100_21658# XM2/a_n158_n134318# 0.00236f
C4708 XM4/w_n358_n132787# XM2/a_100_n321474# 0.103341f
C4709 XM1/a_n100_n91883# XM2/a_n158_n247666# 0.005074f
C4710 XM1/a_n100_n71779# XM2/a_n100_n226675# 1.55e-20
C4711 XM2/a_n100_n44791# XM4/w_n358_n132787# 0.012279f
C4712 XM2/a_100_n223942# XM3/a_n158_n17494# 0.073242f
C4713 XM1/a_n100_n66035# XM2/a_100_n218670# 7.26e-20
C4714 XM3/a_n100_n48671# XM4/a_n100_n48671# 0.009521f
C4715 XM2/a_n100_n229311# XM4/a_100_n22674# 2.56e-20
C4716 XM2/a_100_n155406# XM3/a_n100_50785# 0.010147f
C4717 XM2/a_100_n266118# XM3/a_n100_n59031# 0.005074f
C4718 XM1/a_100_n73118# XM2/a_n100_n226675# 0.005074f
C4719 XM1/a_n100_97669# XM2/a_100_n55238# 7.26e-20
C4720 XM1/a_100_60430# XM2/a_n158_n92142# 0.01677f
C4721 XM4/a_n100_n131551# XM3/a_n100_n131551# 0.009521f
C4722 XM1/a_n158_150898# XM2/a_n100_n2615# 7.26e-20
C4723 XM2/a_100_n78962# XM3/a_n100_126413# 0.010147f
C4724 XM4/a_n100_109837# m1_1634_n2388# 0.072015f
C4725 XM4/w_n358_n132787# XM3/a_n100_n39347# 0.009001f
C4726 XM4/a_100_n24746# m1_1634_n2388# 6.1e-20
C4727 XM1/a_n100_n176607# XM2/a_n158_n332018# 0.005074f
C4728 XM2/a_n100_n305755# XM3/a_n100_n99435# 4.1e-19
C4729 XM1/a_100_n100402# XM3/a_n158_n48574# 0.00544f
C4730 XM4/w_n358_n132787# XM4/a_n100_n98399# -0.004445f
C4731 XM3/a_n158_n69294# m1_1634_n2388# 6.1e-20
C4732 XM2/a_n100_n115963# XM4/a_100_91286# 2.56e-20
C4733 XM1/a_n158_87714# XM2/a_n158_n65782# 4.64e-21
C4734 XM1/a_100_n144918# XM2/a_100_n297750# 4.64e-21
C4735 XM4/w_n358_n132787# XM1/a_100_145154# 0.053546f
C4736 XM1/a_n100_n103371# XM3/a_n100_n51779# 9.88e-19
C4737 XM1/a_100_n63066# XM2/a_n100_n218767# 0.005074f
C4738 XM4/w_n358_n132787# XM3/a_n100_55965# 0.008991f
C4739 XM2/a_100_n297750# XM3/a_n158_n93122# 0.061169f
C4740 XM2/a_n100_n303119# XM4/a_100_n98302# 2.11e-20
C4741 XM1/a_100_40326# XM3/a_n100_92225# 2.85e-20
C4742 XM4/w_n358_n132787# XM2/a_n100_n260943# 0.025089f
C4743 XM1/a_n100_n64599# m1_1634_n2388# 9.68e-20
C4744 XM2/a_n100_n213495# XM3/a_n100_n6195# 0.005189f
C4745 XM3/a_n100_n68355# XM4/a_n100_n68355# 0.009521f
C4746 XM4/w_n358_n132787# XM3/a_n158_1154# 0.038462f
C4747 XM1/a_n100_120645# XM4/w_n358_n132787# 0.012195f
C4748 XM3/a_n158_117186# m1_1634_n2388# 6.1e-20
C4749 XM2/a_n158_n139590# XM3/a_n100_64253# 3.17e-20
C4750 XM1/a_100_37454# XM3/a_n100_88081# 2.85e-20
C4751 XM4/a_n100_70469# m1_1634_n2388# 0.072015f
C4752 XM4/w_n358_n132787# XM3/a_n100_n78715# 0.009186f
C4753 XM4/a_100_n64114# m1_1634_n2388# 6.1e-20
C4754 XM1/a_100_84842# XM2/a_100_n68418# 4.64e-21
C4755 XM1/a_n100_n155067# XM3/a_n100_n102543# 9.11e-19
C4756 XM1/a_100_n7062# XM2/a_n158_n160678# 0.116862f
C4757 XM3/a_n100_118125# XM4/a_n100_118125# 0.009521f
C4758 XM1/a_100_28838# m1_1634_n2388# 0.002487f
C4759 XM1/a_100_n179382# XM2/a_n158_n332018# 0.023001f
C4760 XM1/a_n100_n60291# XM3/a_n158_n9206# 2.85e-20
C4761 XM3/a_n158_n108662# m1_1634_n2388# 6.1e-20
C4762 XM1/a_n158_33146# XM3/a_n100_83937# 1.94e-20
C4763 XM1/a_n100_77565# XM3/a_n158_129618# 2.85e-20
C4764 XM2/a_100_n247666# XM3/a_n100_n41419# 0.007234f
C4765 XM1/a_100_n5626# XM2/a_n100_n160775# 0.005074f
C4766 XM1/a_100_28838# XM3/a_n100_79793# 2.85e-20
C4767 XM2/a_n100_n245127# XM3/a_n158_n40286# 0.00216f
C4768 XM2/a_n100_n18431# XM1/a_100_136538# 0.003566f
C4769 XM2/a_n158_n18334# XM1/a_n100_135005# 0.005074f
C4770 XM1/a_100_117870# XM2/a_n158_n36786# 0.116862f
C4771 XM3/a_n100_94297# m1_1634_n2388# 0.072015f
C4772 XM1/a_n100_n156503# XM2/a_100_n310930# 1.45e-19
C4773 XM1/a_n100_n124911# XM3/a_n100_n74571# 7.8e-19
C4774 XM1/a_100_n78862# XM2/a_n158_n234486# 0.036633f
C4775 XM4/w_n358_n132787# XM3/a_n158_n14386# 0.038462f
C4776 XM1/a_n100_n43059# XM3/a_n158_7370# 9.33e-21
C4777 XM1/a_n158_113562# XM2/a_n158_n42058# 4.64e-21
C4778 XM1/a_n100_41665# XM2/a_n158_n110594# 0.003994f
C4779 XM2/a_100_n129046# m1_1634_n2388# 0.017213f
C4780 XM3/a_n100_39389# m1_1634_n2388# 0.072014f
C4781 XM4/w_n358_n132787# XM1/a_n100_130697# 0.012279f
C4782 XM1/a_n158_60430# XM3/a_n100_110873# 1.94e-20
C4783 XM1/a_100_56122# XM3/a_n158_106826# 0.001549f
C4784 XM3/a_n100_n88039# XM4/a_n100_n88039# 0.009521f
C4785 XM4/w_n358_n132787# XM2/a_n158_n197582# 0.106008f
C4786 XM1/a_100_80534# XM3/a_n100_131593# 2.85e-20
C4787 XM1/a_100_n129122# XM2/a_100_n281934# 4.64e-21
C4788 XM1/a_n100_34485# XM4/w_n358_n132787# 0.013522f
C4789 XM4/a_n100_31101# m1_1634_n2388# 0.072015f
C4790 XM4/w_n358_n132787# XM3/a_n100_n118083# 0.009186f
C4791 XM4/a_100_n103482# m1_1634_n2388# 6.1e-20
C4792 XM1/a_n158_160950# XM2/a_n100_5293# 7.26e-20
C4793 XM3/a_n100_80829# XM4/a_n100_80829# 0.009521f
C4794 XM2/a_n158_n126410# XM3/a_n100_78757# 1.45e-19
C4795 XM1/a_n100_51717# m1_1634_n2388# 1.3e-19
C4796 XM4/w_n358_n132787# XM3/a_n158_80926# 0.034422f
C4797 XM1/a_n100_12945# XM3/a_n158_65386# 2.85e-20
C4798 XM1/a_n100_4329# XM3/a_n100_55965# 7.93e-19
C4799 XM1/a_n100_n22955# XM2/a_n100_n176591# 0.003193f
C4800 XM4/w_n358_n132787# XM3/a_n158_115114# 0.037075f
C4801 XM1/a_n100_n176607# XM3/a_n100_n126371# 2.18e-19
C4802 XM1/a_100_n109018# XM3/a_n100_n57995# 2.85e-20
C4803 XM2/a_100_n321474# XM3/a_n100_n117047# 0.005074f
C4804 XM4/w_n358_n132787# XM3/a_n158_26018# 0.032295f
C4805 XM2/a_n158_n168586# XM3/a_n100_36281# 1.45e-19
C4806 XM1/a_n158_173874# XM2/a_n100_21109# 7.26e-20
C4807 XM4/w_n358_n132787# XM4/a_n100_125377# -0.004445f
C4808 XM1/a_n158_34582# XM2/a_n158_n118502# 4.64e-21
C4809 XM1/a_n100_104849# XM2/a_100_n49966# 7.26e-20
C4810 XM2/a_100_n121138# XM3/a_n158_84034# 0.077916f
C4811 XM1/a_100_n182254# XM2/a_n158_n334654# 2.3e-20
C4812 XM1/a_n158_n44398# XM3/a_n100_7273# 1.94e-20
C4813 XM2/a_100_n23606# XM1/a_100_132230# 4.64e-21
C4814 XM1/a_n100_106285# XM4/w_n358_n132787# 0.012279f
C4815 XM2/a_n100_n97511# XM3/a_n100_108801# 1.4e-19
C4816 XM1/a_n158_11606# XM3/a_n100_63217# 1.94e-20
C4817 XM1/a_100_n2754# XM3/a_n100_47677# 2.85e-20
C4818 XM4/w_n358_n132787# XM3/a_n158_n53754# 0.039197f
C4819 XM4/a_n100_n40383# m1_1634_n2388# 0.072015f
C4820 XM2/a_n100_n171319# XM4/a_100_33270# 2.56e-20
C4821 XM2/a_100_n163314# XM3/a_n158_41558# 0.077916f
C4822 XM1/a_n100_14381# m1_1634_n2388# 1.3e-19
C4823 XM3/a_n100_n107723# XM4/a_n100_n107723# 0.009521f
C4824 XM1/a_n158_79098# XM2/a_n158_n76326# 4.64e-21
C4825 XM3/a_n100_101549# XM4/a_n100_101549# 0.009521f
C4826 XM2/a_100_n229214# XM3/a_n100_n23807# 0.010147f
C4827 XM1/a_100_103510# XM2/a_n100_n50063# 0.005074f
C4828 XM1/a_100_n154970# XM3/a_n100_n103579# 5.78e-19
C4829 XM1/a_100_n60194# XM2/a_100_n213398# 4.64e-21
C4830 XM4/w_n358_n132787# XM2/a_100_n134318# 0.104135f
C4831 XM2/a_n100_n226675# XM3/a_n158_n22674# 2.49e-20
C4832 XM2/a_n100_n276759# XM4/a_n100_n70427# 2.71e-20
C4833 XM2/a_100_n252938# m1_1634_n2388# 0.017213f
C4834 XM1/a_n158_n41526# XM3/a_n100_9345# 1.94e-20
C4835 XM1/a_100_n93222# XM4/w_n358_n132787# 0.048442f
C4836 XM2/a_n158_n113230# XM3/a_n100_93261# 7.26e-20
C4837 XM1/a_100_21658# XM2/a_n100_n134415# 0.005074f
C4838 XM4/w_n358_n132787# XM2/a_n158_n321474# 0.101988f
C4839 XM3/a_n158_64350# m1_1634_n2388# 6.1e-20
C4840 XM4/w_n358_n132787# XM4/a_n100_86009# -0.004445f
C4841 XM2/a_n158_n223942# XM3/a_n158_n17494# 4.64e-21
C4842 XM1/a_n100_n66035# XM2/a_n158_n218670# 0.005074f
C4843 XM2/a_n158_n155406# XM3/a_n100_50785# 1.45e-19
C4844 XM1/a_n100_58897# XM2/a_100_n94778# 1.45e-19
C4845 XM1/a_100_n156406# XM2/a_n158_n310930# 0.116862f
C4846 XM3/a_n100_n20699# m1_1634_n2388# 0.072015f
C4847 XM2/a_n158_n266118# XM3/a_n100_n59031# 7.26e-20
C4848 XM3/a_n158_9442# m1_1634_n2388# 6.1e-20
C4849 XM1/a_100_60430# XM2/a_n100_n92239# 0.005074f
C4850 XM2/a_100_n107958# XM3/a_n158_98538# 0.068569f
C4851 XM1/a_100_20222# XM4/w_n358_n132787# 0.048442f
C4852 XM1/a_100_n144918# XM4/w_n358_n132787# 0.054703f
C4853 XM4/a_n100_1057# m1_1634_n2388# 0.072015f
C4854 XM2/a_n158_n78962# XM3/a_n100_126413# 1.45e-19
C4855 XM4/w_n358_n132787# XM3/a_n158_n93122# 0.037006f
C4856 XM4/a_n100_n79751# m1_1634_n2388# 0.072015f
C4857 XM1/a_100_94894# XM2/a_n158_n57874# 0.035854f
C4858 XM1/a_n100_n113423# XM4/w_n358_n132787# 0.013538f
C4859 XM1/a_n100_132133# XM2/a_n158_n20970# 0.005074f
C4860 XM1/a_n158_90586# XM2/a_n158_n63146# 9.28e-21
C4861 XM2/a_100_n150134# XM3/a_n158_56062# 0.077916f
C4862 XM3/a_n100_n127407# XM4/a_n100_n127407# 0.009521f
C4863 XM1/a_n100_n61727# XM3/a_n158_n9206# 2.23e-20
C4864 XM1/a_100_n24294# XM3/a_n100_26957# 5.71e-20
C4865 XM1/a_n100_127825# XM2/a_n158_n26242# 0.010147f
C4866 XM1/a_n158_n110454# XM2/a_n158_n266118# 4.64e-21
C4867 XM2/a_100_n192310# XM3/a_n158_13586# 0.077916f
C4868 XM1/a_100_92022# XM4/w_n358_n132787# 0.053546f
C4869 XM1/a_100_n144918# XM2/a_n158_n297750# 0.042085f
C4870 XM1/a_100_n182254# XM3/a_n158_n130418# 0.00544f
C4871 XM1/a_n100_n132091# XM2/a_100_n284570# 7.26e-20
C4872 XM1/a_n100_n93319# XM4/w_n358_n132787# 0.01363f
C4873 XM1/a_100_n63066# XM2/a_100_n216034# 4.64e-21
C4874 XM2/a_n100_n192407# m1_1634_n2388# 0.003216f
C4875 XM1/a_100_n21422# XM3/a_n100_30065# 3.4e-20
C4876 XM4/a_100_120294# m1_1634_n2388# 6.1e-20
C4877 XM2/a_n158_n297750# XM3/a_n158_n93122# 4.64e-21
C4878 XM4/w_n358_n132787# XM4/a_n100_46641# -0.004445f
C4879 XM4/w_n358_n132787# XM2/a_100_n258210# 0.103342f
C4880 XM1/a_n100_n73215# m1_1634_n2388# 1.19e-20
C4881 XM2/a_100_n210762# XM3/a_n100_n6195# 0.005074f
C4882 XM1/a_100_116434# XM2/a_n100_n36883# 0.005074f
C4883 XM3/a_n100_n60067# m1_1634_n2388# 0.072015f
C4884 XM3/a_n100_117089# m1_1634_n2388# 0.072015f
C4885 XM1/a_n158_36018# XM3/a_n100_87045# 1.94e-20
C4886 XM2/a_n100_n139687# XM3/a_n100_64253# 0.002458f
C4887 XM4/w_n358_n132787# XM3/a_n158_n132490# 0.032295f
C4888 XM4/a_n100_n119119# m1_1634_n2388# 0.072015f
C4889 XM2/a_100_n295114# XM3/a_n158_n87942# 0.002749f
C4890 XM2/a_n100_n300483# XM4/a_100_n93122# 8.7e-21
C4891 XM1/a_n100_31613# XM3/a_n100_82901# 1.17e-19
C4892 XM1/a_100_n179382# XM2/a_n100_n332115# 0.005074f
C4893 XM1/a_n100_156545# XM4/w_n358_n132787# 0.012279f
C4894 XM1/a_100_n136302# XM3/a_n100_n84931# 5.71e-20
C4895 XM1/a_n100_n58855# XM3/a_n100_n7231# 9.5e-19
C4896 XM1/a_n158_n24294# XM3/a_n100_26957# 3.89e-20
C4897 XM1/a_n158_120742# XM2/a_n158_n34150# 4.64e-21
C4898 XM1/a_n100_68949# m1_1634_n2388# 9.31e-20
C4899 XM2/a_n158_n247666# XM3/a_n100_n41419# 1.18e-19
C4900 XM4/w_n358_n132787# XM4/a_n100_n24843# -0.004445f
C4901 XM1/a_100_n5626# XM2/a_100_n158042# 4.64e-21
C4902 XM1/a_100_4426# XM4/w_n358_n132787# 0.048442f
C4903 XM1/a_n100_n156503# XM2/a_n158_n310930# 0.010147f
C4904 XM1/a_100_n98966# XM4/w_n358_n132787# 0.048442f
C4905 XM3/a_n100_48713# XM4/a_n100_48713# 0.009521f
C4906 XM1/a_n100_41665# XM2/a_n100_n110691# 0.001461f
C4907 XM4/a_100_80926# m1_1634_n2388# 6.1e-20
C4908 XM1/a_100_n78862# XM2/a_n100_n234583# 0.005074f
C4909 XM1/a_100_113562# XM2/a_n100_n39519# 0.005074f
C4910 XM1/a_100_n25730# XM3/a_n158_24982# 0.004082f
C4911 XM4/w_n358_n132787# XM3/a_n100_74613# 0.007706f
C4912 XM1/a_n100_22997# m1_1634_n2388# 5.75e-19
C4913 XM1/a_100_56122# XM3/a_n100_106729# 2.85e-20
C4914 XM3/a_n100_n99435# m1_1634_n2388# 0.072015f
C4915 XM4/w_n358_n132787# XM2/a_n100_n197679# 0.023772f
C4916 XM1/a_100_n129122# XM2/a_n158_n281934# 0.040138f
C4917 XM2/a_n100_n242491# XM3/a_n158_n35106# 1.93e-19
C4918 XM2/a_n100_n316299# m1_1634_n2388# 7.61e-19
C4919 XM1/a_n100_n40187# XM2/a_n100_n192407# 5.6e-19
C4920 XM4/w_n358_n132787# XM3/a_n100_19705# 0.009119f
C4921 XM1/a_n158_172438# XM2/a_n158_18570# 9.28e-21
C4922 XM1/a_100_n42962# XM3/a_n100_9345# 2.82e-20
C4923 XM1/a_100_173874# XM2/a_n158_21206# 0.026117f
C4924 XM1/a_n158_n120506# XM2/a_n158_n274026# 4.64e-21
C4925 XM4/w_n358_n132787# XM3/a_n100_115017# 0.008259f
C4926 XM1/a_n158_n107582# XM3/a_n100_n56959# 1.62e-20
C4927 XM2/a_n158_n321474# XM3/a_n100_n117047# 7.26e-20
C4928 XM4/w_n358_n132787# XM3/a_n100_n5159# 0.009186f
C4929 XM1/a_n100_n133527# XM3/a_n158_n81726# 2.85e-20
C4930 XM1/a_n100_n2851# XM3/a_n100_48713# 7.07e-19
C4931 XM1/a_n158_34582# XM2/a_n100_n118599# 7.26e-20
C4932 XM1/a_100_11606# XM3/a_n100_62181# 2.85e-20
C4933 XM1/a_100_n182254# XM2/a_n100_n334751# 0.005074f
C4934 XM1/a_100_n87478# XM3/a_n100_n36239# 5.71e-20
C4935 XM1/a_n100_n80395# XM3/a_n100_n27951# 5.72e-19
C4936 XM1/a_100_158078# XM2/a_n158_2754# 0.065842f
C4937 XM4/w_n358_n132787# XM4/a_n100_n64211# -0.004445f
C4938 XM3/a_n158_n35106# m1_1634_n2388# 6.1e-20
C4939 XM1/a_n100_n54547# XM3/a_n158_n1954# 1.09e-21
C4940 XM2/a_100_n276662# XM3/a_n158_n70330# 0.077916f
C4941 XM2/a_n158_n73690# XM4/w_n358_n132787# 0.107093f
C4942 XM2/a_n100_n282031# XM4/a_100_n75510# 6.33e-21
C4943 XM4/a_100_41558# m1_1634_n2388# 6.1e-20
C4944 XM2/a_100_n318838# XM3/a_n100_n111867# 0.005074f
C4945 XM1/a_n158_n31474# XM2/a_n158_n187038# 4.64e-21
C4946 XM1/a_100_118# XM3/a_n158_51918# 0.002495f
C4947 XM1/a_n100_n30135# XM4/w_n358_n132787# 0.01363f
C4948 XM1/a_n158_79098# XM2/a_n100_n76423# 7.26e-20
C4949 XM2/a_n158_n229214# XM3/a_n100_n23807# 1.45e-19
C4950 XM1/a_100_n60194# XM2/a_n158_n213398# 0.078305f
C4951 XM3/a_n100_58037# m1_1634_n2388# 0.072015f
C4952 XM2/a_n100_n208223# XM3/a_n158_n918# 0.004917f
C4953 XM4/w_n358_n132787# XM2/a_n158_n134318# 0.107093f
C4954 XM2/a_n100_n168683# XM4/a_100_38450# 2.56e-20
C4955 XM4/a_n100_104657# m1_1634_n2388# 0.072015f
C4956 XM4/w_n358_n132787# XM3/a_n158_99574# 0.032295f
C4957 XM1/a_100_21658# XM2/a_100_n131682# 4.64e-21
C4958 XM1/a_n100_n167991# m1_1634_n2388# 7.81e-20
C4959 XM4/w_n358_n132787# XM2/a_n100_n321571# 0.025185f
C4960 XM4/w_n358_n132787# XM3/a_n100_n44527# 0.00903f
C4961 XM1/a_n100_n91883# XM2/a_100_n245030# 7.26e-20
C4962 XM4/a_100_n29926# m1_1634_n2388# 6.1e-20
C4963 XM1/a_n158_n152098# XM3/a_n100_n101507# 1.94e-20
C4964 XM1/a_100_n47270# XM3/a_n100_4165# 4.93e-20
C4965 XM2/a_n100_n224039# XM3/a_n158_n17494# 0.001457f
C4966 XM1/a_n100_58897# XM2/a_n158_n94778# 0.010147f
C4967 XM4/w_n358_n132787# XM4/a_n100_n103579# -0.004445f
C4968 XM3/a_n158_n74474# m1_1634_n2388# 6.1e-20
C4969 XM4/w_n358_n132787# XM3/a_n158_44666# 0.032295f
C4970 XM1/a_100_53250# XM4/w_n358_n132787# 0.055208f
C4971 XM2/a_n158_n107958# XM3/a_n158_98538# 4.64e-21
C4972 XM2/a_100_n78962# XM3/a_n158_127546# 0.0674f
C4973 XM1/a_n100_61769# XM4/w_n358_n132787# 0.013398f
C4974 XM1/a_n100_n176607# XM2/a_100_n329382# 7.26e-20
C4975 XM1/a_n158_n165022# XM2/a_n158_n318838# 9.28e-21
C4976 XM1/a_100_n86042# XM2/a_n158_n239758# 0.116862f
C4977 XM1/a_n100_84745# XM2/a_n158_n71054# 0.005074f
C4978 XM1/a_n158_n140610# XM2/a_n158_n295114# 9.28e-21
C4979 XM1/a_n100_n101935# XM4/w_n358_n132787# 0.013347f
C4980 XM1/a_100_n53014# XM3/a_n158_n918# 0.00514f
C4981 XM1/a_100_89150# XM2/a_n100_n65879# 0.005074f
C4982 XM4/a_n100_n132587# m1_1634_n2388# 0.036019f
C4983 XM1/a_n158_n110454# XM2/a_n100_n266215# 7.26e-20
C4984 XM2/a_100_n258210# XM3/a_n158_n52718# 0.077916f
C4985 XM1/a_100_n67374# XM3/a_n100_n16555# 2.85e-20
C4986 XM1/a_100_n144918# XM2/a_n100_n297847# 0.005074f
C4987 XM2/a_100_n300386# XM3/a_n100_n94255# 0.010147f
C4988 XM1/a_100_15914# XM4/w_n358_n132787# 0.054609f
C4989 XM1/a_n100_n132091# XM2/a_n158_n284570# 0.005074f
C4990 XM1/a_100_n63066# XM2/a_n158_n216034# 0.055327f
C4991 XM2/a_100_n189674# m1_1634_n2388# 0.019131f
C4992 XM4/a_n100_65289# m1_1634_n2388# 0.072015f
C4993 XM2/a_n100_n297847# XM3/a_n158_n93122# 0.005074f
C4994 XM4/w_n358_n132787# XM3/a_n100_n83895# 0.008899f
C4995 XM4/a_100_n69294# m1_1634_n2388# 6.1e-20
C4996 XM4/w_n358_n132787# XM2/a_n158_n258210# 0.101988f
C4997 XM1/a_n158_n93222# XM3/a_n100_n42455# 1.94e-20
C4998 XM2/a_n158_n210762# XM3/a_n100_n6195# 7.26e-20
C4999 XM1/a_n100_122081# XM2/a_100_n31514# 1.41e-19
C5000 XM3/a_n158_82998# m1_1634_n2388# 6.1e-20
C5001 XM3/a_n158_n113842# m1_1634_n2388# 6.1e-20
C5002 XM1/a_n158_46070# XM3/a_n100_97405# 3.89e-20
C5003 XM3/a_n158_n2990# m1_1634_n2388# 6.1e-20
C5004 XM2/a_n158_n295114# XM3/a_n158_n87942# 4.64e-21
C5005 XM3/a_n158_28090# m1_1634_n2388# 6.1e-20
C5006 XM1/a_n100_153673# XM2/a_n100_21# 0.001471f
C5007 XM3/a_n100_16597# XM4/a_n100_16597# 0.009521f
C5008 XM1/a_n100_80437# XM4/w_n358_n132787# 0.012786f
C5009 XM2/a_n100_n184499# XM3/a_n100_22813# 0.005368f
C5010 XM1/a_n158_n124814# XM3/a_n100_n72499# 1.7e-20
C5011 XM1/a_n100_163725# XM4/w_n358_n132787# 0.012279f
C5012 XM1/a_100_160950# XM2/a_n158_8026# 0.051043f
C5013 XM4/w_n358_n132787# XM3/a_n158_n19566# 0.03921f
C5014 XM4/a_n100_n6195# m1_1634_n2388# 0.072015f
C5015 XM2/a_n100_n247763# XM3/a_n100_n41419# 0.001266f
C5016 XM1/a_100_n5626# XM2/a_n158_n158042# 0.001581f
C5017 XM2/a_n158_29114# XM1/a_n100_182393# 0.005074f
C5018 XM2/a_n100_29017# XM1/a_n158_182490# 7.26e-20
C5019 XM1/a_100_n116198# XM2/a_100_n271390# 4.64e-21
C5020 XM2/a_100_n202854# XM3/a_n100_4165# 0.005074f
C5021 XM4/a_n100_25921# m1_1634_n2388# 0.072015f
C5022 XM1/a_100_n9934# XM2/a_n100_n166047# 0.004756f
C5023 XM4/w_n358_n132787# XM3/a_n100_n123263# 0.009186f
C5024 XM4/a_100_n108662# m1_1634_n2388# 6.1e-20
C5025 XM1/a_100_n78862# XM2/a_100_n231850# 4.64e-21
C5026 XM1/a_n100_155109# XM2/a_n158_118# 0.005074f
C5027 XM2/a_n100_n129143# m1_1634_n2388# 0.001163f
C5028 XM1/a_n100_n74651# XM4/w_n358_n132787# 0.01363f
C5029 XM4/w_n358_n132787# XM2/a_100_n194946# 0.103342f
C5030 XM1/a_100_n129122# XM2/a_n100_n282031# 0.005074f
C5031 XM2/a_n100_n245127# XM4/a_100_n40286# 1.48e-20
C5032 XM2/a_100_n239758# XM3/a_n158_n35106# 0.063506f
C5033 XM1/a_100_n35782# XM2/a_n158_n189674# 0.116862f
C5034 XM2/a_100_n313566# m1_1634_n2388# 0.020684f
C5035 XM4/w_n358_n132787# XM4/a_n100_120197# -0.004445f
C5036 XM1/a_100_27402# XM3/a_n100_78757# 5.71e-20
C5037 XM2/a_100_n281934# XM3/a_n100_n76643# 0.010147f
C5038 XM1/a_n158_n120506# XM2/a_n100_n274123# 6.38e-20
C5039 XM1/a_n158_n48706# XM2/a_n158_n202854# 9.28e-21
C5040 XM2/a_n100_n73787# XM4/a_100_130654# 2.56e-20
C5041 XM1/a_n100_18689# XM3/a_n158_70566# 2.85e-20
C5042 XM1/a_n158_n144918# XM3/a_n100_n93219# 6.61e-21
C5043 XM4/w_n358_n132787# XM3/a_n158_n58934# 0.038462f
C5044 XM4/a_n100_n45563# m1_1634_n2388# 0.072015f
C5045 XM1/a_100_n50142# XM3/a_n158_1154# 0.00544f
C5046 XM2/a_n158_n318838# XM3/a_n100_n111867# 7.26e-20
C5047 XM1/a_n158_n31474# XM2/a_n100_n187135# 7.26e-20
C5048 XM1/a_n100_n159375# XM3/a_n158_n108662# 2.85e-20
C5049 XM1/a_n100_n175171# XM3/a_n158_n124202# 2.85e-20
C5050 XM1/a_100_n31474# XM3/a_n100_20741# 2.85e-20
C5051 XM4/w_n358_n132787# XM3/a_n100_93261# 0.008158f
C5052 XM1/a_100_n60194# XM2/a_n100_n213495# 0.005074f
C5053 XM1/a_n100_n22955# XM4/w_n358_n132787# 0.013358f
C5054 XM1/a_n100_n103371# m1_1634_n2388# 3.43e-19
C5055 XM2/a_100_n205490# XM3/a_n158_n918# 0.055716f
C5056 XM4/w_n358_n132787# XM4/a_n100_80829# -0.004445f
C5057 XM1/a_n158_25966# XM2/a_n158_n129046# 4.64e-21
C5058 XM4/w_n358_n132787# XM2/a_n100_n134415# 0.025779f
C5059 XM2/a_n100_n253035# m1_1634_n2388# 0.002555f
C5060 XM3/a_n100_n25879# m1_1634_n2388# 0.072015f
C5061 XM4/w_n358_n132787# XM3/a_n100_38353# 0.009055f
C5062 XM3/a_n100_3129# m1_1634_n2388# 0.072015f
C5063 XM2/a_100_n110594# XM3/a_n100_93261# 0.003644f
C5064 XM4/w_n358_n132787# XM2/a_100_n318838# 0.106157f
C5065 XM1/a_100_21658# XM2/a_n158_n131682# 0.091547f
C5066 XM4/w_n358_n132787# XM3/a_n158_n98302# 0.034127f
C5067 XM4/a_n100_n84931# m1_1634_n2388# 0.072015f
C5068 XM1/a_n100_n91883# XM2/a_n158_n245030# 0.005074f
C5069 XM1/a_n100_n87575# XM2/a_100_n242394# 7.26e-20
C5070 XM1/a_n100_n71779# XM2/a_n100_n224039# 0.004619f
C5071 XM2/a_n100_n226675# XM4/a_100_n22674# 2.64e-22
C5072 XM1/a_100_n61630# XM4/w_n358_n132787# 0.048442f
C5073 XM1/a_n158_n150662# XM3/a_n158_n98302# 1.14e-21
C5074 XM2/a_100_n263482# XM3/a_n100_n59031# 0.005074f
C5075 XM2/a_n100_n108055# XM3/a_n158_98538# 0.005055f
C5076 XM1/a_n158_n169330# XM3/a_n100_n119119# 1e-21
C5077 XM1/a_n100_n107679# m1_1634_n2388# 1.3e-19
C5078 XM2/a_n158_n78962# XM3/a_n158_127546# 4.64e-21
C5079 XM2/a_100_n78962# XM3/a_n100_127449# 0.005074f
C5080 XM1/a_n158_n87478# XM2/a_n158_n242394# 4.64e-21
C5081 XM1/a_n158_159514# XM2/a_n158_5390# 9.28e-21
C5082 XM2/a_n158_n26242# XM4/w_n358_n132787# 0.107093f
C5083 XM1/a_100_94894# XM4/w_n358_n132787# 0.053546f
C5084 sw_b iout_n 0.001928f
C5085 XM1/a_n100_n176607# XM2/a_n158_n329382# 0.005074f
C5086 XM2/a_n100_n15795# XM1/a_100_139410# 0.005074f
C5087 XM4/a_100_115114# m1_1634_n2388# 6.1e-20
C5088 XM1/a_100_n74554# XM4/w_n358_n132787# 0.048442f
C5089 XM1/a_n158_160950# XM2/a_n158_8026# 4.64e-21
C5090 XM4/a_n100_7273# m1_1634_n2388# 0.072015f
C5091 XM4/w_n358_n132787# XM4/a_n100_41461# -0.004445f
C5092 XM2/a_n100_n113327# XM4/a_100_91286# 2.56e-20
C5093 XM1/a_n158_n116198# XM3/a_n100_n65247# 1.94e-20
C5094 XM1/a_n100_87617# XM2/a_100_n65782# 7.26e-20
C5095 XM3/a_n100_76685# m1_1634_n2388# 0.072015f
C5096 XM3/a_n100_n65247# m1_1634_n2388# 0.072015f
C5097 XM2/a_n158_n300386# XM3/a_n100_n94255# 1.45e-19
C5098 XM1/a_100_n63066# XM2/a_n100_n216131# 0.005074f
C5099 XM1/a_n100_43101# XM4/w_n358_n132787# 0.013334f
C5100 XM3/a_n100_69433# XM4/a_n100_69433# 0.009521f
C5101 XM2/a_n158_n189674# m1_1634_n2388# 2.36e-21
C5102 XM4/a_n100_n124299# m1_1634_n2388# 0.072015f
C5103 XM1/a_100_n32910# XM3/a_n100_17633# 2.85e-20
C5104 XM3/a_n100_21777# m1_1634_n2388# 0.072015f
C5105 XM4/w_n358_n132787# XM2/a_n100_n258307# 0.025738f
C5106 XM3/a_n100_n14483# XM4/a_n100_n14483# 0.009521f
C5107 XM1/a_n158_81970# XM2/a_n158_n71054# 4.64e-21
C5108 XM3/a_n158_118222# m1_1634_n2388# 6.1e-20
C5109 XM1/a_n100_43101# XM2/a_100_n110594# 1.45e-19
C5110 XM1/a_100_n45834# XM2/a_n158_n200218# 0.116862f
C5111 XM2/a_100_n139590# XM3/a_n100_65289# 0.010147f
C5112 XM4/w_n358_n132787# XM3/a_n158_63314# 0.032295f
C5113 XM2/a_n100_n295211# XM3/a_n158_n87942# 0.005074f
C5114 XM4/w_n358_n132787# XM4/a_n100_n30023# -0.004445f
C5115 XM1/a_n100_n12903# XM2/a_100_n168586# 7.26e-20
C5116 XM1/a_n100_n2851# XM2/a_100_n158042# 7.26e-20
C5117 XM1/a_n100_n106243# XM2/a_100_n260846# 1.45e-19
C5118 XM2/a_100_n181766# XM3/a_n100_22813# 0.005074f
C5119 XM2/a_n158_21206# XM4/w_n358_n132787# 0.107093f
C5120 XM1/a_n100_n77523# XM4/w_n358_n132787# 0.013462f
C5121 XM4/a_100_75746# m1_1634_n2388# 6.1e-20
C5122 XM1/a_100_148026# XM2/a_n158_n5154# 0.075968f
C5123 XM1/a_n100_n129219# XM2/a_100_n284570# 7.26e-20
C5124 XM1/a_100_n84606# XM3/a_n100_n34167# 2.85e-20
C5125 XM3/a_n100_n104615# m1_1634_n2388# 0.072015f
C5126 XM1/a_n100_n143579# XM2/a_100_n297750# 1.45e-19
C5127 XM2/a_n158_n202854# XM3/a_n100_4165# 7.26e-20
C5128 XM1/a_100_n5626# XM2/a_n100_n158139# 0.005074f
C5129 XM1/a_100_n159278# XM4/w_n358_n132787# 0.048442f
C5130 XM1/a_100_n116198# XM2/a_n158_n271390# 0.078695f
C5131 XM2/a_n100_n179227# XM3/a_n158_28090# 0.004675f
C5132 XM1/a_n100_117773# XM2/a_100_n36786# 1.45e-19
C5133 XM1/a_100_n9934# XM2/a_100_n163314# 4.64e-21
C5134 XM2/a_n158_n7790# XM1/a_100_145154# 0.05299f
C5135 XM2/a_n100_n7887# XM1/a_n158_145154# 7.26e-20
C5136 XM1/a_n100_35921# XM2/a_100_n118502# 1.45e-19
C5137 XM2/a_100_n329382# XM3/a_n158_n123166# 0.077916f
C5138 XM1/a_100_n78862# XM2/a_n158_n231850# 0.057274f
C5139 XM3/a_n100_n34167# XM4/a_n100_n34167# 0.009521f
C5140 XM1/a_100_n12806# XM4/w_n358_n132787# 0.054609f
C5141 XM2/a_100_n126410# m1_1634_n2388# 0.020445f
C5142 XM1/a_100_n51578# XM2/a_n158_n205490# 0.116862f
C5143 XM1/a_100_n8498# XM3/a_n158_43630# 6.06e-19
C5144 XM1/a_n100_162289# XM4/w_n358_n132787# 0.012279f
C5145 XM1/a_n158_60430# XM3/a_n100_111909# 2.42e-20
C5146 XM4/w_n358_n132787# XM2/a_n158_n194946# 0.101988f
C5147 XM2/a_n158_n13062# XM1/a_100_142282# 0.063895f
C5148 XM2/a_100_n13062# XM1/a_n100_140749# 1.45e-19
C5149 XM2/a_n158_n239758# XM3/a_n158_n35106# 4.64e-21
C5150 XM4/w_n358_n132787# XM3/a_n100_n10339# 0.009186f
C5151 XM2/a_n158_23842# XM1/a_100_179618# 0.021833f
C5152 XM1/a_n158_110690# XM2/a_n158_n42058# 4.64e-21
C5153 XM2/a_n158_n313566# m1_1634_n2388# 2.36e-21
C5154 XM1/a_n158_n127686# XM2/a_n158_n281934# 9.28e-21
C5155 XM1/a_n100_n183787# m1_1634_n2388# 6.48e-20
C5156 XM2/a_n158_n281934# XM3/a_n100_n76643# 1.45e-19
C5157 XM2/a_100_n126410# XM3/a_n100_79793# 0.010147f
C5158 XM4/w_n358_n132787# XM4/a_n100_n69391# -0.004445f
C5159 XM3/a_n158_n40286# m1_1634_n2388# 6.1e-20
C5160 XM4/w_n358_n132787# XM3/a_n158_116150# 0.032295f
C5161 XM1/a_100_18786# XM3/a_n158_69530# 0.001549f
C5162 XM3/a_n158_46738# m1_1634_n2388# 6.1e-20
C5163 XM1/a_100_110690# XM2/a_n100_n42155# 0.005074f
C5164 XM1/a_100_31710# XM4/w_n358_n132787# 0.054609f
C5165 XM4/a_100_36378# m1_1634_n2388# 6.1e-20
C5166 XM2/a_n100_n242491# XM4/a_100_n35106# 2.37e-21
C5167 XM2/a_100_n237122# XM3/a_n158_n29926# 4.13e-19
C5168 XM2/a_100_n168586# XM3/a_n100_37317# 0.010147f
C5169 XM1/a_100_150898# XM2/a_n100_n2615# 0.005074f
C5170 XM1/a_n158_n9934# XM3/a_n100_40425# 1.12e-20
C5171 XM2/a_n100_n97511# XM3/a_n100_109837# 0.003753f
C5172 XM2/a_100_n94778# XM3/a_n158_109934# 0.069348f
C5173 XM1/a_100_n162150# XM3/a_n100_n109795# 1.4e-20
C5174 XM1/a_n100_163725# XM2/a_100_8026# 7.26e-20
C5175 XM1/a_n100_n127783# m1_1634_n2388# 1.05e-19
C5176 XM3/a_n100_n53851# XM4/a_n100_n53851# 0.009521f
C5177 XM1/a_n100_101977# XM4/w_n358_n132787# 0.012279f
C5178 XM1/a_n100_67513# XM3/a_n158_118222# 2.85e-20
C5179 XM1/a_100_100638# XM2/a_100_n55238# 4.64e-21
C5180 XM4/a_n100_99477# m1_1634_n2388# 0.072015f
C5181 XM1/a_n158_64738# XM3/a_n100_115017# 1.46e-20
C5182 XM4/w_n358_n132787# XM3/a_n100_n49707# 0.009186f
C5183 XM4/a_100_n35106# m1_1634_n2388# 6.1e-20
C5184 XM2/a_n158_n205490# XM3/a_n158_n918# 4.64e-21
C5185 XM1/a_n100_64641# XM3/a_n158_117186# 1.52e-20
C5186 XM1/a_n158_25966# XM2/a_n100_n129143# 7.26e-20
C5187 XM4/w_n358_n132787# XM2/a_100_n131682# 0.103404f
C5188 XM1/a_n100_10073# m1_1634_n2388# 1.27e-19
C5189 XM1/a_100_77662# XM2/a_n158_n76326# 0.116862f
C5190 XM4/w_n358_n132787# XM4/a_n100_n108759# -0.004445f
C5191 XM3/a_n158_n79654# m1_1634_n2388# 6.1e-20
C5192 XM2/a_100_n250302# m1_1634_n2388# 0.01937f
C5193 XM1/a_n158_n58758# XM3/a_n100_n7231# 1.94e-20
C5194 XM1/a_100_152334# XM2/a_n158_n2518# 0.111799f
C5195 XM2/a_100_n310930# XM3/a_n158_n105554# 0.077916f
C5196 XM1/a_n100_91925# XM2/a_n158_n60510# 0.005074f
C5197 XM2/a_n158_n110594# XM3/a_n100_93261# 4.06e-20
C5198 XM4/w_n358_n132787# XM2/a_n158_n318838# 0.106642f
C5199 XM1/a_100_21658# XM2/a_n100_n131779# 0.005074f
C5200 XM1/a_n100_n87575# XM2/a_n158_n242394# 0.005074f
C5201 XM2/a_n100_n42155# XM4/w_n358_n132787# 0.012279f
C5202 XM1/a_n158_n121942# XM3/a_n100_n70427# 1.94e-20
C5203 XM1/a_n100_n41623# XM4/w_n358_n132787# 0.01278f
C5204 XM2/a_n158_n263482# XM3/a_n100_n59031# 7.26e-20
C5205 XM2/a_n100_n79059# XM3/a_n158_127546# 0.005074f
C5206 XM2/a_n158_n78962# XM3/a_n100_127449# 7.26e-20
C5207 XM1/a_n158_n87478# XM2/a_n100_n242491# 7.26e-20
C5208 XM2/a_100_n197582# XM3/a_n100_9345# 0.005074f
C5209 XM3/a_n100_37317# XM4/a_n100_37317# 0.009521f
C5210 XM1/a_n100_n167991# XM3/a_n158_n115914# 2.85e-20
C5211 XM3/a_n100_n73535# XM4/a_n100_n73535# 0.009521f
C5212 XM1/a_n158_166694# XM2/a_n158_13298# 4.64e-21
C5213 XM2/a_n100_n224039# XM4/a_100_n17494# 1.27e-20
C5214 XM2/a_100_n218670# XM3/a_n158_n12314# 0.077916f
C5215 XM1/a_100_18786# XM4/w_n358_n132787# 0.055022f
C5216 XM4/a_n100_60109# m1_1634_n2388# 0.072015f
C5217 XM4/w_n358_n132787# XM3/a_n100_n89075# 0.008979f
C5218 XM4/a_100_n74474# m1_1634_n2388# 6.1e-20
C5219 XM2/a_100_n260846# XM3/a_n100_n53851# 0.005074f
C5220 XM1/a_100_48942# XM3/a_n100_99477# 2.85e-20
C5221 XM1/a_n158_n110454# XM2/a_n158_n263482# 4.64e-21
C5222 XM1/a_100_n109018# XM2/a_n158_n263482# 0.116862f
C5223 XM1/a_100_n71682# XM3/a_n100_n20699# 2.85e-20
C5224 XM3/a_n158_n119022# m1_1634_n2388# 6.1e-20
C5225 XM1/a_n158_n60194# XM3/a_n100_n9303# 1.94e-20
C5226 XM2/a_n100_n189771# m1_1634_n2388# 0.002489f
C5227 XM1/a_100_158078# XM2/a_100_5390# 4.64e-21
C5228 XM4/w_n358_n132787# XM3/a_n100_57001# 0.008281f
C5229 XM4/w_n358_n132787# XM2/a_100_n255574# 0.105283f
C5230 XM2/a_n100_n110691# XM4/a_100_96466# 2.56e-20
C5231 XM4/w_n358_n132787# XM1/a_n100_n143579# 0.013401f
C5232 XM1/a_n100_166597# XM4/w_n358_n132787# 0.011792f
C5233 XM3/a_n100_118125# m1_1634_n2388# 0.072015f
C5234 XM1/a_n100_43101# XM2/a_n158_n110594# 0.010147f
C5235 XM4/w_n358_n132787# XM3/a_n158_n24746# 0.038462f
C5236 XM4/a_n100_n11375# m1_1634_n2388# 0.072015f
C5237 XM1/a_n158_61866# XM2/a_n158_n92142# 9.28e-21
C5238 XM2/a_n158_n139590# XM3/a_n100_65289# 1.45e-19
C5239 XM4/w_n358_n132787# XM1/a_n100_n133527# 0.01363f
C5240 XM1/a_100_37454# XM3/a_n100_89117# 2.85e-20
C5241 XM2/a_100_n292478# XM3/a_n158_n87942# 0.052211f
C5242 XM1/a_n100_n84703# m1_1634_n2388# 9.43e-20
C5243 XM2/a_n100_n297847# XM4/a_100_n93122# 2.56e-20
C5244 XM3/a_n100_n93219# XM4/a_n100_n93219# 0.009521f
C5245 XM1/a_n100_n12903# XM2/a_n158_n168586# 0.005074f
C5246 XM1/a_n100_n2851# XM2/a_n158_n158042# 0.005074f
C5247 XM2/a_100_n334654# XM3/a_n100_n129479# 0.010147f
C5248 XM1/a_n100_n106243# XM2/a_n158_n260846# 0.010147f
C5249 XM2/a_n158_n181766# XM3/a_n100_22813# 7.26e-20
C5250 XM1/a_n100_n24391# XM2/a_100_n179130# 7.26e-20
C5251 XM4/a_n100_20741# m1_1634_n2388# 0.072015f
C5252 XM1/a_n158_33146# XM3/a_n100_84973# 1.94e-20
C5253 XM4/w_n358_n132787# XM3/a_n100_n128443# 0.008845f
C5254 XM4/a_100_n113842# m1_1634_n2388# 6.1e-20
C5255 XM1/a_n100_n110551# XM2/a_100_n266118# 7.26e-20
C5256 XM1/a_100_119306# XM2/a_100_n34150# 4.64e-21
C5257 XM2/a_100_n134318# XM3/a_n158_70566# 0.077916f
C5258 XM1/a_n100_n15775# XM4/w_n358_n132787# 0.01363f
C5259 XM1/a_n100_n129219# XM2/a_n158_n284570# 0.005074f
C5260 XM1/a_100_n96094# XM4/w_n358_n132787# 0.048442f
C5261 XM1/a_n100_n143579# XM2/a_n158_n297750# 0.010147f
C5262 XM1/a_100_28838# XM3/a_n100_80829# 4.7e-19
C5263 XM1/a_100_n116198# XM2/a_n100_n271487# 0.005074f
C5264 XM2/a_100_n176494# XM3/a_n158_28090# 0.056885f
C5265 XM3/a_n100_95333# m1_1634_n2388# 0.072015f
C5266 XM1/a_100_n9934# XM2/a_n158_n163314# 0.095442f
C5267 XM4/w_n358_n132787# XM4/a_n100_115017# -0.004445f
C5268 XM1/a_n100_35921# XM2/a_n158_n118502# 0.010147f
C5269 XM1/a_100_n78862# XM2/a_n100_n231947# 0.005074f
C5270 XM1/a_n158_113562# XM2/a_n158_n39422# 4.64e-21
C5271 XM2/a_n158_n126410# m1_1634_n2388# 2.36e-21
C5272 XM1/a_100_n166458# XM2/a_100_n321474# 4.64e-21
C5273 XM1/a_n100_n136399# XM3/a_n100_n83895# 0.001171f
C5274 XM1/a_100_104946# XM4/w_n358_n132787# 0.05072f
C5275 XM1/a_n158_25966# XM3/a_n100_76685# 1.94e-20
C5276 XM1/a_n100_20125# XM3/a_n158_72638# 2.46e-20
C5277 XM2/a_100_n242394# XM3/a_n100_n36239# 0.010147f
C5278 XM3/a_n100_40425# m1_1634_n2388# 0.072015f
C5279 XM1/a_100_56122# XM3/a_n100_107765# 2.85e-20
C5280 XM4/w_n358_n132787# XM2/a_n100_n195043# 0.025193f
C5281 XM3/a_n100_125377# XM4/a_n100_125377# 0.009521f
C5282 XM4/w_n358_n132787# XM3/a_n158_n64114# 0.036903f
C5283 XM1/a_n158_n113326# XM2/a_n158_n268754# 4.64e-21
C5284 XM4/a_n100_n50743# m1_1634_n2388# 0.072015f
C5285 XM2/a_n100_n239855# XM3/a_n158_n35106# 0.005074f
C5286 XM1/a_n158_n167894# XM3/a_n158_n116950# 1.14e-21
C5287 XM2/a_n100_n313663# m1_1634_n2388# 0.001179f
C5288 XM1/a_n158_77662# XM2/a_n158_n76326# 9.28e-21
C5289 XM4/w_n358_n132787# XM3/a_n158_81962# 0.032295f
C5290 XM2/a_n158_n126410# XM3/a_n100_79793# 1.45e-19
C5291 XM3/a_n100_n112903# XM4/a_n100_n112903# 0.009521f
C5292 XM4/w_n358_n132787# XM3/a_n100_116053# 0.009186f
C5293 XM1/a_n100_n37315# m1_1634_n2388# 1.3e-19
C5294 XM2/a_n158_n237122# XM3/a_n158_n29926# 4.64e-21
C5295 XM2/a_n158_n168586# XM3/a_n100_37317# 1.45e-19
C5296 XM1/a_n100_n169427# XM3/a_n158_n119022# 2.27e-21
C5297 XM4/w_n358_n132787# XM3/a_n158_27054# 0.032295f
C5298 XM1/a_100_n104710# XM4/w_n358_n132787# 0.050569f
C5299 XM2/a_100_n20970# XM1/a_100_132230# 4.64e-21
C5300 XM2/a_100_n121138# XM3/a_n158_85070# 0.077916f
C5301 XM3/a_n100_n1015# XM4/a_n100_n1015# 0.009521f
C5302 XM1/a_n158_169566# XM2/a_n158_15934# 9.28e-21
C5303 XM2/a_100_n94778# XM3/a_n100_109837# 0.005074f
C5304 XM2/a_n158_n94778# XM3/a_n158_109934# 4.64e-21
C5305 XM1/a_100_n2754# XM3/a_n100_48713# 3.99e-20
C5306 XM4/w_n358_n132787# XM4/a_n100_75649# -0.004445f
C5307 XM2/a_100_n316202# XM3/a_n100_n111867# 0.005074f
C5308 XM1/a_n158_n31474# XM2/a_n158_n184402# 4.64e-21
C5309 XM2/a_100_n163314# XM3/a_n158_42594# 0.077916f
C5310 XM1/a_100_79098# XM2/a_100_n76326# 4.64e-21
C5311 XM3/a_n100_n31059# m1_1634_n2388# 0.072015f
C5312 XM3/a_n100_1057# XM4/a_n100_1057# 0.009521f
C5313 XM1/a_n100_24433# XM4/w_n358_n132787# 0.013171f
C5314 XM1/a_100_69046# XM3/a_n158_120294# 0.00544f
C5315 XM4/w_n358_n132787# XM3/a_n158_n103482# 0.032295f
C5316 XM4/a_n100_n90111# m1_1634_n2388# 0.072015f
C5317 XM2/a_n100_n205587# XM3/a_n158_n918# 0.005074f
C5318 XM2/a_n158_23842# XM1/a_n100_178085# 0.010147f
C5319 XM1/a_n100_64641# XM3/a_n100_117089# 6.24e-19
C5320 XM4/w_n358_n132787# XM2/a_n158_n131682# 0.102535f
C5321 XM1/a_100_n175074# XM4/w_n358_n132787# 0.048442f
C5322 XM1/a_n100_n110551# XM3/a_n100_n57995# 4.94e-19
C5323 XM1/a_n158_n74554# XM3/a_n100_n23807# 1.94e-20
C5324 XM4/w_n358_n132787# XM3/a_n100_8309# 0.009186f
C5325 XM2/a_n158_n250302# m1_1634_n2388# 2.36e-21
C5326 XM1/a_n158_n41526# XM3/a_n100_10381# 1.94e-20
C5327 XM2/a_n100_n166047# XM4/a_100_38450# 2.56e-20
C5328 XM1/a_n158_63302# XM2/a_n158_n92142# 4.64e-21
C5329 XM1/a_100_127922# XM2/a_n158_n26242# 0.116862f
C5330 XM2/a_n100_n110691# XM3/a_n100_93261# 0.00171f
C5331 XM3/a_n100_90153# XM4/a_n100_90153# 0.009521f
C5332 XM4/w_n358_n132787# XM2/a_n100_n318935# 0.024581f
C5333 XM2/a_100_n223942# XM3/a_n100_n18627# 0.010147f
C5334 XM1/a_n100_162289# XM2/a_100_8026# 1.45e-19
C5335 XM1/a_100_163822# XM2/a_n100_7929# 0.005074f
C5336 XM3/a_n158_65386# m1_1634_n2388# 6.1e-20
C5337 XM2/a_n100_n208223# XM4/a_100_n918# 2.35e-20
C5338 XM4/a_100_109934# m1_1634_n2388# 6.1e-20
C5339 XM1/a_n100_n159375# XM2/a_100_n313566# 1.45e-19
C5340 XM1/a_n158_n146354# XM2/a_n158_n300386# 9.28e-21
C5341 XM1/a_n100_n43059# XM4/w_n358_n132787# 0.013401f
C5342 XM1/a_n100_n153631# XM4/w_n358_n132787# 0.013508f
C5343 XM3/a_n158_10478# m1_1634_n2388# 6.1e-20
C5344 XM4/w_n358_n132787# XM4/a_n100_36281# -0.004445f
C5345 XM3/a_n100_108801# XM4/a_n100_108801# 0.009521f
C5346 XM1/a_100_n100402# XM3/a_n100_n49707# 2.85e-20
C5347 XM1/a_n158_n81734# XM3/a_n100_n30023# 1.94e-20
C5348 XM2/a_n158_n197582# XM3/a_n100_9345# 7.26e-20
C5349 XM3/a_n100_n70427# m1_1634_n2388# 0.072015f
C5350 XM1/a_100_n57322# XM2/a_n100_n213495# 0.001183f
C5351 XM1/a_100_48942# XM4/w_n358_n132787# 0.048442f
C5352 XM1/a_n100_n145015# XM3/a_n158_n93122# 2.85e-20
C5353 XM1/a_n100_n87575# m1_1634_n2388# 4.31e-20
C5354 XM1/a_100_n24294# XM3/a_n100_27993# 1.02e-19
C5355 XM4/a_n100_n129479# m1_1634_n2388# 0.072015f
C5356 XM2/a_n158_n260846# XM3/a_n100_n53851# 7.26e-20
C5357 XM1/a_100_n157842# XM3/a_n158_n106590# 0.00544f
C5358 XM1/a_n158_n110454# XM2/a_n100_n263579# 7.26e-20
C5359 XM1/a_n100_n84703# XM2/a_100_n239758# 7.26e-20
C5360 XM2/a_100_n192310# XM3/a_n158_14622# 0.026117f
C5361 XM1/a_100_125050# XM2/a_n158_n28878# 0.116862f
C5362 XM4/w_n358_n132787# XM1/a_100_137974# 0.048442f
C5363 XM1/a_n100_n134963# XM2/a_100_n289842# 7.26e-20
C5364 XM2/a_100_n187038# m1_1634_n2388# 0.017213f
C5365 XM1/a_n100_n24391# m1_1634_n2388# 3.94e-20
C5366 XM4/w_n358_n132787# XM4/a_n100_n35203# -0.004445f
C5367 XM4/w_n358_n132787# XM2/a_n158_n255574# 0.105364f
C5368 XM3/a_n158_n6098# m1_1634_n2388# 6.1e-20
C5369 XM1/a_100_11606# XM4/w_n358_n132787# 0.048442f
C5370 XM1/a_100_7298# XM2/a_n158_n147498# 0.116862f
C5371 XM4/a_100_70566# m1_1634_n2388# 6.1e-20
C5372 XM1/a_n100_n20083# XM3/a_n100_31101# 0.001054f
C5373 XM1/a_n158_36018# XM3/a_n100_88081# 1.94e-20
C5374 XM1/a_n100_86181# XM2/a_100_n68418# 1.45e-19
C5375 XM2/a_n158_n292478# XM3/a_n158_n87942# 4.64e-21
C5376 XM1/a_n100_n80395# XM4/w_n358_n132787# 0.013401f
C5377 XM1/a_100_n40090# XM3/a_n158_11514# 0.001549f
C5378 XM3/a_n100_n109795# m1_1634_n2388# 0.072015f
C5379 XM1/a_n158_n50142# XM3/a_n100_1057# 3.87e-20
C5380 XM2/a_n158_n334654# XM3/a_n100_n129479# 1.45e-19
C5381 XM1/a_n100_n24391# XM2/a_n158_n179130# 0.005074f
C5382 XM1/a_n100_n110551# XM2/a_n158_n266118# 0.005074f
C5383 XM1/a_n100_n40187# XM3/a_n158_10478# 2.85e-20
C5384 XM1/a_n158_n24294# XM3/a_n100_27993# 1.54e-20
C5385 XM1/a_n158_79098# XM2/a_n158_n73690# 4.64e-21
C5386 XM3/a_n158_4262# m1_1634_n2388# 6.1e-20
C5387 XM2/a_n100_n295211# XM4/a_100_n87942# 2.56e-20
C5388 XM2/a_100_n289842# XM3/a_n158_n82762# 0.011707f
C5389 XM1/a_100_n55886# XM4/w_n358_n132787# 0.050001f
C5390 XM1/a_100_n180818# XM3/a_n100_n128443# 8.15e-21
C5391 XM1/a_100_n98966# XM3/a_n100_n48671# 2.7e-20
C5392 XM2/a_100_n200218# XM3/a_n100_4165# 0.005074f
C5393 XM1/a_100_n116198# XM2/a_100_n268754# 4.64e-21
C5394 XM1/a_100_n100402# XM2/a_100_n255574# 4.64e-21
C5395 XM4/w_n358_n132787# XM3/a_n100_n15519# 0.009186f
C5396 XM2/a_n158_n176494# XM3/a_n158_28090# 4.64e-21
C5397 XM1/a_100_n9934# XM2/a_n100_n163411# 0.005074f
C5398 XM1/a_100_n94658# XM3/a_n158_n43394# 0.00544f
C5399 XM1/a_100_n15678# m1_1634_n2388# 3.03e-19
C5400 XM1/a_n100_n11467# XM3/a_n158_39486# 2.85e-20
C5401 XM2/a_n100_n126507# m1_1634_n2388# 0.001337f
C5402 XM4/w_n358_n132787# XM3/a_n100_75649# 0.007858f
C5403 XM1/a_100_n166458# XM2/a_n158_n321474# 0.095831f
C5404 XM4/w_n358_n132787# XM4/a_n100_n74571# -0.004445f
C5405 XM3/a_n158_n45466# m1_1634_n2388# 6.1e-20
C5406 XM2/a_n158_n242394# XM3/a_n100_n36239# 1.45e-19
C5407 XM4/w_n358_n132787# XM2/a_100_n192310# 0.103929f
C5408 XM4/a_100_31198# m1_1634_n2388# 6.1e-20
C5409 XM1/a_n100_157981# XM2/a_n158_2754# 0.005074f
C5410 XM1/a_n158_n113326# XM2/a_n100_n268851# 7.26e-20
C5411 XM1/a_100_n14242# XM2/a_n158_n168586# 0.116862f
C5412 XM2/a_100_n310930# m1_1634_n2388# 0.017213f
C5413 XM1/a_n100_n140707# XM3/a_n158_n88978# 1.02e-20
C5414 XM4/w_n358_n132787# XM3/a_n100_20741# 0.009186f
C5415 XM1/a_n100_n127783# XM3/a_n158_n76546# 1.84e-20
C5416 XM1/a_100_n120506# XM3/a_n100_n69391# 2.93e-20
C5417 XM2/a_n100_n237219# XM3/a_n158_n29926# 0.005074f
C5418 XM1/a_100_11606# XM3/a_n100_63217# 2.85e-20
C5419 XM1/a_100_106382# XM4/w_n358_n132787# 0.048442f
C5420 XM4/a_n100_94297# m1_1634_n2388# 0.072015f
C5421 XM1/a_100_n97530# XM4/w_n358_n132787# 0.054932f
C5422 XM2/a_n158_n94778# XM3/a_n100_109837# 7.26e-20
C5423 XM2/a_n100_n94875# XM3/a_n158_109934# 0.004897f
C5424 XM4/w_n358_n132787# XM3/a_n100_n54887# 0.009186f
C5425 XM4/a_100_n40286# m1_1634_n2388# 6.1e-20
C5426 XM2/a_n158_n71054# XM4/w_n358_n132787# 0.107093f
C5427 XM2/a_n158_n316202# XM3/a_n100_n111867# 7.26e-20
C5428 XM1/a_n158_n31474# XM2/a_n100_n184499# 7.26e-20
C5429 XM1/a_100_79098# XM2/a_n158_n76326# 0.056106f
C5430 XM3/a_n100_58037# XM4/a_n100_58037# 0.009521f
C5431 XM4/w_n358_n132787# XM4/a_n100_n113939# -0.004445f
C5432 XM3/a_n158_n84834# m1_1634_n2388# 6.1e-20
C5433 XM1/a_n100_n80395# XM2/a_100_n234486# 1.45e-19
C5434 XM1/a_100_63302# XM3/a_n100_113981# 2.85e-20
C5435 XM1/a_100_69046# XM3/a_n100_120197# 4.35e-20
C5436 XM2/a_100_n271390# XM3/a_n158_n65150# 0.077916f
C5437 XM3/a_n100_59073# m1_1634_n2388# 0.072015f
C5438 XM1/a_n100_n38751# XM3/a_n100_12453# 0.001668f
C5439 XM4/w_n358_n132787# XM2/a_n100_n131779# 0.0242f
C5440 XM2/a_100_n313566# XM3/a_n100_n106687# 0.005074f
C5441 XM2/a_n100_n250399# m1_1634_n2388# 0.002627f
C5442 XM1/a_100_n75990# XM4/w_n358_n132787# 0.054609f
C5443 XM1/a_n100_n106243# XM3/a_n158_n53754# 2.85e-20
C5444 XM1/a_n100_n71779# XM3/a_n158_n20602# 2.85e-20
C5445 XM1/a_n158_63302# XM2/a_n100_n92239# 7.26e-20
C5446 XM4/w_n358_n132787# XM2/a_100_n316202# 0.103341f
C5447 XM2/a_n158_n223942# XM3/a_n100_n18627# 1.45e-19
C5448 XM1/a_n100_n163683# m1_1634_n2388# 1.3e-19
C5449 XM1/a_n158_171002# XM2/a_n100_15837# 7.26e-20
C5450 XM1/a_n100_n159375# XM2/a_n158_n313566# 0.010147f
C5451 XM4/w_n358_n132787# XM3/a_n158_45702# 0.032295f
C5452 XM2/a_n100_n155503# XM3/a_n100_51821# 0.005548f
C5453 XM4/a_n100_54929# m1_1634_n2388# 0.072015f
C5454 XM4/a_100_1154# m1_1634_n2388# 6.1e-20
C5455 XM2/a_n100_n163411# XM4/a_100_43630# 2.56e-20
C5456 XM4/w_n358_n132787# XM3/a_n100_n94255# 0.009186f
C5457 XM4/a_100_n79654# m1_1634_n2388# 6.1e-20
C5458 XM1/a_n100_35921# m1_1634_n2388# 1.15e-19
C5459 XM1/a_n100_123517# XM2/a_100_n31514# 7.26e-20
C5460 XM1/a_100_90586# XM2/a_n158_n63146# 0.116862f
C5461 XM3/a_n158_n124202# m1_1634_n2388# 6.1e-20
C5462 XM1/a_100_n57322# XM2/a_100_n210762# 4.64e-21
C5463 XM1/a_n100_n166555# XM2/a_100_n321474# 7.26e-20
C5464 XM1/a_n100_84745# XM2/a_n158_n68418# 0.005074f
C5465 XM1/a_n100_n84703# XM2/a_n158_n239758# 0.005074f
C5466 XM2/a_n158_n192310# XM3/a_n158_14622# 4.64e-21
C5467 XM1/a_n158_129358# XM2/a_n100_n26339# 7.26e-20
C5468 XM1/a_100_n182254# XM3/a_n100_n131551# 2.85e-20
C5469 XM1/a_100_n176510# XM3/a_n100_n125335# 5.05e-20
C5470 XM1/a_100_n146354# XM2/a_n158_n300386# 0.116862f
C5471 XM1/a_n100_n134963# XM2/a_n158_n289842# 0.005074f
C5472 XM4/w_n358_n132787# XM3/a_n158_n29926# 0.038462f
C5473 XM4/a_n100_n16555# m1_1634_n2388# 0.072015f
C5474 XM1/a_n100_n15775# XM2/a_100_n171222# 7.26e-20
C5475 XM1/a_n100_n5723# m1_1634_n2388# 9.25e-20
C5476 XM1/a_n100_n58855# m1_1634_n2388# 8.08e-20
C5477 XM4/w_n358_n132787# XM2/a_n100_n255671# 0.024356f
C5478 XM1/a_n158_163822# XM2/a_n100_7929# 7.26e-20
C5479 XM2/a_100_n252938# XM3/a_n158_n47538# 0.077916f
C5480 XM1/a_100_n51578# XM3/a_n100_n1015# 2.85e-20
C5481 XM1/a_n158_46070# XM3/a_n100_98441# 5.81e-21
C5482 XM1/a_100_43198# XM4/w_n358_n132787# 0.048442f
C5483 XM3/a_n158_84034# m1_1634_n2388# 6.1e-20
C5484 XM4/a_n100_15561# m1_1634_n2388# 0.072014f
C5485 XM3/a_n158_119258# m1_1634_n2388# 6.1e-20
C5486 XM4/a_100_n119022# m1_1634_n2388# 6.1e-20
C5487 XM2/a_100_n295114# XM3/a_n100_n89075# 0.010147f
C5488 XM1/a_n158_168130# XM2/a_n158_13298# 4.64e-21
C5489 XM3/a_n158_n1954# m1_1634_n2388# 6.1e-20
C5490 XM2/a_n100_n292575# XM3/a_n158_n87942# 0.005074f
C5491 XM3/a_n158_29126# m1_1634_n2388# 6.1e-20
C5492 XM1/a_n100_n12903# XM2/a_100_n165950# 7.26e-20
C5493 XM1/a_n100_n2851# XM2/a_100_n155406# 7.26e-20
C5494 XM1/a_n100_n24391# XM2/a_n100_n179227# 0.003193f
C5495 XM1/a_100_76226# m1_1634_n2388# 0.002487f
C5496 XM4/w_n358_n132787# XM4/a_n100_109837# -0.004445f
C5497 XM1/a_n100_n129219# XM2/a_100_n281934# 7.26e-20
C5498 XM1/a_100_n2754# XM2/a_100_n158042# 4.64e-21
C5499 XM1/a_100_114998# XM4/w_n358_n132787# 0.048442f
C5500 XM2/a_n158_n289842# XM3/a_n158_n82762# 4.64e-21
C5501 XM1/a_100_n100402# XM2/a_n158_n255574# 0.080642f
C5502 XM2/a_n158_n200218# XM3/a_n100_4165# 7.26e-20
C5503 XM4/w_n358_n132787# XM3/a_n158_n69294# 0.033785f
C5504 XM1/a_100_n116198# XM2/a_n158_n268754# 0.015212f
C5505 XM4/a_n100_n55923# m1_1634_n2388# 0.072015f
C5506 XM2/a_n100_n176591# XM3/a_n158_28090# 0.005074f
C5507 XM2/a_100_n123774# m1_1634_n2388# 0.017213f
C5508 XM1/a_100_n166458# XM2/a_n100_n321571# 0.005074f
C5509 XM1/a_100_17350# XM3/a_n100_68397# 2.85e-20
C5510 XM1/a_n100_n63163# m1_1634_n2388# 1.3e-19
C5511 XM4/w_n358_n132787# XM2/a_n158_n192310# 0.103073f
C5512 XM1/a_100_27402# XM3/a_n100_79793# 3.44e-21
C5513 XM1/a_n158_n47270# XM3/a_n100_4165# 3.31e-20
C5514 XM1/a_n158_80534# XM4/w_n358_n132787# 5.68e-32
C5515 XM1/a_100_n86042# XM4/w_n358_n132787# 0.048442f
C5516 XM1/a_n100_n64599# XM4/w_n358_n132787# 0.013474f
C5517 XM1/a_n100_n37315# XM3/a_n158_13586# 2.85e-20
C5518 XM4/w_n358_n132787# XM3/a_n158_117186# 0.038462f
C5519 XM1/a_n158_n35782# XM2/a_n158_n189674# 9.28e-21
C5520 XM3/a_n100_25921# XM4/a_n100_25921# 0.009521f
C5521 XM2/a_100_n234486# XM3/a_n158_n29926# 0.054548f
C5522 XM4/w_n358_n132787# XM4/a_n100_70469# -0.004445f
C5523 XM1/a_n100_n87575# XM3/a_n158_n37178# 1.99e-22
C5524 XM2/a_n100_n239855# XM4/a_100_n35106# 2.56e-20
C5525 XM1/a_100_n61630# XM3/a_n100_n9303# 2.23e-20
C5526 XM1/a_100_107818# XM2/a_n158_n47330# 0.082979f
C5527 XM3/a_n100_n36239# m1_1634_n2388# 0.072014f
C5528 XM1/a_100_28838# XM4/w_n358_n132787# 0.055058f
C5529 XM2/a_100_n276662# XM3/a_n100_n71463# 0.010147f
C5530 XM2/a_100_n94778# XM3/a_n158_110970# 0.077916f
C5531 XM2/a_n100_n94875# XM3/a_n100_109837# 1.4e-19
C5532 XM4/w_n358_n132787# XM3/a_n158_n108662# 0.032295f
C5533 XM4/a_n100_n95291# m1_1634_n2388# 0.072015f
C5534 XM1/a_100_79098# XM2/a_n100_n76423# 0.005074f
C5535 XM1/a_n100_67513# XM3/a_n158_119258# 1.49e-20
C5536 XM1/a_n100_n90447# XM3/a_n158_n39250# 2.85e-20
C5537 XM1/a_n100_n80395# XM2/a_n158_n234486# 0.010147f
C5538 XM1/a_n158_64738# XM3/a_n100_116053# 3.89e-20
C5539 XM4/w_n358_n132787# XM3/a_n100_94297# 0.008928f
C5540 XM1/a_n100_n77523# XM2/a_100_n231850# 1.45e-19
C5541 XM1/a_n100_n44495# XM3/a_n158_6334# 2.85e-20
C5542 XM1/a_n158_25966# XM2/a_n100_n126507# 5.46e-20
C5543 XM4/w_n358_n132787# XM2/a_100_n129046# 0.103342f
C5544 XM2/a_n158_n313566# XM3/a_n100_n106687# 7.26e-20
C5545 XM1/a_n100_n116295# XM2/a_100_n271390# 7.26e-20
C5546 XM2/a_100_n247666# m1_1634_n2388# 0.019664f
C5547 XM4/w_n358_n132787# XM3/a_n100_39389# 0.009186f
C5548 XM4/a_100_104754# m1_1634_n2388# 6.1e-20
C5549 XM1/a_n158_n182254# XM2/a_n158_n337290# 4.64e-21
C5550 XM2/a_100_n110594# XM3/a_n100_94297# 0.010147f
C5551 XM1/a_100_n170766# XM2/a_100_n326746# 4.64e-21
C5552 XM4/w_n358_n132787# XM2/a_n158_n316202# 0.107093f
C5553 XM4/w_n358_n132787# XM4/a_n100_31101# -0.004445f
C5554 XM1/a_n100_n74651# XM3/a_n158_n23710# 2.85e-20
C5555 XM1/a_n100_89053# XM2/a_100_n65782# 7.26e-20
C5556 XM3/a_n100_n75607# m1_1634_n2388# 0.072015f
C5557 XM1/a_100_n38654# XM2/a_n158_n192310# 0.116862f
C5558 XM2/a_100_n152770# XM3/a_n100_51821# 0.005074f
C5559 XM1/a_n100_51717# XM4/w_n358_n132787# 0.01363f
C5560 XM1/a_n158_132230# XM2/a_n158_n23606# 4.64e-21
C5561 XM3/a_n100_n19663# XM4/a_n100_n19663# 0.009521f
C5562 XM1/a_100_66174# XM4/w_n358_n132787# 0.054609f
C5563 XM2/a_100_n194946# XM3/a_n100_9345# 0.005074f
C5564 XM1/a_n100_n27263# XM2/a_100_n181766# 1.45e-19
C5565 XM2/a_n158_n23606# XM4/w_n358_n132787# 0.107093f
C5566 XM1/a_n158_n86042# XM3/a_n100_n35203# 1.94e-20
C5567 XM1/a_100_n57322# XM2/a_n158_n210762# 0.101283f
C5568 XM2/a_n158_n13062# XM1/a_n158_142282# 4.64e-21
C5569 XM2/a_n100_n13159# XM1/a_100_139410# 0.005074f
C5570 XM1/a_n100_n166555# XM2/a_n158_n321474# 0.005074f
C5571 XM1/a_n100_n27263# XM3/a_n100_23849# 5.85e-20
C5572 XM2/a_n100_n150231# XM3/a_n158_57098# 0.004433f
C5573 XM2/a_100_n258210# XM3/a_n100_n53851# 0.005074f
C5574 XM4/a_100_n132490# m1_1634_n2388# 3.05e-20
C5575 XM1/a_n100_n91883# m1_1634_n2388# 8.78e-20
C5576 XM4/w_n358_n132787# XM4/a_n100_n40383# -0.004445f
C5577 XM1/a_n100_160853# XM2/a_n158_5390# 0.005074f
C5578 XM3/a_n158_n11278# m1_1634_n2388# 6.1e-20
C5579 XM1/a_n100_14381# XM4/w_n358_n132787# 0.01363f
C5580 XM2/a_n100_n192407# XM3/a_n158_14622# 0.005074f
C5581 XM3/a_n100_77721# m1_1634_n2388# 0.072015f
C5582 XM4/a_100_65386# m1_1634_n2388# 6.1e-20
C5583 XM1/a_100_n144918# XM3/a_n100_n93219# 9.08e-19
C5584 XM1/a_n100_n124911# XM2/a_100_n279298# 1.45e-19
C5585 XM2/a_n100_n187135# m1_1634_n2388# 0.002354f
C5586 XM1/a_n100_n15775# XM2/a_n158_n171222# 0.005074f
C5587 XM1/a_n100_n64599# XM3/a_n158_n13350# 1.49e-20
C5588 XM1/a_100_n55886# XM3/a_n100_n4123# 2.85e-20
C5589 XM1/a_100_n32910# XM3/a_n100_18669# 2.85e-20
C5590 XM3/a_n100_22813# m1_1634_n2388# 0.072015f
C5591 XM1/a_n158_69046# XM2/a_n158_n86870# 4.64e-21
C5592 XM3/a_n100_n114975# m1_1634_n2388# 0.072015f
C5593 XM4/w_n358_n132787# XM2/a_100_n252938# 0.103341f
C5594 XM2/a_n100_n108055# XM4/a_100_96466# 2.56e-20
C5595 XM1/a_n100_150801# XM2/a_n100_n5251# 0.001959f
C5596 XM1/a_n158_1554# XM2/a_n158_n152770# 9.28e-21
C5597 XM3/a_n100_119161# m1_1634_n2388# 0.072014f
C5598 XM1/a_n158_n160714# XM3/a_n100_n108759# 1.94e-20
C5599 XM2/a_n158_n295114# XM3/a_n100_n89075# 1.45e-19
C5600 XM2/a_100_n139590# XM3/a_n100_66325# 0.010147f
C5601 XM4/w_n358_n132787# XM3/a_n158_64350# 0.03704f
C5602 XM3/a_n100_n39347# XM4/a_n100_n39347# 0.009521f
C5603 XM1/a_100_87714# XM4/w_n358_n132787# 0.050354f
C5604 XM1/a_n100_168033# XM4/w_n358_n132787# 0.012765f
C5605 XM4/a_n100_128485# m1_1634_n2388# 0.072015f
C5606 XM1/a_n158_n129122# XM3/a_n100_n77679# 3.15e-20
C5607 XM1/a_n100_n100499# XM3/a_n158_n49610# 2.85e-20
C5608 XM1/a_n158_n98966# XM3/a_n100_n46599# 6.61e-21
C5609 XM1/a_n100_n12903# XM2/a_n158_n165950# 0.005074f
C5610 XM1/a_n100_n2851# XM2/a_n158_n155406# 0.005074f
C5611 XM1/a_100_43198# XM2/a_n158_n110594# 0.116862f
C5612 XM4/w_n358_n132787# XM3/a_n100_n20699# 0.008937f
C5613 XM4/a_100_n6098# m1_1634_n2388# 6.1e-20
C5614 XM2/a_100_n181766# XM3/a_n100_23849# 0.010147f
C5615 XM2/a_n158_23842# XM4/w_n358_n132787# 0.107093f
C5616 XM4/w_n358_n132787# XM4/a_n100_1057# -0.004445f
C5617 XM4/w_n358_n132787# XM3/a_n158_9442# 0.038652f
C5618 XM4/w_n358_n132787# XM4/a_n100_n79751# -0.004445f
C5619 XM1/a_n100_n110551# XM2/a_100_n263482# 7.26e-20
C5620 XM1/a_100_159514# XM2/a_n158_5390# 0.116862f
C5621 XM1/a_n100_n129219# XM2/a_n158_n281934# 0.005074f
C5622 XM3/a_n158_n50646# m1_1634_n2388# 6.1e-20
C5623 XM1/a_100_n2754# XM2/a_n158_n158042# 0.069347f
C5624 XM2/a_n100_n289939# XM3/a_n158_n82762# 0.005074f
C5625 XM4/a_100_26018# m1_1634_n2388# 6.1e-20
C5626 XM1/a_100_n100402# XM2/a_n100_n255671# 0.005074f
C5627 XM1/a_100_n116198# XM2/a_n100_n268851# 0.005074f
C5628 XM3/a_n100_78757# XM4/a_n100_78757# 0.009521f
C5629 XM1/a_n158_n83170# XM3/a_n100_n31059# 1.94e-20
C5630 XM1/a_n100_n44495# XM2/a_100_n200218# 7.26e-20
C5631 XM4/w_n358_n132787# XM2/a_n100_n192407# 0.027332f
C5632 XM2/a_n158_n10426# XM1/a_100_142282# 0.030012f
C5633 XM2/a_n100_n311027# m1_1634_n2388# 0.001347f
C5634 XM1/a_n158_n113326# XM2/a_n158_n266118# 4.64e-21
C5635 XM2/a_n158_26478# XM1/a_100_179618# 0.072074f
C5636 XM1/a_n100_103413# XM2/a_100_n49966# 7.26e-20
C5637 XM3/a_n100_n59031# XM4/a_n100_n59031# 0.009521f
C5638 XM1/a_100_n4190# XM4/w_n358_n132787# 0.048442f
C5639 XM2/a_100_n324110# XM3/a_n158_n117986# 0.077916f
C5640 XM1/a_n100_n73215# XM4/w_n358_n132787# 0.012251f
C5641 XM4/a_n100_89117# m1_1634_n2388# 0.072015f
C5642 XM1/a_n158_10170# XM3/a_n100_61145# 1.94e-20
C5643 XM4/w_n358_n132787# XM3/a_n100_117089# 0.009033f
C5644 XM1/a_100_48942# XM3/a_n100_100513# 2.85e-20
C5645 XM4/w_n358_n132787# XM3/a_n100_n60067# 0.009186f
C5646 XM4/a_100_n45466# m1_1634_n2388# 6.1e-20
C5647 XM3/a_n158_47774# m1_1634_n2388# 6.1e-20
C5648 XM2/a_n158_n234486# XM3/a_n158_n29926# 4.64e-21
C5649 XM2/a_100_n168586# XM3/a_n100_38353# 0.005074f
C5650 XM4/w_n358_n132787# XM4/a_n100_n119119# -0.004445f
C5651 XM3/a_n158_n90014# m1_1634_n2388# 6.1e-20
C5652 XM2/a_n158_n276662# XM3/a_n100_n71463# 1.45e-19
C5653 XM1/a_n158_n9934# XM3/a_n100_41461# 3.39e-20
C5654 XM1/a_n100_n182351# m1_1634_n2388# 1.3e-19
C5655 XM2/a_100_n94778# XM3/a_n100_110873# 0.010147f
C5656 XM2/a_100_n231850# XM3/a_n158_n24746# 0.00937f
C5657 XM1/a_n100_163725# XM2/a_100_10662# 7.26e-20
C5658 XM1/a_n100_68949# XM4/w_n358_n132787# 0.013474f
C5659 XM2/a_n100_n237219# XM4/a_100_n29926# 2.56e-20
C5660 XM1/a_n100_67513# XM3/a_n100_119161# 6.37e-19
C5661 XM1/a_100_63302# XM3/a_n158_115114# 0.003891f
C5662 XM1/a_n158_n101838# XM3/a_n100_n50743# 1.94e-20
C5663 XM1/a_100_100638# XM2/a_100_n52602# 4.64e-21
C5664 XM1/a_n100_n77523# XM2/a_n158_n231850# 0.010147f
C5665 XM3/a_n100_n78715# XM4/a_n100_n78715# 0.009521f
C5666 XM1/a_n100_n116295# XM2/a_n158_n271390# 0.005074f
C5667 XM4/w_n358_n132787# XM2/a_n158_n129046# 0.101988f
C5668 XM1/a_n100_22997# XM4/w_n358_n132787# 0.012874f
C5669 XM4/a_n100_49749# m1_1634_n2388# 0.072015f
C5670 XM1/a_100_n87478# XM2/a_100_n242394# 4.64e-21
C5671 XM1/a_n158_63302# XM2/a_n158_n89506# 4.64e-21
C5672 XM1/a_n158_n182254# XM2/a_n100_n337387# 7.26e-20
C5673 XM4/w_n358_n132787# XM3/a_n100_n99435# 0.008977f
C5674 XM4/a_100_n84834# m1_1634_n2388# 6.1e-20
C5675 XM2/a_n158_n110594# XM3/a_n100_94297# 1.45e-19
C5676 XM1/a_100_n170766# XM2/a_n158_n326746# 0.00197f
C5677 XM4/w_n358_n132787# XM2/a_n100_n316299# 0.025738f
C5678 XM1/a_n100_n87575# XM2/a_n100_n239855# 0.005487f
C5679 XM1/a_n158_n176510# XM3/a_n100_n124299# 1.94e-20
C5680 XM2/a_100_n200218# XM3/a_n158_5298# 0.077916f
C5681 XM2/a_n100_n39519# XM4/w_n358_n132787# 0.012279f
C5682 XM3/a_n158_n129382# m1_1634_n2388# 6.1e-20
C5683 XM1/a_n158_n150662# XM3/a_n100_n99435# 3.55e-20
C5684 XM1/a_100_n106146# XM3/a_n100_n55923# 5.8e-21
C5685 XM1/a_100_n60194# XM3/a_n100_n8267# 2.85e-20
C5686 XM2/a_n100_n205587# XM4/a_100_n918# 2.56e-20
C5687 XM2/a_n158_n152770# XM3/a_n100_51821# 7.26e-20
C5688 XM1/a_n100_n34443# m1_1634_n2388# 1.3e-19
C5689 XM2/a_100_n305658# XM3/a_n158_n100374# 0.077916f
C5690 XM2/a_100_n105322# XM3/a_n158_99574# 0.077916f
C5691 XM2/a_100_n76326# XM3/a_n158_128582# 0.077916f
C5692 XM2/a_n100_n76423# XM3/a_n100_127449# 0.005177f
C5693 XM1/a_n158_18786# XM2/a_n158_n136954# 4.64e-21
C5694 XM2/a_n158_n194946# XM3/a_n100_9345# 7.26e-20
C5695 XM1/a_n100_n27263# XM2/a_n158_n181766# 0.010147f
C5696 XM1/a_n100_157981# XM2/a_100_5390# 7.26e-20
C5697 XM1/a_100_n57322# XM2/a_n100_n210859# 0.005074f
C5698 XM4/w_n358_n132787# XM3/a_n158_n35106# 0.037323f
C5699 XM4/a_n100_n21735# m1_1634_n2388# 0.072014f
C5700 XM4/a_100_7370# m1_1634_n2388# 6.1e-20
C5701 XM2/a_100_n147498# XM3/a_n158_57098# 0.058053f
C5702 XM2/a_n158_n258210# XM3/a_n100_n53851# 7.26e-20
C5703 XM1/a_n100_n123475# XM3/a_n158_n72402# 2.85e-20
C5704 XM1/a_n158_n106146# XM3/a_n100_n55923# 3.41e-21
C5705 XM1/a_n100_n78959# XM3/a_n158_n27854# 2.85e-20
C5706 XM1/a_n100_45973# XM3/a_n158_96466# 2.82e-20
C5707 XM3/a_n100_n98399# XM4/a_n100_n98399# 0.009521f
C5708 XM1/a_n100_n84703# XM2/a_100_n237122# 7.26e-20
C5709 XM4/a_n100_10381# m1_1634_n2388# 0.072015f
C5710 XM2/a_100_n189674# XM3/a_n158_14622# 0.028843f
C5711 XM1/a_n100_124953# XM2/a_100_n28878# 1.45e-19
C5712 XM1/a_n100_71821# XM2/a_n100_n84331# 0.002666f
C5713 XM2/a_100_n213398# XM3/a_n158_n7134# 0.077916f
C5714 XM4/a_100_n124202# m1_1634_n2388# 6.1e-20
C5715 XM1/a_n100_n134963# XM2/a_100_n287206# 3.17e-20
C5716 XM1/a_n100_n124911# XM2/a_n158_n279298# 0.010147f
C5717 XM2/a_100_n184402# m1_1634_n2388# 0.021879f
C5718 XM1/a_100_120742# XM2/a_100_n34150# 4.64e-21
C5719 XM4/w_n358_n132787# XM3/a_n100_58037# 0.009186f
C5720 XM2/a_100_n255574# XM3/a_n100_n48671# 0.005074f
C5721 XM1/a_n158_n42962# XM3/a_n100_9345# 1.86e-20
C5722 XM1/a_n100_160853# XM4/w_n358_n132787# 0.012279f
C5723 XM1/a_n158_69046# XM2/a_n100_n86967# 7.26e-20
C5724 XM4/w_n358_n132787# XM2/a_n158_n252938# 0.107093f
C5725 XM1/a_n158_n71682# XM3/a_n158_n19566# 1.14e-21
C5726 XM2/a_n100_7929# XM4/w_n358_n132787# 0.012279f
C5727 XM4/w_n358_n132787# XM1/a_100_142282# 0.053546f
C5728 XM1/a_n100_76129# m1_1634_n2388# 9.25e-20
C5729 XM1/a_n100_n156503# XM3/a_n158_n105554# 2.85e-20
C5730 XM1/a_n100_n76087# m1_1634_n2388# 9.07e-20
C5731 XM1/a_n100_n25827# XM3/a_n158_24982# 1.61e-19
C5732 XM4/w_n358_n132787# XM4/a_n100_104657# -0.004445f
C5733 XM4/w_n358_n132787# XM1/a_n100_n167991# 0.012864f
C5734 XM2/a_n158_n139590# XM3/a_n100_66325# 1.45e-19
C5735 XM1/a_100_n12806# XM2/a_100_n168586# 4.64e-21
C5736 XM1/a_n100_116337# XM4/w_n358_n132787# 0.012279f
C5737 XM1/a_100_n110454# XM4/w_n358_n132787# 0.054609f
C5738 XM1/a_n100_33049# XM3/a_n158_84034# 2.85e-20
C5739 XM2/a_n100_n105419# XM4/a_100_101646# 2.56e-20
C5740 XM4/w_n358_n132787# XM3/a_n158_n74474# 0.032295f
C5741 XM4/a_n100_n61103# m1_1634_n2388# 0.072015f
C5742 XM2/a_n158_n181766# XM3/a_n100_23849# 1.45e-19
C5743 XM3/a_n100_46641# XM4/a_n100_46641# 0.009521f
C5744 XM1/a_100_24530# m1_1634_n2388# 4.87e-19
C5745 XM1/a_n100_n110551# XM2/a_n158_n263482# 0.005074f
C5746 XM2/a_100_n134318# XM3/a_n158_71602# 0.077916f
C5747 XM3/a_n100_n118083# XM4/a_n100_n118083# 0.009521f
C5748 XM1/a_100_n2754# XM2/a_n100_n158139# 0.005074f
C5749 XM2/a_n100_n292575# XM4/a_100_n87942# 2.56e-20
C5750 XM2/a_100_n287206# XM3/a_n158_n82762# 0.043253f
C5751 XM1/a_n158_n45834# XM3/a_n100_5201# 1.94e-20
C5752 XM1/a_n100_79001# XM3/a_n158_129618# 2.85e-20
C5753 XM1/a_100_n100402# XM2/a_100_n252938# 4.64e-21
C5754 XM3/a_n100_96369# m1_1634_n2388# 0.072015f
C5755 XM2/a_100_n329382# XM3/a_n100_n124299# 0.010147f
C5756 XM2/a_100_n176494# XM3/a_n158_29126# 0.077916f
C5757 XM1/a_n100_113465# XM2/a_100_n42058# 7.26e-20
C5758 XM4/a_n100_n132587# XM4/w_n358_n132787# -3.9e-19
C5759 XM1/a_100_159514# XM4/w_n358_n132787# 0.048442f
C5760 XM2/a_n100_n123871# m1_1634_n2388# 7.61e-19
C5761 XM1/a_n158_25966# XM3/a_n100_77721# 1.94e-20
C5762 XM1/a_n100_n44495# XM2/a_n158_n200218# 0.005074f
C5763 XM3/a_n100_41461# m1_1634_n2388# 0.072015f
C5764 XM4/w_n358_n132787# XM2/a_100_n189674# 0.103667f
C5765 XM4/w_n358_n132787# XM4/a_n100_65289# -0.004445f
C5766 XM2/a_100_n308294# m1_1634_n2388# 0.017936f
C5767 XM1/a_n158_n113326# XM2/a_n100_n266215# 7.26e-20
C5768 XM1/a_n158_n64502# XM3/a_n100_n12411# 1.94e-20
C5769 XM1/a_n100_n50239# XM2/a_100_n205490# 7.26e-20
C5770 XM3/a_n100_n41419# m1_1634_n2388# 0.072015f
C5771 XM4/w_n358_n132787# XM3/a_n158_82998# 0.038462f
C5772 XM2/a_100_n237122# XM3/a_n100_n31059# 0.010147f
C5773 XM4/w_n358_n132787# XM3/a_n158_n113842# 0.032295f
C5774 XM4/a_n100_n100471# m1_1634_n2388# 0.072015f
C5775 XM2/a_n100_n234583# XM3/a_n158_n29926# 0.005074f
C5776 XM4/w_n358_n132787# XM3/a_n158_n2990# 0.032295f
C5777 XM1/a_n158_n77426# XM3/a_n100_n26915# 1.94e-20
C5778 XM4/w_n358_n132787# XM3/a_n158_28090# 0.038311f
C5779 XM2/a_n158_n168586# XM3/a_n100_38353# 7.26e-20
C5780 XM1/a_100_n107582# XM3/a_n100_n55923# 2.85e-20
C5781 XM2/a_n158_n94778# XM3/a_n100_110873# 1.45e-19
C5782 XM4/w_n358_n132787# XM4/a_n100_n6195# -0.004445f
C5783 XM2/a_n158_n231850# XM3/a_n158_n24746# 4.64e-21
C5784 XM1/a_100_n37218# XM2/a_100_n192310# 4.64e-21
C5785 XM2/a_100_n163314# XM3/a_n158_43630# 0.024949f
C5786 XM1/a_100_63302# XM3/a_n100_115017# 6.54e-19
C5787 XM4/a_100_99574# m1_1634_n2388# 6.1e-20
C5788 XM1/a_100_n31474# XM2/a_100_n187038# 4.64e-21
C5789 XM1/a_100_69046# XM3/a_n100_121233# 2.85e-20
C5790 XM4/w_n358_n132787# XM4/a_n100_25921# -0.004445f
C5791 XM3/a_n100_n80787# m1_1634_n2388# 0.072015f
C5792 XM4/w_n358_n132787# XM2/a_n100_n129143# 0.023764f
C5793 XM2/a_100_n310930# XM3/a_n100_n106687# 0.005074f
C5794 XM2/a_n100_n247763# m1_1634_n2388# 0.003351f
C5795 XM1/a_100_n87478# XM2/a_n158_n242394# 0.105567f
C5796 XM1/a_n158_63302# XM2/a_n100_n89603# 7.26e-20
C5797 XM1/a_100_n170766# XM2/a_n100_n326843# 0.005074f
C5798 XM4/w_n358_n132787# XM2/a_100_n313566# 0.104499f
C5799 XM1/a_100_n124814# XM3/a_n100_n74571# 1.17e-20
C5800 XM1/a_100_163822# XM2/a_n100_10565# 0.005074f
C5801 XM3/a_n158_66422# m1_1634_n2388# 6.1e-20
C5802 XM1/a_n100_n84703# XM3/a_n100_n33131# 7.68e-19
C5803 XM1/a_n158_n130558# XM3/a_n100_n78715# 1.94e-20
C5804 XM1/a_n100_n74651# XM2/a_100_n229214# 1.45e-19
C5805 XM2/a_n100_n160775# XM4/a_100_43630# 2.56e-20
C5806 XM1/a_n100_165161# XM2/a_n158_10662# 0.010147f
C5807 XM1/a_n100_60333# XM2/a_100_n94778# 7.26e-20
C5808 XM1/a_100_n146354# XM4/w_n358_n132787# 0.048442f
C5809 XM4/w_n358_n132787# XM4/a_n100_n45563# -0.004445f
C5810 XM3/a_n158_11514# m1_1634_n2388# 6.1e-20
C5811 XM3/a_n158_n16458# m1_1634_n2388# 6.1e-20
C5812 XM2/a_100_n218670# XM3/a_n100_n13447# 0.010147f
C5813 XM1/a_n100_119209# XM4/w_n358_n132787# 0.011718f
C5814 XM1/a_n100_90489# XM2/a_100_n63146# 1.45e-19
C5815 XM2/a_100_n76326# XM3/a_n100_128485# 0.010147f
C5816 XM1/a_n158_18786# XM2/a_n100_n137051# 7.26e-20
C5817 XM4/a_100_60206# m1_1634_n2388# 6.1e-20
C5818 XM1/a_n100_n166555# XM2/a_100_n318838# 5.76e-20
C5819 XM2/a_n158_n147498# XM3/a_n158_57098# 4.64e-21
C5820 XM3/a_n100_n120155# m1_1634_n2388# 0.072015f
C5821 XM1/a_n100_n84703# XM2/a_n158_n237122# 0.005074f
C5822 XM2/a_n158_n189674# XM3/a_n158_14622# 4.64e-21
C5823 XM4/w_n358_n132787# XM1/a_n100_136441# 0.013155f
C5824 XM1/a_n100_71821# XM2/a_100_n81598# 7.26e-20
C5825 XM1/a_n100_n134963# XM2/a_n158_n287206# 0.002589f
C5826 XM2/a_n158_n184402# m1_1634_n2388# 2.36e-21
C5827 XM1/a_100_61866# XM4/w_n358_n132787# 0.048442f
C5828 XM1/a_100_n142046# XM3/a_n158_n91050# 0.00544f
C5829 XM2/a_n158_n255574# XM3/a_n100_n48671# 7.26e-20
C5830 XM1/a_n100_n15775# XM2/a_100_n168586# 7.26e-20
C5831 XM1/a_n100_n103371# XM4/w_n358_n132787# 0.012508f
C5832 XM3/a_n100_14525# XM4/a_n100_14525# 0.009521f
C5833 XM4/a_n100_123305# m1_1634_n2388# 0.072015f
C5834 XM3/a_n100_99477# XM4/a_n100_99477# 0.009521f
C5835 XM1/a_n100_35921# XM3/a_n158_87142# 2.32e-20
C5836 XM4/w_n358_n132787# XM2/a_n100_n253035# 0.024857f
C5837 XM4/w_n358_n132787# XM3/a_n100_n25879# 0.009017f
C5838 XM4/a_100_n11278# m1_1634_n2388# 6.1e-20
C5839 XM1/a_n100_n48803# XM3/a_n158_3226# 2.85e-20
C5840 XM3/a_n100_116053# XM4/a_n100_116053# 0.009521f
C5841 XM4/w_n358_n132787# XM3/a_n100_3129# 0.009186f
C5842 XM3/a_n158_120294# m1_1634_n2388# 6.1e-20
C5843 XM4/w_n358_n132787# XM4/a_n100_n84931# -0.004445f
C5844 XM1/a_n100_n134963# XM3/a_n158_n83798# 2.85e-20
C5845 XM3/a_n158_n55826# m1_1634_n2388# 6.1e-20
C5846 XM1/a_100_n12806# XM2/a_n158_n168586# 0.021444f
C5847 XM1/a_n100_63205# m1_1634_n2388# 1.3e-19
C5848 XM4/a_100_20838# m1_1634_n2388# 6.1e-20
C5849 XM1/a_100_n83170# XM3/a_n100_n32095# 2.85e-20
C5850 XM1/a_100_n75990# XM2/a_100_n231850# 4.64e-21
C5851 XM1/a_n100_120645# XM2/a_100_n34150# 7.26e-20
C5852 XM1/a_100_31710# XM3/a_n100_82901# 5.52e-20
C5853 XM1/a_n100_n40187# XM3/a_n158_11514# 7.95e-22
C5854 XM1/a_n100_n24391# XM3/a_n100_25921# 0.001145f
C5855 XM1/a_n100_116337# XM2/a_100_n39422# 7.26e-20
C5856 XM1/a_n100_n170863# XM2/a_100_n326746# 7.26e-20
C5857 XM1/a_n100_n107679# XM4/w_n358_n132787# 0.01363f
C5858 XM2/a_n158_n287206# XM3/a_n158_n82762# 4.64e-21
C5859 XM1/a_100_n2754# XM2/a_100_n155406# 4.64e-21
C5860 XM4/w_n358_n132787# XM1/a_n100_176649# 0.012279f
C5861 XM1/a_100_n100402# XM2/a_n158_n252938# 0.013265f
C5862 XM1/a_100_n34346# XM3/a_n158_17730# 0.001211f
C5863 XM1/a_100_36018# XM2/a_n158_n118502# 0.116862f
C5864 XM2/a_n158_n329382# XM3/a_n100_n124299# 1.45e-19
C5865 XM1/a_n100_n147887# XM3/a_n100_n96327# 6.76e-19
C5866 XM4/w_n358_n132787# XM4/a_n100_7273# -0.004445f
C5867 XM1/a_n100_n43059# XM3/a_n100_9345# 5.2e-20
C5868 XM1/a_n100_n147887# XM2/a_100_n303022# 7.26e-20
C5869 XM1/a_n100_n11467# XM3/a_n158_40522# 2.85e-20
C5870 XM2/a_100_n121138# m1_1634_n2388# 0.023369f
C5871 XM4/a_n100_83937# m1_1634_n2388# 0.072015f
C5872 XM4/w_n358_n132787# XM3/a_n100_76685# 0.009186f
C5873 XM1/a_100_n166458# XM2/a_n100_n318935# 0.004675f
C5874 XM2/a_100_n284570# XM3/a_n158_n77582# 0.020665f
C5875 sw_bn iout_n 0.046619f
C5876 XM2/a_n100_n289939# XM4/a_100_n82762# 2.56e-20
C5877 XM4/w_n358_n132787# XM3/a_n100_n65247# 0.008918f
C5878 XM4/a_100_n50646# m1_1634_n2388# 6.1e-20
C5879 XM4/w_n358_n132787# XM2/a_n158_n189674# 0.107093f
C5880 XM4/w_n358_n132787# XM4/a_n100_n124299# -0.004445f
C5881 XM2/a_n158_n308294# m1_1634_n2388# 2.36e-21
C5882 XM1/a_n100_n50239# XM2/a_n158_n205490# 0.005074f
C5883 XM4/w_n358_n132787# XM3/a_n100_21777# 0.009186f
C5884 XM3/a_n158_n95194# m1_1634_n2388# 6.1e-20
C5885 XM1/a_n100_160853# XM2/a_100_8026# 7.26e-20
C5886 XM2/a_n100_n126507# XM3/a_n100_80829# 0.00499f
C5887 XM2/a_n158_n237122# XM3/a_n100_n31059# 1.45e-19
C5888 XM4/w_n358_n132787# XM3/a_n158_118222# 0.032295f
C5889 XM2/a_n158_23842# XM1/a_n158_178182# 9.28e-21
C5890 XM1/a_n100_166597# XM2/a_100_10662# 4.86e-20
C5891 XM1/a_n100_152237# XM4/w_n358_n132787# 0.013902f
C5892 XM1/a_n100_n117731# XM3/a_n158_n65150# 4.62e-21
C5893 XM1/a_100_n11370# XM4/w_n358_n132787# 0.048442f
C5894 XM2/a_100_n94778# XM3/a_n158_112006# 0.040527f
C5895 XM1/a_n100_n104807# m1_1634_n2388# 9.61e-20
C5896 XM1/a_n158_n68810# XM3/a_n100_n17591# 2.91e-20
C5897 XM1/a_100_n51578# XM3/a_n100_21# 2.85e-20
C5898 XM2/a_n158_n68418# XM4/w_n358_n132787# 0.1039f
C5899 XM2/a_n100_n231947# XM3/a_n158_n24746# 0.005074f
C5900 XM1/a_n158_n17114# XM3/a_n100_33173# 1.62e-20
C5901 XM1/a_n100_126389# XM4/w_n358_n132787# 0.012279f
C5902 XM1/a_n100_101977# XM2/a_n158_n52602# 0.010147f
C5903 XM1/a_100_n37218# XM2/a_n158_n192310# 0.088431f
C5904 XM2/a_n158_n163314# XM3/a_n158_43630# 4.64e-21
C5905 XM4/a_n100_44569# m1_1634_n2388# 0.072015f
C5906 XM1/a_100_n31474# XM2/a_n158_n187038# 0.042475f
C5907 XM4/w_n358_n132787# XM3/a_n100_n104615# 0.007926f
C5908 XM4/a_100_n90014# m1_1634_n2388# 6.1e-20
C5909 XM1/a_n158_64738# XM3/a_n100_117089# 9.82e-21
C5910 XM3/a_n100_60109# m1_1634_n2388# 0.072015f
C5911 XM1/a_n100_n116295# XM2/a_100_n268754# 7.26e-20
C5912 XM4/w_n358_n132787# XM2/a_100_n126410# 0.104368f
C5913 XM1/a_n158_n167894# XM2/a_n158_n321474# 4.64e-21
C5914 XM2/a_n158_n310930# XM3/a_n100_n106687# 7.26e-20
C5915 XM2/a_100_n245030# m1_1634_n2388# 0.017213f
C5916 XM1/a_100_n87478# XM2/a_n100_n242491# 0.005074f
C5917 XM1/a_n158_n182254# XM2/a_n158_n334654# 4.64e-21
C5918 XM1/a_n158_123614# XM2/a_n158_n31514# 4.64e-21
C5919 XM1/a_100_n170766# XM2/a_100_n324110# 4.64e-21
C5920 XM4/w_n358_n132787# XM2/a_n158_n313566# 0.107093f
C5921 XM2/a_100_n266118# XM3/a_n158_n59970# 0.077916f
C5922 XM1/a_n100_91925# XM4/w_n358_n132787# 0.012279f
C5923 XM1/a_n100_n183787# XM4/w_n358_n132787# 0.011821f
C5924 XM1/a_n100_n156503# m1_1634_n2388# 1.3e-19
C5925 XM1/a_100_181054# XM4/w_n358_n132787# 0.048442f
C5926 XM1/a_n158_171002# XM2/a_n100_18473# 7.26e-20
C5927 XM2/a_100_n308294# XM3/a_n100_n101507# 0.005074f
C5928 XM4/a_n100_n26915# m1_1634_n2388# 0.072015f
C5929 XM1/a_n100_93361# XM2/a_100_n60510# 1.45e-19
C5930 XM1/a_n100_n147887# m1_1634_n2388# 9.43e-20
C5931 XM4/w_n358_n132787# XM3/a_n158_n40286# 0.033682f
C5932 XM4/w_n358_n132787# XM3/a_n158_46738# 0.032893f
C5933 XM1/a_n100_1457# m1_1634_n2388# 8.14e-20
C5934 XM1/a_n100_n153631# XM3/a_n158_n102446# 2.85e-20
C5935 XM1/a_n100_n74651# XM2/a_n158_n229214# 0.010147f
C5936 XM1/a_n100_60333# XM2/a_n158_n94778# 0.005074f
C5937 XM2/a_n158_n218670# XM3/a_n100_n13447# 1.45e-19
C5938 XM2/a_n158_n76326# XM3/a_n100_128485# 1.45e-19
C5939 XM1/a_n100_123517# XM2/a_100_n28878# 7.26e-20
C5940 XM1/a_100_n87478# m1_1634_n2388# 6.08e-20
C5941 XM4/a_100_n129382# m1_1634_n2388# 6.1e-20
C5942 XM1/a_n100_n166555# XM2/a_n158_n318838# 0.004675f
C5943 XM3/a_n100_67361# XM4/a_n100_67361# 0.009521f
C5944 XM2/a_n100_n147595# XM3/a_n158_57098# 0.005074f
C5945 XM2/a_n100_n158139# XM4/a_100_48810# 2.56e-20
C5946 XM1/a_n158_84842# XM2/a_n158_n71054# 4.64e-21
C5947 XM1/a_n100_n127783# XM4/w_n358_n132787# 0.013513f
C5948 XM1/a_n100_n103371# XM3/a_n158_n52718# 2.85e-20
C5949 XM1/a_n158_129358# XM2/a_n100_n23703# 7.26e-20
C5950 XM2/a_n100_n189771# XM3/a_n158_14622# 0.005074f
C5951 XM1/a_n100_71821# XM2/a_n158_n81598# 0.005074f
C5952 XM4/w_n358_n132787# XM4/a_n100_99477# -0.004445f
C5953 XM1/a_n100_n134963# XM2/a_n100_n287303# 0.002458f
C5954 XM2/a_n100_n184499# m1_1634_n2388# 0.001625f
C5955 XM3/a_n100_n7231# m1_1634_n2388# 0.072015f
C5956 XM1/a_n100_n15775# XM2/a_n158_n168586# 0.005074f
C5957 XM1/a_n100_10073# XM4/w_n358_n132787# 0.013542f
C5958 XM1/a_n158_69046# XM2/a_n158_n84234# 4.64e-21
C5959 XM4/w_n358_n132787# XM2/a_100_n250302# 0.103711f
C5960 XM1/a_n158_163822# XM2/a_n100_10565# 7.26e-20
C5961 XM3/a_n158_85070# m1_1634_n2388# 6.1e-20
C5962 XM4/w_n358_n132787# XM3/a_n158_n79654# 0.032295f
C5963 XM4/a_n100_n66283# m1_1634_n2388# 0.072015f
C5964 XM3/a_n100_120197# m1_1634_n2388# 0.072015f
C5965 XM1/a_n100_n122039# XM3/a_n100_n70427# 0.001161f
C5966 XM1/a_100_n117634# XM3/a_n100_n67319# 2.85e-20
C5967 XM1/a_100_n12806# XM2/a_n100_n168683# 0.005074f
C5968 XM3/a_n158_30162# m1_1634_n2388# 6.1e-20
C5969 XM2/a_100_n247666# XM3/a_n158_n42358# 0.077916f
C5970 XM1/a_100_79098# XM2/a_n158_n73690# 0.037801f
C5971 XM1/a_100_n75990# XM2/a_n158_n231850# 0.013654f
C5972 XM2/a_100_n289842# XM3/a_n100_n83895# 0.010147f
C5973 XM1/a_n100_n170863# XM2/a_n158_n326746# 0.005074f
C5974 XM1/a_n100_n143579# XM3/a_n100_n93219# 5.2e-19
C5975 XM2/a_n100_n287303# XM3/a_n158_n82762# 0.005074f
C5976 XM1/a_n158_n103274# XM3/a_n100_n52815# 1.94e-20
C5977 XM1/a_100_n27166# XM3/a_n100_23849# 2.85e-20
C5978 XM1/a_100_n2754# XM2/a_n158_n155406# 0.024559f
C5979 XM1/a_100_n100402# XM2/a_n100_n253035# 0.005074f
C5980 XM1/a_n100_n17211# m1_1634_n2388# 8.14e-20
C5981 XM1/a_100_60430# XM3/a_n100_110873# 2.85e-20
C5982 XM4/w_n358_n132787# XM4/a_n100_60109# -0.004445f
C5983 XM1/a_n100_n54547# m1_1634_n2388# 5.14e-20
C5984 XM3/a_n100_n46599# m1_1634_n2388# 0.072015f
C5985 XM1/a_n100_n147887# XM2/a_n158_n303022# 0.005074f
C5986 XM2/a_n158_n121138# m1_1634_n2388# 5.91e-22
C5987 XM1/a_100_n152098# XM2/a_100_n305658# 4.64e-21
C5988 XM2/a_n158_n284570# XM3/a_n158_n77582# 4.64e-21
C5989 XM1/a_n100_n44495# XM2/a_100_n197582# 7.26e-20
C5990 XM4/w_n358_n132787# XM3/a_n158_n119022# 0.032295f
C5991 XM4/a_n100_n105651# m1_1634_n2388# 0.072015f
C5992 XM3/a_n100_n5159# XM4/a_n100_n5159# 0.009521f
C5993 XM1/a_100_17350# XM3/a_n100_69433# 2.85e-20
C5994 XM1/a_100_n169330# XM3/a_n100_n119119# 2.27e-21
C5995 XM4/w_n358_n132787# XM2/a_n100_n189771# 0.025565f
C5996 XM2/a_n100_n308391# m1_1634_n2388# 0.001429f
C5997 XM1/a_100_n104710# XM3/a_n100_n53851# 2.85e-20
C5998 XM1/a_100_n74554# XM2/a_n158_n229214# 0.116862f
C5999 XM1/a_n158_1554# XM3/a_n100_51821# 1.22e-20
C6000 XM2/a_100_n123774# XM3/a_n100_80829# 0.005074f
C6001 XM1/a_n100_n37315# XM3/a_n158_14622# 2.85e-20
C6002 XM4/w_n358_n132787# XM3/a_n100_118125# 0.009186f
C6003 XM4/w_n358_n132787# XM4/a_n100_n11375# -0.004445f
C6004 XM1/a_100_107818# XM2/a_n158_n44694# 0.010928f
C6005 XM1/a_n100_n84703# XM4/w_n358_n132787# 0.013481f
C6006 XM2/a_100_n165950# XM3/a_n100_38353# 0.005074f
C6007 XM4/a_100_94394# m1_1634_n2388# 6.1e-20
C6008 XM2/a_n100_n121235# XM3/a_n158_86106# 0.003994f
C6009 XM1/a_n100_12945# m1_1634_n2388# 9.25e-20
C6010 XM4/w_n358_n132787# XM4/a_n100_20741# -0.004445f
C6011 XM2/a_n158_n94778# XM3/a_n158_112006# 4.64e-21
C6012 XM2/a_100_n94778# XM3/a_n100_111909# 0.005074f
C6013 XM1/a_n158_n88914# XM3/a_n100_n37275# 1.94e-20
C6014 XM3/a_n100_n85967# m1_1634_n2388# 0.072015f
C6015 XM2/a_100_n229214# XM3/a_n158_n24746# 0.04559f
C6016 XM1/a_100_n44398# XM3/a_n100_7273# 2.85e-20
C6017 XM1/a_n158_30274# XM2/a_n158_n123774# 9.28e-21
C6018 XM2/a_n100_n234583# XM4/a_100_n29926# 2.56e-20
C6019 XM1/a_100_n37218# XM2/a_n100_n192407# 0.005074f
C6020 XM2/a_n100_n163411# XM3/a_n158_43630# 0.005074f
C6021 XM1/a_100_n154970# XM3/a_n158_n104518# 4.55e-19
C6022 XM2/a_100_n271390# XM3/a_n100_n66283# 0.010147f
C6023 XM1/a_100_n31474# XM2/a_n100_n187135# 0.005074f
C6024 XM3/a_n100_n24843# XM4/a_n100_n24843# 0.009521f
C6025 XM1/a_100_73354# XM4/w_n358_n132787# 0.052982f
C6026 XM4/w_n358_n132787# XM3/a_n100_95333# 0.009186f
C6027 XM1/a_100_n179382# XM3/a_n158_n127310# 0.001739f
C6028 XM1/a_n100_180957# XM4/w_n358_n132787# 0.012279f
C6029 XM1/a_n100_175213# XM4/w_n358_n132787# 0.012279f
C6030 XM1/a_100_162386# XM4/w_n358_n132787# 0.048442f
C6031 XM1/a_n100_n116295# XM2/a_n158_n268754# 0.005074f
C6032 XM1/a_100_171002# XM2/a_n158_15934# 0.090768f
C6033 XM4/w_n358_n132787# XM2/a_n158_n126410# 0.106546f
C6034 XM1/a_n158_n167894# XM2/a_n100_n321571# 1.5e-20
C6035 XM4/w_n358_n132787# XM3/a_n100_40425# 0.00985f
C6036 XM1/a_n158_73354# XM2/a_n158_n81598# 4.64e-21
C6037 XM1/a_n100_n27263# m1_1634_n2388# 1.23e-19
C6038 XM1/a_n158_n182254# XM2/a_n100_n334751# 7.26e-20
C6039 XM4/w_n358_n132787# XM4/a_n100_n50743# -0.004445f
C6040 XM1/a_100_n73118# XM3/a_n100_n21735# 5.71e-20
C6041 XM2/a_100_n110594# XM3/a_n100_95333# 0.010147f
C6042 XM1/a_100_n170766# XM2/a_n158_n324110# 0.091936f
C6043 XM4/w_n358_n132787# XM2/a_n100_n313663# 0.025024f
C6044 XM3/a_n158_n21638# m1_1634_n2388# 6.1e-20
C6045 XM3/a_n100_35245# XM4/a_n100_35245# 0.009521f
C6046 XM4/a_100_55026# m1_1634_n2388# 6.1e-20
C6047 XM1/a_n100_n180915# XM2/a_100_n334654# 1.45e-19
C6048 XM2/a_n158_n308294# XM3/a_n100_n101507# 7.26e-20
C6049 XM2/a_100_n152770# XM3/a_n100_52857# 0.010147f
C6050 XM1/a_n100_n37315# XM4/w_n358_n132787# 0.01363f
C6051 XM1/a_n158_132230# XM2/a_n158_n20970# 4.64e-21
C6052 XM1/a_n100_n86139# XM3/a_n158_n35106# 2.85e-20
C6053 XM3/a_n100_n125335# m1_1634_n2388# 0.072014f
C6054 XM2/a_100_n76326# XM3/a_n158_129618# 0.077916f
C6055 XM1/a_n158_18786# XM2/a_n158_n134318# 4.64e-21
C6056 XM2/a_100_n194946# XM3/a_n100_10381# 0.010147f
C6057 XM2/a_n158_n20970# XM4/w_n358_n132787# 0.105871f
C6058 XM2/a_n158_n10426# XM1/a_n158_142282# 4.64e-21
C6059 XM1/a_n158_92022# XM2/a_n100_n63243# 7.26e-20
C6060 XM1/a_n100_n166555# XM2/a_n100_n318935# 6.21e-19
C6061 XM3/a_n100_n44527# XM4/a_n100_n44527# 0.009521f
C6062 XM1/a_n158_175310# XM2/a_n158_21206# 9.28e-21
C6063 XM1/a_100_53250# XM2/a_100_n102686# 4.64e-21
C6064 XM1/a_n100_155109# XM4/w_n358_n132787# 0.012279f
C6065 XM4/a_n100_118125# m1_1634_n2388# 0.072015f
C6066 XM4/w_n358_n132787# XM3/a_n100_n31059# 0.009186f
C6067 XM4/a_100_n16458# m1_1634_n2388# 6.1e-20
C6068 XM3/a_n100_78757# m1_1634_n2388# 0.072015f
C6069 XM1/a_n100_71821# XM2/a_n100_n81695# 4.51e-19
C6070 XM4/w_n358_n132787# XM4/a_n100_n90111# -0.004445f
C6071 XM2/a_100_n181766# m1_1634_n2388# 0.017213f
C6072 XM3/a_n158_n61006# m1_1634_n2388# 6.1e-20
C6073 XM2/a_100_n252938# XM3/a_n100_n48671# 0.005074f
C6074 XM4/a_100_15658# m1_1634_n2388# 6.1e-20
C6075 XM3/a_n100_23849# m1_1634_n2388# 0.072015f
C6076 XM1/a_n158_69046# XM2/a_n100_n84331# 7.26e-20
C6077 XM4/w_n358_n132787# XM2/a_n158_n250302# 0.107093f
C6078 XM2/a_100_n337290# XM3/a_n158_n130418# 0.031959f
C6079 XM1/a_100_n136302# XM3/a_n158_n85870# 4.93e-19
C6080 XM1/a_100_n80298# XM3/a_n100_n27951# 1.64e-20
C6081 XM1/a_n158_n61630# XM3/a_n100_n11375# 9.82e-21
C6082 XM1/a_n100_n58855# XM3/a_n158_n8170# 2.85e-20
C6083 XM2/a_100_n139590# XM3/a_n100_67361# 0.005074f
C6084 XM4/w_n358_n132787# XM3/a_n158_65386# 0.032295f
C6085 XM1/a_100_n12806# XM2/a_100_n165950# 4.64e-21
C6086 XM2/a_n100_n102783# XM4/a_100_101646# 2.56e-20
C6087 XM1/a_n100_n45931# m1_1634_n2388# 1.1e-19
C6088 XM1/a_100_n75990# XM2/a_n100_n231947# 0.005074f
C6089 XM4/w_n358_n132787# XM3/a_n158_10478# 0.032295f
C6090 XM2/a_100_n181766# XM3/a_n100_24885# 0.005074f
C6091 XM2/a_n158_26478# XM4/w_n358_n132787# 0.106835f
C6092 XM2/a_n158_n289842# XM3/a_n100_n83895# 1.45e-19
C6093 XM3/a_n100_n64211# XM4/a_n100_n64211# 0.009521f
C6094 XM1/a_100_2990# XM4/w_n358_n132787# 0.054609f
C6095 XM1/a_n100_113465# XM4/w_n358_n132787# 0.012279f
C6096 XM1/a_100_n27166# XM2/a_n158_n181766# 0.116862f
C6097 XM4/a_n100_78757# m1_1634_n2388# 0.072015f
C6098 XM1/a_n100_n183787# XM3/a_n158_n131454# 2.85e-20
C6099 XM4/a_100_n55826# m1_1634_n2388# 6.1e-20
C6100 XM1/a_100_n2754# XM2/a_n100_n155503# 0.005074f
C6101 XM1/a_n100_58897# XM3/a_n158_109934# 2.85e-20
C6102 XM4/w_n358_n132787# XM3/a_n100_n70427# 0.008912f
C6103 XM1/a_n100_n87575# XM4/w_n358_n132787# 0.012336f
C6104 XM4/w_n358_n132787# XM4/a_n100_n129479# -0.004445f
C6105 XM1/a_n158_n166458# XM2/a_n158_n321474# 4.64e-21
C6106 XM3/a_n158_n100374# m1_1634_n2388# 6.1e-20
C6107 XM1/a_100_n68810# XM2/a_100_n223942# 4.64e-21
C6108 XM1/a_n158_n12806# XM3/a_n100_38353# 3.07e-20
C6109 XM2/a_n100_n121235# m1_1634_n2388# 0.001091f
C6110 XM1/a_100_n152098# XM2/a_n158_n305658# 0.112967f
C6111 XM2/a_n100_n284667# XM3/a_n158_n77582# 0.005074f
C6112 XM1/a_n100_n44495# XM2/a_n158_n197582# 0.005074f
C6113 XM4/w_n358_n132787# XM2/a_100_n187038# 0.103341f
C6114 XM2/a_100_n305658# m1_1634_n2388# 0.019664f
C6115 XM1/a_n100_n50239# XM2/a_100_n202854# 7.26e-20
C6116 XM1/a_n100_n24391# XM4/w_n358_n132787# 0.013882f
C6117 XM1/a_n158_n149226# XM2/a_n158_n303022# 9.28e-21
C6118 XM4/w_n358_n132787# XM3/a_n158_n6098# 0.036335f
C6119 XM1/a_n100_33049# XM2/a_100_n121138# 1.45e-19
C6120 XM1/a_n100_n114859# XM2/a_100_n268754# 1.45e-19
C6121 XM2/a_n158_n123774# XM3/a_n100_80829# 7.26e-20
C6122 XM1/a_n158_10170# XM3/a_n100_62181# 1.94e-20
C6123 XM3/a_n158_48810# m1_1634_n2388# 6.1e-20
C6124 XM3/a_n100_n83895# XM4/a_n100_n83895# 0.009521f
C6125 XM2/a_n158_n165950# XM3/a_n100_38353# 7.26e-20
C6126 XM4/a_n100_39389# m1_1634_n2388# 0.072014f
C6127 XM1/a_n100_n10031# XM3/a_n158_40522# 8.73e-20
C6128 XM1/a_n100_n5723# XM3/a_n100_44569# 7.04e-19
C6129 XM1/a_100_73354# XM3/a_n100_124341# 2.85e-20
C6130 XM2/a_100_n318838# XM3/a_n158_n112806# 0.077916f
C6131 XM4/w_n358_n132787# XM3/a_n100_n109795# 0.008335f
C6132 XM4/a_100_n95194# m1_1634_n2388# 6.1e-20
C6133 XM2/a_100_n118502# XM3/a_n158_86106# 0.059221f
C6134 XM2/a_n100_n94875# XM3/a_n158_112006# 0.005074f
C6135 XM2/a_n158_n94778# XM3/a_n100_111909# 7.26e-20
C6136 XM1/a_n158_n173638# XM3/a_n100_n122227# 2.75e-20
C6137 XM1/a_n158_n109018# XM3/a_n100_n56959# 1.94e-20
C6138 XM2/a_n158_n229214# XM3/a_n158_n24746# 4.64e-21
C6139 XM4/w_n358_n132787# XM3/a_n158_4262# 0.038462f
C6140 XM1/a_100_n37218# XM2/a_100_n189674# 4.64e-21
C6141 XM2/a_100_n160678# XM3/a_n158_43630# 0.030012f
C6142 XM1/a_n100_n175171# m1_1634_n2388# 1.3e-19
C6143 XM2/a_n158_n271390# XM3/a_n100_n66283# 1.45e-19
C6144 XM1/a_100_n31474# XM2/a_100_n184402# 4.64e-21
C6145 XM4/w_n358_n132787# XM1/a_100_n139174# 0.054609f
C6146 XM3/a_n100_88081# XM4/a_n100_88081# 0.009521f
C6147 XM1/a_100_n15678# XM4/w_n358_n132787# 0.054697f
C6148 XM1/a_n158_n114762# XM2/a_n158_n268754# 9.28e-21
C6149 XM4/w_n358_n132787# XM3/a_n158_n45466# 0.032295f
C6150 XM4/a_n100_n32095# m1_1634_n2388# 0.072015f
C6151 XM2/a_100_n226578# XM3/a_n158_n19566# 0.018328f
C6152 XM4/w_n358_n132787# XM2/a_n100_n126507# 0.024496f
C6153 XM1/a_n158_n162150# XM2/a_n158_n316202# 9.28e-21
C6154 XM2/a_n100_n245127# m1_1634_n2388# 0.002404f
C6155 XM2/a_n100_n231947# XM4/a_100_n24746# 2.56e-20
C6156 XM1/a_n158_73354# XM2/a_n100_n81695# 7.26e-20
C6157 XM1/a_n100_5765# m1_1634_n2388# 8.6e-20
C6158 XM4/w_n358_n132787# XM1/a_100_n130558# 0.048442f
C6159 XM1/a_n158_n117634# XM3/a_n100_n65247# 2.6e-21
C6160 XM1/a_n100_n81831# XM3/a_n158_n30962# 2.85e-20
C6161 XM2/a_n158_n110594# XM3/a_n100_95333# 1.45e-19
C6162 XM1/a_100_n170766# XM2/a_n100_n324207# 0.005074f
C6163 XM4/w_n358_n132787# XM2/a_100_n310930# 0.103342f
C6164 XM3/a_n100_n103579# XM4/a_n100_n103579# 0.009521f
C6165 XM2/a_n100_n36883# XM4/w_n358_n132787# 0.011718f
C6166 XM1/a_n100_n180915# XM2/a_n158_n334654# 0.010147f
C6167 XM2/a_n158_n152770# XM3/a_n100_52857# 1.45e-19
C6168 XM1/a_n100_60333# XM2/a_100_n92142# 7.26e-20
C6169 XM1/a_100_n28602# XM3/a_n158_22910# 0.002948f
C6170 XM2/a_100_n76326# XM3/a_n100_129521# 0.010147f
C6171 XM1/a_n158_18786# XM2/a_n100_n134415# 7.26e-20
C6172 XM2/a_n158_n194946# XM3/a_n100_10381# 1.45e-19
C6173 XM4/w_n358_n132787# XM4/a_n100_94297# -0.004445f
C6174 XM2/a_100_n147498# XM3/a_n158_58134# 0.077916f
C6175 XM2/a_100_n300386# XM3/a_n158_n95194# 0.077916f
C6176 XM3/a_n100_n12411# m1_1634_n2388# 0.072014f
C6177 XM1/a_100_53250# XM2/a_n158_n102686# 0.006254f
C6178 XM1/a_n100_179521# XM2/a_100_23842# 7.26e-20
C6179 XM1/a_n100_n179479# XM2/a_100_n334654# 7.26e-20
C6180 XM4/a_n100_n71463# m1_1634_n2388# 0.072015f
C6181 XM4/w_n358_n132787# XM3/a_n158_n84834# 0.032295f
C6182 XM2/a_100_n189674# XM3/a_n158_15658# 0.077916f
C6183 XM1/a_n158_n15678# XM2/a_n158_n171222# 4.64e-21
C6184 XM1/a_100_48942# XM2/a_n158_n105322# 0.116862f
C6185 XM1/a_n158_5862# XM2/a_n158_n150134# 4.64e-21
C6186 XM4/w_n358_n132787# XM3/a_n100_59073# 0.009186f
C6187 XM3/a_n100_n123263# XM4/a_n100_n123263# 0.009521f
C6188 XM2/a_n158_n252938# XM3/a_n100_n48671# 7.26e-20
C6189 XM4/w_n358_n132787# XM2/a_n100_n250399# 0.025351f
C6190 XM1/a_100_1554# XM2/a_n158_n152770# 0.116862f
C6191 XM1/a_n100_n25827# XM3/a_n158_26018# 2.85e-20
C6192 XM2/a_n100_10565# XM4/w_n358_n132787# 0.011792f
C6193 XM3/a_n158_121330# m1_1634_n2388# 6.1e-20
C6194 XM2/a_n158_n337290# XM3/a_n158_n130418# 4.64e-21
C6195 XM4/w_n358_n132787# XM1/a_n100_n163683# 0.01363f
C6196 XM4/a_100_128582# m1_1634_n2388# 6.1e-20
C6197 XM2/a_n158_n139590# XM3/a_n100_67361# 7.26e-20
C6198 XM2/a_100_n250302# XM3/a_n100_n43491# 0.005074f
C6199 XM1/a_100_n12806# XM2/a_n158_n165950# 0.072463f
C6200 XM1/a_100_38890# XM3/a_n100_89117# 6.97e-21
C6201 XM1/a_n100_33049# XM3/a_n158_85070# 2.85e-20
C6202 XM4/w_n358_n132787# XM4/a_n100_54929# -0.004445f
C6203 XM1/a_100_n75990# XM2/a_100_n229214# 4.64e-21
C6204 XM2/a_n158_n181766# XM3/a_n100_24885# 7.26e-20
C6205 XM1/a_n100_n149323# XM3/a_n158_n98302# 2.85e-20
C6206 XM3/a_n100_n51779# m1_1634_n2388# 0.072015f
C6207 XM1/a_n100_35921# XM4/w_n358_n132787# 0.013564f
C6208 XM1/a_n100_n170863# XM2/a_100_n324110# 7.26e-20
C6209 XM2/a_100_n134318# XM3/a_n158_72638# 0.02378f
C6210 XM1/a_n158_n32910# XM2/a_n158_n187038# 9.28e-21
C6211 XM4/w_n358_n132787# XM3/a_n158_n124202# 0.032295f
C6212 XM4/a_n100_n110831# m1_1634_n2388# 0.072015f
C6213 XM1/a_n100_79001# XM3/a_n100_130557# 6.5e-19
C6214 XM2/a_n100_n100147# XM4/a_100_106826# 2.56e-20
C6215 XM4/a_n100_21# m1_1634_n2388# 0.072015f
C6216 XM1/a_n158_n7062# XM2/a_n158_n160678# 9.28e-21
C6217 XM1/a_n100_113465# XM2/a_100_n39422# 7.26e-20
C6218 XM1/a_100_60430# XM3/a_n158_112006# 0.00544f
C6219 XM3/a_n100_97405# m1_1634_n2388# 0.072015f
C6220 XM1/a_n100_n180915# XM3/a_n158_n130418# 2.85e-20
C6221 XM2/a_100_n176494# XM3/a_n158_30162# 0.05299f
C6222 XM1/a_n100_n14339# XM3/a_n100_37317# 5.33e-19
C6223 XM1/a_n100_25869# XM3/a_n158_76782# 2.85e-20
C6224 XM1/a_n100_15817# XM3/a_n100_67361# 2.98e-19
C6225 XM1/a_n158_n166458# XM2/a_n100_n321571# 7.26e-20
C6226 XM1/a_n100_n147887# XM2/a_100_n300386# 7.26e-20
C6227 XM1/a_100_n68810# XM2/a_n158_n223942# 0.084537f
C6228 XM2/a_100_n118502# m1_1634_n2388# 0.017213f
C6229 XM1/a_100_n152098# XM2/a_n100_n305755# 8.19e-19
C6230 XM1/a_n100_n146451# XM3/a_n158_n95194# 1.26e-20
C6231 XM2/a_100_n281934# XM3/a_n158_n77582# 0.034296f
C6232 XM3/a_n100_42497# m1_1634_n2388# 0.072015f
C6233 XM1/a_n100_173777# XM2/a_n158_18570# 0.005074f
C6234 XM2/a_n100_n287303# XM4/a_100_n82762# 2.56e-20
C6235 XM4/w_n358_n132787# XM4/a_n100_n16555# -0.004445f
C6236 XM2/a_100_n324110# XM3/a_n100_n119119# 0.010147f
C6237 XM4/w_n358_n132787# XM2/a_n158_n187038# 0.107093f
C6238 XM1/a_n100_n5723# XM4/w_n358_n132787# 0.013471f
C6239 XM1/a_100_53250# XM3/a_n158_103718# 1.53e-19
C6240 XM1/a_n100_n58855# XM4/w_n358_n132787# 0.013398f
C6241 XM1/a_n100_n50239# XM2/a_n158_n202854# 0.005074f
C6242 XM4/a_100_89214# m1_1634_n2388# 6.1e-20
C6243 XM1/a_100_5862# XM3/a_n158_57098# 0.004233f
C6244 XM1/a_n100_33049# XM2/a_n158_n121138# 0.010147f
C6245 XM1/a_n100_n114859# XM2/a_n158_n268754# 0.010147f
C6246 XM1/a_n158_n45834# XM2/a_n158_n200218# 9.28e-21
C6247 XM1/a_n100_66077# XM3/a_n158_117186# 2.85e-20
C6248 XM4/w_n358_n132787# XM3/a_n158_84034# 0.032295f
C6249 XM4/w_n358_n132787# XM4/a_n100_15561# -0.004445f
C6250 XM4/w_n358_n132787# XM3/a_n158_119258# 0.032295f
C6251 XM3/a_n100_n91147# m1_1634_n2388# 0.072015f
C6252 XM4/w_n358_n132787# XM3/a_n158_n1954# 0.032295f
C6253 XM4/w_n358_n132787# XM3/a_n158_29126# 0.032295f
C6254 XM3/a_n100_55965# XM4/a_n100_55965# 0.009521f
C6255 XM2/a_n158_n18334# XM1/a_100_135102# 0.100894f
C6256 XM1/a_100_76226# XM4/w_n358_n132787# 0.054997f
C6257 XM2/a_n158_n118502# XM3/a_n158_86106# 4.64e-21
C6258 XM2/a_100_n231850# XM3/a_n100_n25879# 0.010147f
C6259 XM2/a_100_n92142# XM3/a_n158_112006# 0.014433f
C6260 XM2/a_n100_n229311# XM3/a_n158_n24746# 0.005074f
C6261 XM1/a_100_n37218# XM2/a_n158_n189674# 0.005476f
C6262 XM2/a_n158_n160678# XM3/a_n158_43630# 4.64e-21
C6263 XM1/a_100_n31474# XM2/a_n158_n184402# 0.051432f
C6264 XM4/w_n358_n132787# XM4/a_n100_n55923# -0.004445f
C6265 XM3/a_n158_n26818# m1_1634_n2388# 6.1e-20
C6266 XM1/a_100_130794# XM4/w_n358_n132787# 0.048442f
C6267 XM1/a_100_27402# XM4/w_n358_n132787# 0.048442f
C6268 XM4/a_100_49846# m1_1634_n2388# 6.1e-20
C6269 XM2/a_n158_n226578# XM3/a_n158_n19566# 4.64e-21
C6270 XM4/w_n358_n132787# XM2/a_100_n123774# 0.103341f
C6271 XM2/a_100_n242394# m1_1634_n2388# 0.023309f
C6272 XM1/a_n100_n63163# XM4/w_n358_n132787# 0.01363f
C6273 XM3/a_n100_n130515# m1_1634_n2388# 0.072015f
C6274 XM4/w_n358_n132787# XM2/a_n158_n310930# 0.107093f
C6275 XM3/a_n158_67458# m1_1634_n2388# 6.1e-20
C6276 XM2/a_100_n305658# XM3/a_n100_n101507# 0.005074f
C6277 XM1/a_n158_n134866# XM3/a_n100_n82859# 1.94e-20
C6278 XM3/a_n158_12550# m1_1634_n2388# 6.1e-20
C6279 XM1/a_n100_n21519# XM3/a_n158_29126# 2.85e-20
C6280 XM1/a_n100_60333# XM2/a_n158_n92142# 0.005074f
C6281 XM4/a_n100_112945# m1_1634_n2388# 0.072015f
C6282 XM4/w_n358_n132787# XM3/a_n100_n36239# 0.009186f
C6283 XM4/a_100_n21638# m1_1634_n2388# 6.1e-20
C6284 XM1/a_100_n30038# XM3/a_n100_20741# 2.85e-20
C6285 XM2/a_n158_n76326# XM3/a_n100_129521# 1.45e-19
C6286 XM1/a_n100_47409# XM3/a_n158_98538# 2.85e-20
C6287 XM1/a_n100_n173735# m1_1634_n2388# 9.25e-20
C6288 XM1/a_n158_14478# XM2/a_n158_n139590# 9.28e-21
C6289 XM4/w_n358_n132787# XM4/a_n100_n95291# -0.004445f
C6290 XM1/a_100_n167894# XM3/a_n100_n116011# 2.85e-20
C6291 XM3/a_n158_n66186# m1_1634_n2388# 6.1e-20
C6292 XM2/a_n100_n155503# XM4/a_100_48810# 2.56e-20
C6293 XM1/a_100_53250# XM2/a_n100_n102783# 0.005074f
C6294 XM4/a_100_10478# m1_1634_n2388# 6.1e-20
C6295 XM1/a_n100_n179479# XM2/a_n158_n334654# 0.005074f
C6296 XM2/a_100_n213398# XM3/a_n100_n8267# 0.010147f
C6297 XM4/w_n358_n132787# XM1/a_n100_135005# 0.011815f
C6298 XM1/a_n158_n133430# XM3/a_n100_n81823# 1.94e-20
C6299 XM1/a_n158_n15678# XM2/a_n100_n171319# 7.26e-20
C6300 XM1/a_n158_5862# XM2/a_n100_n150231# 7.26e-20
C6301 XM1/a_n158_n71682# XM3/a_n100_n20699# 1.94e-20
C6302 XM2/a_n100_n181863# m1_1634_n2388# 7.61e-19
C6303 XM1/a_n158_148026# XM2/a_n100_n7887# 7.26e-20
C6304 XM1/a_n100_n162247# XM3/a_n158_n111770# 2.35e-20
C6305 XM1/a_n158_41762# XM3/a_n100_92225# 1.94e-20
C6306 XM1/a_n100_35921# XM3/a_n158_88178# 2.85e-20
C6307 XM4/w_n358_n132787# XM2/a_100_n247666# 0.103894f
C6308 XM1/a_n100_114901# XM2/a_n158_n39422# 0.010147f
C6309 XM3/a_n100_121233# m1_1634_n2388# 0.072015f
C6310 XM2/a_n100_n337387# XM3/a_n158_n130418# 0.005074f
C6311 XM4/a_n100_73577# m1_1634_n2388# 0.072015f
C6312 XM4/w_n358_n132787# XM3/a_n100_n75607# 0.008666f
C6313 XM4/a_100_n61006# m1_1634_n2388# 6.1e-20
C6314 XM2/a_n158_n250302# XM3/a_n100_n43491# 7.26e-20
C6315 XM1/a_100_n12806# XM2/a_n100_n166047# 0.005074f
C6316 XM1/a_n100_n15775# XM3/a_n158_35342# 2.85e-20
C6317 XM1/a_n100_79001# XM2/a_100_n73690# 7.26e-20
C6318 XM1/a_100_n75990# XM2/a_n158_n229214# 0.080252f
C6319 XM1/a_100_31710# XM3/a_n100_83937# 2.85e-20
C6320 XM3/a_n158_n105554# m1_1634_n2388# 6.1e-20
C6321 XM1/a_n100_116337# XM2/a_100_n36786# 7.26e-20
C6322 XM1/a_n100_n170863# XM2/a_n158_n324110# 0.005074f
C6323 XM2/a_n158_n134318# XM3/a_n158_72638# 4.64e-21
C6324 XM1/a_100_n48706# XM3/a_n100_2093# 2.85e-20
C6325 XM1/a_100_83406# XM4/w_n358_n132787# 0.048442f
C6326 XM3/a_n100_123305# XM4/a_n100_123305# 0.009521f
C6327 XM1/a_100_60430# XM3/a_n100_111909# 3.64e-20
C6328 XM1/a_n100_n91883# XM4/w_n358_n132787# 0.013446f
C6329 XM2/a_n158_n176494# XM3/a_n158_30162# 4.64e-21
C6330 XM4/w_n358_n132787# XM3/a_n158_n11278# 0.033579f
C6331 XM1/a_n100_n147887# XM2/a_n158_n300386# 0.005074f
C6332 XM1/a_100_n68810# XM2/a_n100_n224039# 0.005074f
C6333 XM4/w_n358_n132787# XM3/a_n100_77721# 0.009186f
C6334 XM2/a_n158_n281934# XM3/a_n158_n77582# 4.64e-21
C6335 XM3/a_n100_23849# XM4/a_n100_23849# 0.009521f
C6336 XM1/a_n158_n11370# XM2/a_n158_n165950# 9.28e-21
C6337 XM1/a_100_23094# XM3/a_n100_73577# 2.85e-20
C6338 XM2/a_n158_n324110# XM3/a_n100_n119119# 1.45e-19
C6339 XM4/w_n358_n132787# XM2/a_n100_n187135# 0.024763f
C6340 XM1/a_100_53250# XM3/a_n100_103621# 3.31e-19
C6341 XM2/a_n100_n305755# m1_1634_n2388# 0.002432f
C6342 XM1/a_n158_n142046# XM3/a_n100_n91147# 1.94e-20
C6343 XM4/w_n358_n132787# XM3/a_n100_22813# 0.008008f
C6344 XM4/a_n100_34209# m1_1634_n2388# 0.072015f
C6345 XM4/a_100_n100374# m1_1634_n2388# 6.1e-20
C6346 XM4/w_n358_n132787# XM3/a_n100_n114975# 0.008117f
C6347 XM1/a_n100_147929# XM2/a_100_n7790# 7.26e-20
C6348 XM1/a_100_47506# m1_1634_n2388# 0.002487f
C6349 XM2/a_100_n279298# XM3/a_n158_n72402# 0.029622f
C6350 XM1/a_100_n117634# XM4/w_n358_n132787# 0.048442f
C6351 XM4/w_n358_n132787# XM3/a_n100_119161# 0.00903f
C6352 XM2/a_n100_n284667# XM4/a_100_n77582# 2.56e-20
C6353 XM1/a_100_n15678# XM2/a_100_n171222# 4.64e-21
C6354 XM1/a_n100_166597# XM2/a_100_13298# 7.26e-20
C6355 XM1/a_100_73354# XM3/a_n158_125474# 0.003891f
C6356 XM4/w_n358_n132787# XM4/a_n100_128485# -0.004445f
C6357 XM2/a_n100_n118599# XM3/a_n158_86106# 0.005074f
C6358 XM2/a_n158_n231850# XM3/a_n100_n25879# 1.45e-19
C6359 XM2/a_n158_n92142# XM3/a_n158_112006# 4.64e-21
C6360 XM2/a_100_n92142# XM3/a_n100_111909# 0.005074f
C6361 XM2/a_n158_n65782# XM4/w_n358_n132787# 0.101988f
C6362 XM1/a_n158_n127686# XM3/a_n100_n76643# 1.94e-20
C6363 XM4/w_n358_n132787# XM3/a_n158_n50646# 0.032295f
C6364 XM4/a_n100_n37275# m1_1634_n2388# 0.072015f
C6365 XM1/a_n158_n17114# XM3/a_n100_34209# 3.89e-20
C6366 XM1/a_100_n123378# XM2/a_100_n279298# 4.64e-21
C6367 XM1/a_100_n37218# XM2/a_n100_n189771# 0.005074f
C6368 XM2/a_n100_n160775# XM3/a_n158_43630# 0.005074f
C6369 XM3/a_n158_118# m1_1634_n2388# 6.1e-20
C6370 XM1/a_100_n31474# XM2/a_n100_n184499# 0.005074f
C6371 XM3/a_n100_61145# m1_1634_n2388# 0.072015f
C6372 XM2/a_n100_n226675# XM3/a_n158_n19566# 0.005074f
C6373 XM4/w_n358_n132787# XM2/a_n158_n123774# 0.107093f
C6374 XM2/a_n158_n242394# m1_1634_n2388# 5.91e-22
C6375 XM1/a_n158_123614# XM2/a_n158_n28878# 4.64e-21
C6376 XM1/a_n158_n120506# XM3/a_n100_n68355# 1.94e-20
C6377 XM3/a_n100_6237# XM4/a_n100_6237# 0.009521f
C6378 XM3/a_n100_106729# XM4/a_n100_106729# 0.009521f
C6379 XM4/w_n358_n132787# XM2/a_n100_n311027# 0.024295f
C6380 XM2/a_n158_n305658# XM3/a_n100_n101507# 7.26e-20
C6381 XM4/w_n358_n132787# XM4/a_n100_89117# -0.004445f
C6382 XM1/a_100_n139174# XM2/a_100_n295114# 4.64e-21
C6383 XM3/a_n100_n17591# m1_1634_n2388# 0.072015f
C6384 XM1/a_n100_n33007# XM3/a_n100_18669# 2.73e-19
C6385 XM4/w_n358_n132787# XM3/a_n158_47774# 0.032295f
C6386 XM2/a_100_n76326# XM3/a_n158_130654# 0.021444f
C6387 XM4/w_n358_n132787# XM3/a_n158_n90014# 0.032295f
C6388 XM4/a_n100_n76643# m1_1634_n2388# 0.072015f
C6389 XM2/a_100_n260846# XM3/a_n158_n54790# 0.077916f
C6390 XM1/a_n100_74693# XM2/a_100_n78962# 1.45e-19
C6391 XM1/a_n100_n182351# XM4/w_n358_n132787# 0.01363f
C6392 XM2/a_100_n303022# XM3/a_n100_n96327# 0.005074f
C6393 XM1/a_100_81970# XM2/a_100_n73690# 4.64e-21
C6394 XM1/a_n100_n73215# XM2/a_100_n229214# 7.48e-22
C6395 XM1/a_n158_n55886# XM3/a_n100_n4123# 1.94e-20
C6396 XM1/a_n100_129261# XM2/a_n158_n26242# 0.005074f
C6397 XM1/a_n100_119209# XM2/a_100_n36786# 3.74e-21
C6398 XM1/a_n158_84842# XM2/a_n158_n68418# 4.64e-21
C6399 XM1/a_100_53250# XM2/a_100_n100050# 4.64e-21
C6400 XM1/a_100_10170# XM2/a_100_n144862# 4.64e-21
C6401 XM1/a_100_165258# XM2/a_n158_10662# 0.116862f
C6402 XM1/a_100_44634# XM3/a_n100_95333# 2.85e-20
C6403 XM2/a_n158_n213398# XM3/a_n100_n8267# 1.45e-19
C6404 XM1/a_n100_n47367# m1_1634_n2388# 1.07e-19
C6405 XM1/a_100_123614# XM2/a_n158_n31514# 0.084926f
C6406 XM1/a_n158_n18550# XM3/a_n100_32137# 1.94e-20
C6407 XM1/a_n100_169469# XM2/a_n100_15837# 0.003522f
C6408 XM1/a_n100_n99063# XM3/a_n158_n48574# 2.7e-20
C6409 XM2/a_100_n179130# m1_1634_n2388# 0.024627f
C6410 XM2/a_n100_n152867# XM4/a_100_53990# 2.56e-20
C6411 XM4/a_100_123402# m1_1634_n2388# 6.1e-20
C6412 XM4/w_n358_n132787# XM2/a_n158_n247666# 0.107093f
C6413 XM4/w_n358_n132787# XM4/a_n100_49749# -0.004445f
C6414 XM3/a_n158_86106# m1_1634_n2388# 6.1e-20
C6415 XM2/a_100_n334654# XM3/a_n158_n130418# 0.023001f
C6416 XM3/a_n100_n56959# m1_1634_n2388# 0.072015f
C6417 XM2/a_100_n136954# XM3/a_n100_67361# 0.005074f
C6418 XM4/a_n100_n116011# m1_1634_n2388# 0.072014f
C6419 XM1/a_n158_n143482# XM3/a_n100_n92183# 3.89e-20
C6420 XM3/a_n158_31198# m1_1634_n2388# 6.1e-20
C6421 XM4/w_n358_n132787# XM3/a_n158_n129382# 0.032295f
C6422 XM3/a_n100_n10339# XM4/a_n100_n10339# 0.009521f
C6423 XM1/a_n100_n34443# XM4/w_n358_n132787# 0.01363f
C6424 XM1/a_100_n75990# XM2/a_n100_n229311# 0.005074f
C6425 XM2/a_100_n179130# XM3/a_n100_24885# 0.005074f
C6426 XM3/a_n100_6237# m1_1634_n2388# 0.072015f
C6427 XM3/a_n100_76685# XM4/a_n100_76685# 0.009521f
C6428 XM2/a_n100_n134415# XM3/a_n158_72638# 0.005074f
C6429 XM1/a_100_n27166# XM3/a_n100_24885# 2.85e-20
C6430 XM1/a_n100_58897# XM3/a_n158_110970# 2.85e-20
C6431 XM4/w_n358_n132787# XM4/a_n100_n21735# -0.004445f
C6432 XM1/a_100_176746# XM2/a_100_21206# 4.64e-21
C6433 XM2/a_100_n242394# XM3/a_n158_n37178# 0.077916f
C6434 XM2/a_n100_n176591# XM3/a_n158_30162# 0.005074f
C6435 XM4/a_100_84034# m1_1634_n2388# 6.1e-20
C6436 XM2/a_100_n284570# XM3/a_n100_n78715# 0.010147f
C6437 XM1/a_100_104946# XM2/a_n158_n49966# 0.105957f
C6438 XM1/a_100_n68810# XM2/a_100_n221306# 4.64e-21
C6439 XM2/a_n100_n118599# m1_1634_n2388# 7.61e-19
C6440 XM1/a_n158_8734# XM3/a_n100_59073# 1.94e-20
C6441 XM2/a_n100_n282031# XM3/a_n158_n77582# 0.005074f
C6442 XM4/w_n358_n132787# XM4/a_n100_10381# -0.004445f
C6443 XM1/a_n100_51717# XM3/a_n158_102682# 2.85e-20
C6444 XM1/a_n100_n111987# XM3/a_n158_n59970# 2.85e-20
C6445 XM3/a_n100_n96327# m1_1634_n2388# 0.072015f
C6446 XM4/a_n100_6237# m1_1634_n2388# 0.072015f
C6447 XM4/w_n358_n132787# XM2/a_100_n184402# 0.105152f
C6448 XM2/a_100_n303022# m1_1634_n2388# 0.017213f
C6449 XM3/a_n100_n30023# XM4/a_n100_n30023# 0.009521f
C6450 XM1/a_n158_1554# XM3/a_n100_52857# 3.89e-20
C6451 XM1/a_n100_76129# XM4/w_n358_n132787# 0.013471f
C6452 XM2/a_100_n123774# XM3/a_n100_81865# 0.010147f
C6453 XM1/a_100_15914# XM3/a_n100_66325# 2.85e-20
C6454 XM2/a_n158_n279298# XM3/a_n158_n72402# 4.64e-21
C6455 XM1/a_n100_n76087# XM4/w_n358_n132787# 0.013462f
C6456 XM1/a_100_n15678# XM2/a_n158_n171222# 0.044422f
C6457 XM1/a_n158_n111890# XM3/a_n100_n61103# 1.94e-20
C6458 XM2/a_100_n165950# XM3/a_n100_39389# 0.010147f
C6459 XM1/a_100_73354# XM3/a_n100_125377# 2.85e-20
C6460 XM1/a_n158_n137738# XM3/a_n100_n87003# 1.94e-20
C6461 XM1/a_n100_106285# XM2/a_n158_n47330# 0.010147f
C6462 XM4/w_n358_n132787# XM4/a_n100_n61103# -0.004445f
C6463 XM3/a_n158_n31998# m1_1634_n2388# 6.1e-20
C6464 XM1/a_100_n4190# XM3/a_n100_46641# 2.85e-20
C6465 XM2/a_n158_n92142# XM3/a_n100_111909# 7.26e-20
C6466 XM2/a_n100_n92239# XM3/a_n158_112006# 0.005074f
C6467 XM1/a_100_n127686# XM2/a_n158_n281934# 0.116862f
C6468 XM1/a_100_24530# XM4/w_n358_n132787# 0.049202f
C6469 XM4/a_100_44666# m1_1634_n2388# 6.1e-20
C6470 XM1/a_100_n123378# XM2/a_n158_n279298# 0.007812f
C6471 XM1/a_n100_n160811# XM2/a_100_n316202# 7.26e-20
C6472 XM4/w_n358_n132787# XM3/a_n100_96369# 0.009173f
C6473 XM1/a_n158_n170766# XM2/a_n158_n326746# 4.64e-21
C6474 XM1/a_n100_182393# XM4/w_n358_n132787# 0.012096f
C6475 XM2/a_100_n223942# XM3/a_n158_n19566# 0.036633f
C6476 XM1/a_100_171002# XM2/a_n158_18570# 0.003139f
C6477 XM4/w_n358_n132787# XM2/a_n100_n123871# 0.025738f
C6478 XM3/a_n100_n49707# XM4/a_n100_n49707# 0.009521f
C6479 XM2/a_n100_n242491# m1_1634_n2388# 0.002646f
C6480 XM2/a_n100_n229311# XM4/a_100_n24746# 2.56e-20
C6481 XM4/w_n358_n132787# XM3/a_n100_41461# 0.009023f
C6482 XM1/a_100_99202# XM4/w_n358_n132787# 0.048442f
C6483 XM1/a_n158_73354# XM2/a_n100_n79059# 1.37e-20
C6484 XM2/a_100_n266118# XM3/a_n100_n61103# 0.010147f
C6485 XM4/a_n100_n132587# XM3/a_n100_n132587# 0.01485f
C6486 XM1/a_100_n80298# XM4/w_n358_n132787# 0.048442f
C6487 XM4/a_n100_107765# m1_1634_n2388# 0.072015f
C6488 XM2/a_100_n110594# XM3/a_n100_96369# 0.005074f
C6489 XM4/w_n358_n132787# XM2/a_100_n308294# 0.103447f
C6490 XM4/w_n358_n132787# XM3/a_n100_n41419# 0.009115f
C6491 XM4/a_100_n26818# m1_1634_n2388# 6.1e-20
C6492 XM4/w_n358_n132787# XM4/a_n100_n100471# -0.004445f
C6493 XM1/a_100_n139174# XM2/a_n158_n295114# 0.005865f
C6494 XM1/a_n100_n66035# XM3/a_n100_n13447# 7.8e-20
C6495 XM2/a_100_n152770# XM3/a_n100_53893# 0.005074f
C6496 XM3/a_n158_n71366# m1_1634_n2388# 6.1e-20
C6497 XM1/a_n100_94797# XM2/a_n158_n60510# 0.005074f
C6498 XM2/a_n158_n76326# XM3/a_n158_130654# 4.64e-21
C6499 XM2/a_100_n76326# XM3/a_n100_130557# 0.005074f
C6500 XM1/a_100_47506# XM3/a_n100_98441# 6.08e-19
C6501 XM1/a_n158_57558# XM2/a_n158_n97414# 4.64e-21
C6502 XM2/a_100_n194946# XM3/a_n100_11417# 0.005074f
C6503 XM2/a_n158_n18334# XM4/w_n358_n132787# 0.101988f
C6504 XM1/a_n100_74693# XM2/a_n158_n78962# 0.010147f
C6505 XM1/a_100_58994# XM4/w_n358_n132787# 0.048442f
C6506 XM2/a_n158_n303022# XM3/a_n100_n96327# 7.26e-20
C6507 XM1/a_n158_92022# XM2/a_n100_n60607# 7.26e-20
C6508 XM1/a_n100_n73215# XM2/a_n158_n229214# 2.49e-20
C6509 XM1/a_100_53250# XM2/a_n158_n100050# 0.087652f
C6510 XM1/a_100_10170# XM2/a_n158_n144862# 0.094273f
C6511 XM1/a_n100_n179479# XM2/a_100_n332018# 7.26e-20
C6512 XM3/a_n100_79793# m1_1634_n2388# 0.072015f
C6513 XM3/a_n100_n69391# XM4/a_n100_n69391# 0.009521f
C6514 XM1/a_n158_n15678# XM2/a_n158_n168586# 4.64e-21
C6515 XM1/a_n158_5862# XM2/a_n158_n147498# 4.64e-21
C6516 XM1/a_n158_n61630# XM2/a_n158_n216034# 9.28e-21
C6517 XM2/a_n158_n179130# m1_1634_n2388# 2.36e-21
C6518 XM4/a_n100_68397# m1_1634_n2388# 0.072015f
C6519 XM4/w_n358_n132787# XM3/a_n100_n80787# 0.008583f
C6520 XM4/a_100_n66186# m1_1634_n2388# 6.1e-20
C6521 XM3/a_n100_24885# m1_1634_n2388# 0.072015f
C6522 XM4/w_n358_n132787# XM2/a_n100_n247763# 0.026677f
C6523 XM1/a_100_n75990# XM3/a_n100_n24843# 4.23e-20
C6524 XM1/a_n158_n57322# XM3/a_n100_n6195# 2e-20
C6525 XM3/a_n100_44569# XM4/a_n100_44569# 0.009521f
C6526 XM3/a_n158_122366# m1_1634_n2388# 6.1e-20
C6527 XM2/a_n158_n334654# XM3/a_n158_n130418# 4.64e-21
C6528 XM3/a_n158_n110734# m1_1634_n2388# 6.1e-20
C6529 XM1/a_100_n159278# XM3/a_n100_n108759# 2.85e-20
C6530 XM2/a_n158_n136954# XM3/a_n100_67361# 7.26e-20
C6531 XM4/w_n358_n132787# XM3/a_n158_66422# 0.032295f
C6532 XM2/a_100_n247666# XM3/a_n100_n43491# 0.005074f
C6533 XM1/a_n100_112029# XM2/a_100_n42058# 1.45e-19
C6534 XM1/a_n158_46070# XM2/a_n158_n107958# 9.28e-21
C6535 XM1/a_n100_170905# XM4/w_n358_n132787# 0.012279f
C6536 XM1/a_n158_n182254# XM3/a_n100_n131551# 1.94e-20
C6537 XM4/w_n358_n132787# XM3/a_n158_11514# 0.033716f
C6538 XM2/a_n158_n179130# XM3/a_n100_24885# 7.26e-20
C6539 XM2/a_n158_29114# XM4/w_n358_n132787# 0.061385f
C6540 XM2/a_100_n332018# XM3/a_n158_n125238# 0.040917f
C6541 XM1/a_100_n152098# XM3/a_n100_n101507# 2.85e-20
C6542 XM4/w_n358_n132787# XM3/a_n158_n16458# 0.032295f
C6543 XM4/a_n100_n3087# m1_1634_n2388# 0.072015f
C6544 XM1/a_n158_118# XM2/a_n158_n155406# 4.64e-21
C6545 XM2/a_100_n131682# XM3/a_n158_72638# 0.03118f
C6546 XM1/a_n100_n40187# m1_1634_n2388# 2.05e-19
C6547 XM3/a_n100_n89075# XM4/a_n100_n89075# 0.009521f
C6548 XM1/a_n100_79001# XM3/a_n100_131593# 2.6e-20
C6549 XM2/a_n100_n97511# XM4/a_100_106826# 2.56e-20
C6550 XM1/a_n100_n133527# XM2/a_100_n287206# 1.45e-19
C6551 XM2/a_100_n173858# XM3/a_n158_30162# 0.00197f
C6552 XM4/a_n100_29029# m1_1634_n2388# 0.072015f
C6553 XM4/w_n358_n132787# XM3/a_n100_n120155# 0.009186f
C6554 XM1/a_n158_n166458# XM2/a_n100_n318935# 5.76e-20
C6555 XM4/a_100_n105554# m1_1634_n2388# 6.1e-20
C6556 XM2/a_n158_n284570# XM3/a_n100_n78715# 1.45e-19
C6557 XM1/a_100_n68810# XM2/a_n158_n221306# 0.00937f
C6558 XM1/a_n158_n12806# XM3/a_n100_39389# 1.94e-20
C6559 XM1/a_n158_66174# XM3/a_n100_117089# 1.94e-20
C6560 XM2/a_100_n115866# m1_1634_n2388# 0.025819f
C6561 XM1/a_n100_n182351# XM3/a_n158_n131454# 2.85e-20
C6562 XM1/a_100_n137738# XM3/a_n100_n87003# 2.85e-20
C6563 XM1/a_n158_n110454# XM3/a_n100_n60067# 1.94e-20
C6564 XM1/a_n100_n169427# m1_1634_n2388# 1.67e-20
C6565 XM4/w_n358_n132787# XM2/a_n158_n184402# 0.107093f
C6566 XM1/a_n100_67513# m1_1634_n2388# 9.68e-20
C6567 XM1/a_100_1554# XM3/a_n100_51821# 1.87e-20
C6568 XM4/w_n358_n132787# XM4/a_n100_123305# -0.004445f
C6569 XM1/a_n158_n28602# XM3/a_n100_21777# 1.94e-20
C6570 XM1/a_n100_n160811# XM3/a_n158_n108662# 2.85e-20
C6571 XM1/a_n100_104849# XM4/w_n358_n132787# 0.011611f
C6572 XM1/a_n100_66077# XM3/a_n158_118222# 2.85e-20
C6573 XM2/a_n158_n123774# XM3/a_n100_81865# 1.45e-19
C6574 XM2/a_n100_n279395# XM3/a_n158_n72402# 0.005074f
C6575 XM1/a_100_n15678# XM2/a_n100_n171319# 0.005074f
C6576 XM3/a_n158_49846# m1_1634_n2388# 6.1e-20
C6577 XM4/w_n358_n132787# XM3/a_n158_120294# 0.038462f
C6578 XM1/a_n158_n37218# XM2/a_n158_n192310# 4.64e-21
C6579 XM4/w_n358_n132787# XM3/a_n158_n55826# 0.032295f
C6580 XM4/a_n100_n42455# m1_1634_n2388# 0.072015f
C6581 XM1/a_n100_63205# XM4/w_n358_n132787# 0.01363f
C6582 XM2/a_n158_n165950# XM3/a_n100_39389# 1.45e-19
C6583 XM1/a_100_n58758# XM3/a_n100_n7231# 2.85e-20
C6584 XM2/a_100_n92142# XM3/a_n158_113042# 0.077916f
C6585 XM2/a_100_n118502# XM3/a_n158_87142# 0.077916f
C6586 XM3/a_n100_n108759# XM4/a_n100_n108759# 0.009521f
C6587 XM1/a_100_30274# XM2/a_n158_n123774# 0.116862f
C6588 XM1/a_100_n123378# XM2/a_n100_n279395# 0.005074f
C6589 XM1/a_n100_n50239# XM3/a_n100_21# 6.5e-19
C6590 XM2/a_100_n160678# XM3/a_n158_44666# 0.077916f
C6591 XM2/a_100_n313566# XM3/a_n158_n107626# 0.077916f
C6592 XM1/a_100_64738# XM2/a_n158_n89506# 0.116862f
C6593 XM1/a_100_n179382# XM3/a_n100_n128443# 4.69e-20
C6594 XM1/a_n100_n160811# XM2/a_n158_n316202# 0.005074f
C6595 XM4/w_n358_n132787# XM1/a_100_n156406# 0.048442f
C6596 XM1/a_n158_n170766# XM2/a_n100_n326843# 7.26e-20
C6597 XM2/a_n158_n223942# XM3/a_n158_n19566# 4.64e-21
C6598 XM4/w_n358_n132787# XM2/a_100_n121138# 0.106121f
C6599 XM4/w_n358_n132787# XM4/a_n100_83937# -0.004445f
C6600 XM2/a_100_n239758# m1_1634_n2388# 0.017213f
C6601 XM3/a_n100_n22771# m1_1634_n2388# 0.072015f
C6602 XM1/a_100_129358# XM4/w_n358_n132787# 0.053546f
C6603 XM1/a_n100_n150759# XM3/a_n158_n98302# 1.75e-19
C6604 XM2/a_n158_n266118# XM3/a_n100_n61103# 1.45e-19
C6605 XM2/a_n158_n110594# XM3/a_n100_96369# 7.26e-20
C6606 XM4/w_n358_n132787# XM2/a_n158_n308294# 0.10292f
C6607 XM4/w_n358_n132787# XM3/a_n158_n95194# 0.032295f
C6608 XM4/a_n100_n81823# m1_1634_n2388# 0.072015f
C6609 XM2/a_n100_n34247# XM4/w_n358_n132787# 0.012203f
C6610 XM2/a_100_n221306# XM3/a_n158_n14386# 0.027285f
C6611 XM1/a_100_n139174# XM2/a_n100_n295211# 0.005074f
C6612 XM1/a_n100_n101935# XM3/a_n158_n49610# 2.85e-20
C6613 XM2/a_n100_n226675# XM4/a_100_n19566# 2.56e-20
C6614 XM1/a_n100_n61727# XM3/a_n158_n11278# 1.52e-20
C6615 XM2/a_n158_n152770# XM3/a_n100_53893# 7.26e-20
C6616 sw_bn iout 0.001766f
C6617 XM3/a_n100_n128443# XM4/a_n100_n128443# 0.009521f
C6618 XM2/a_n100_n76423# XM3/a_n158_130654# 0.005074f
C6619 XM2/a_n158_n76326# XM3/a_n100_130557# 7.26e-20
C6620 XM1/a_100_92022# XM2/a_n100_n63243# 0.005074f
C6621 XM1/a_n158_57558# XM2/a_n100_n97511# 7.26e-20
C6622 XM2/a_n158_n194946# XM3/a_n100_11417# 7.26e-20
C6623 XM1/a_100_90586# XM4/w_n358_n132787# 0.048442f
C6624 XM1/a_100_n139174# XM3/a_n100_n88039# 3.87e-20
C6625 XM1/a_100_129358# XM2/a_n100_n26339# 0.005074f
C6626 XM1/a_n100_51717# XM2/a_100_n102686# 1.45e-19
C6627 XM1/a_100_n172202# XM3/a_n100_n120155# 2.85e-20
C6628 XM1/a_100_n110454# XM3/a_n100_n59031# 5.29e-20
C6629 XM1/a_n100_n104807# XM4/w_n358_n132787# 0.013028f
C6630 XM1/a_n100_n73215# XM2/a_n100_n229311# 0.005067f
C6631 XM4/a_100_118222# m1_1634_n2388# 6.1e-20
C6632 XM2/a_100_n147498# XM3/a_n158_59170# 0.051822f
C6633 XM1/a_100_53250# XM2/a_n100_n100147# 0.005074f
C6634 XM3/a_n100_97405# XM4/a_n100_97405# 0.009521f
C6635 XM1/a_100_10170# XM2/a_n100_n144959# 0.005074f
C6636 XM3/a_n100_12453# XM4/a_n100_12453# 0.009521f
C6637 XM1/a_n100_n7159# m1_1634_n2388# 7.54e-20
C6638 XM1/a_n100_179521# XM2/a_100_26478# 7.26e-20
C6639 XM1/a_n100_45973# XM3/a_n158_98538# 9.33e-21
C6640 XM1/a_n100_n179479# XM2/a_n158_n332018# 0.005074f
C6641 XM4/w_n358_n132787# XM4/a_n100_44569# -0.004445f
C6642 XM1/a_100_5862# XM2/a_100_n150134# 4.64e-21
C6643 XM3/a_n100_n62139# m1_1634_n2388# 0.072015f
C6644 XM2/a_100_n189674# XM3/a_n158_16694# 0.077916f
C6645 XM1/a_n158_n15678# XM2/a_n100_n168683# 7.26e-20
C6646 XM1/a_n158_5862# XM2/a_n100_n147595# 7.26e-20
C6647 XM2/a_n100_n179227# m1_1634_n2388# 8.58e-19
C6648 XM4/w_n358_n132787# XM3/a_n100_60109# 0.009186f
C6649 XM4/a_n100_n121191# m1_1634_n2388# 0.072015f
C6650 XM2/a_100_n295114# XM3/a_n158_n90014# 0.077916f
C6651 XM1/a_100_n160714# XM2/a_100_n316202# 4.64e-21
C6652 XM1/a_n100_41665# XM3/a_n158_92322# 2.85e-20
C6653 XM2/a_100_n337290# XM3/a_n100_n131551# 0.010147f
C6654 XM4/w_n358_n132787# XM2/a_100_n245030# 0.103341f
C6655 XM1/a_n158_n114762# XM3/a_n100_n63175# 1.94e-20
C6656 XM2/a_n100_13201# XM4/w_n358_n132787# 0.012074f
C6657 XM3/a_n100_122269# m1_1634_n2388# 0.072015f
C6658 XM2/a_n100_n334751# XM3/a_n158_n130418# 0.005074f
C6659 XM4/w_n358_n132787# XM1/a_n100_n156503# 0.01363f
C6660 XM2/a_n158_n247666# XM3/a_n100_n43491# 7.26e-20
C6661 XM4/w_n358_n132787# XM1/a_n100_n147887# 0.013481f
C6662 XM4/w_n358_n132787# XM4/a_n100_n26915# -0.004445f
C6663 XM1/a_n158_n73118# XM3/a_n100_n22771# 2e-22
C6664 XM1/a_n100_n53111# XM2/a_100_n208126# 7.26e-20
C6665 XM1/a_100_38890# XM3/a_n100_90153# 5.71e-20
C6666 XM1/a_n100_1457# XM4/w_n358_n132787# 0.013401f
C6667 XM1/a_n158_118# XM2/a_n100_n155503# 7.26e-20
C6668 XM4/a_100_78854# m1_1634_n2388# 6.1e-20
C6669 XM2/a_n158_n332018# XM3/a_n158_n125238# 4.64e-21
C6670 XM1/a_100_n80298# XM2/a_n158_n234486# 0.116862f
C6671 XM2/a_n158_n131682# XM3/a_n158_72638# 4.64e-21
C6672 XM2/a_100_n245030# XM3/a_n100_n38311# 0.005074f
C6673 XM1/a_100_n87478# XM4/w_n358_n132787# 0.051502f
C6674 XM3/a_n100_n101507# m1_1634_n2388# 0.072015f
C6675 XM3/a_n100_98441# m1_1634_n2388# 0.072015f
C6676 XM1/a_n100_n133527# XM2/a_n158_n287206# 0.010147f
C6677 XM1/a_n100_n120603# m1_1634_n2388# 1.08e-19
C6678 XM2/a_n158_n173858# XM3/a_n158_30162# 4.64e-21
C6679 XM1/a_n100_25869# XM3/a_n158_77818# 1.17e-19
C6680 XM1/a_n100_15817# XM3/a_n100_68397# 1.82e-19
C6681 XM1/a_100_n68810# XM2/a_n100_n221403# 0.005074f
C6682 XM1/a_n158_n153534# XM2/a_n158_n308294# 9.28e-21
C6683 XM2/a_n100_n202951# XM4/a_100_4262# 2.56e-20
C6684 XM3/a_n100_43533# m1_1634_n2388# 0.072015f
C6685 XM1/a_n100_173777# XM2/a_n158_21206# 0.005074f
C6686 XM1/a_100_n176510# XM4/w_n358_n132787# 0.054609f
C6687 XM2/a_n100_n94875# XM4/a_100_112006# 2.56e-20
C6688 XM4/w_n358_n132787# XM3/a_n100_n7231# 0.008953f
C6689 XM4/w_n358_n132787# XM2/a_n100_n184499# 0.024367f
C6690 XM1/a_100_53250# XM3/a_n100_104657# 3.44e-19
C6691 XM2/a_n100_n303119# m1_1634_n2388# 0.001171f
C6692 XM1/a_n100_n80395# XM3/a_n100_n30023# 3.64e-19
C6693 XM1/a_100_n70246# XM3/a_n100_n18627# 2.85e-20
C6694 XM4/w_n358_n132787# XM4/a_n100_n66283# -0.004445f
C6695 XM3/a_n158_n37178# m1_1634_n2388# 6.1e-20
C6696 XM4/w_n358_n132787# XM3/a_n158_85070# 0.032295f
C6697 XM2/a_100_n276662# XM3/a_n158_n72402# 0.025338f
C6698 XM1/a_n158_n37218# XM2/a_n100_n192407# 7.26e-20
C6699 XM1/a_100_n15678# XM2/a_100_n168586# 4.64e-21
C6700 XM4/w_n358_n132787# XM3/a_n100_120197# 0.00903f
C6701 XM2/a_n100_n282031# XM4/a_100_n77582# 2.56e-20
C6702 XM4/a_100_39486# m1_1634_n2388# 6.1e-20
C6703 XM1/a_n158_7298# XM3/a_n100_58037# 1.94e-20
C6704 XM2/a_100_n318838# XM3/a_n100_n113939# 0.010147f
C6705 XM1/a_n158_n162150# XM3/a_n100_n109795# 9.02e-21
C6706 XM1/a_100_n124814# XM2/a_n158_n279298# 0.116862f
C6707 XM4/w_n358_n132787# XM3/a_n158_30162# 0.038462f
C6708 XM1/a_n100_168033# XM2/a_100_13298# 7.26e-20
C6709 XM2/a_100_n92142# XM3/a_n100_112945# 0.010147f
C6710 XM1/a_100_n123378# XM2/a_100_n276662# 4.64e-21
C6711 XM1/a_n100_99105# XM2/a_100_n55238# 1.45e-19
C6712 XM1/a_n100_n54547# XM4/w_n358_n132787# 0.013139f
C6713 XM1/a_n100_n17211# XM4/w_n358_n132787# 0.013401f
C6714 XM4/a_n100_102585# m1_1634_n2388# 0.072015f
C6715 XM4/w_n358_n132787# XM3/a_n100_n46599# 0.009203f
C6716 XM4/a_100_n31998# m1_1634_n2388# 6.1e-20
C6717 XM2/a_100_n226578# XM3/a_n100_n20699# 0.010147f
C6718 XM2/a_n100_n224039# XM3/a_n158_n19566# 0.005074f
C6719 XM1/a_100_99202# XM2/a_n158_n55238# 0.116862f
C6720 XM4/w_n358_n132787# XM2/a_n158_n121138# 0.107093f
C6721 XM4/w_n358_n132787# XM4/a_n100_n105651# -0.004445f
C6722 XM3/a_n158_n76546# m1_1634_n2388# 6.1e-20
C6723 XM3/a_n158_7370# m1_1634_n2388# 6.1e-20
C6724 XM4/w_n358_n132787# XM2/a_n100_n308391# 0.02493f
C6725 XM3/a_n158_68494# m1_1634_n2388# 6.1e-20
C6726 XM1/a_100_69046# XM4/w_n358_n132787# 0.054609f
C6727 XM2/a_n158_n221306# XM3/a_n158_n14386# 4.64e-21
C6728 XM1/a_n100_17253# XM2/a_100_n136954# 1.45e-19
C6729 XM1/a_100_n139174# XM2/a_100_n292478# 4.64e-21
C6730 XM1/a_n100_n114859# XM3/a_n100_n63175# 1.69e-19
C6731 XM1/a_n100_n104807# XM3/a_n158_n52718# 2.85e-20
C6732 XM3/a_n100_65289# XM4/a_n100_65289# 0.009521f
C6733 XM3/a_n158_13586# m1_1634_n2388# 6.1e-20
C6734 XM1/a_n158_n21422# XM2/a_n158_n176494# 4.64e-21
C6735 XM1/a_n100_n8595# m1_1634_n2388# 7.54e-20
C6736 XM1/a_100_n30038# XM3/a_n100_21777# 2.85e-20
C6737 XM2/a_n100_n195043# XM3/a_n100_11417# 0.001572f
C6738 XM1/a_100_116434# XM4/w_n358_n132787# 0.053546f
C6739 XM1/a_n100_47409# XM3/a_n158_99574# 2.85e-20
C6740 XM2/a_100_n300386# XM3/a_n100_n96327# 0.005074f
C6741 XM1/a_n100_51717# XM2/a_n158_n102686# 0.010147f
C6742 XM1/a_n100_12945# XM4/w_n358_n132787# 0.013471f
C6743 XM1/a_n100_n73215# XM2/a_100_n226578# 7.26e-20
C6744 XM4/a_n100_63217# m1_1634_n2388# 0.072015f
C6745 XM2/a_n158_n147498# XM3/a_n158_59170# 4.64e-21
C6746 XM4/w_n358_n132787# XM3/a_n100_n85967# 0.008564f
C6747 XM4/a_100_n71366# m1_1634_n2388# 6.1e-20
C6748 XM1/a_100_5862# XM2/a_n158_n150134# 4.13e-19
C6749 XM1/a_n100_44537# XM3/a_n158_95430# 2.85e-20
C6750 XM1/a_n100_33049# m1_1634_n2388# 1.3e-19
C6751 XM1/a_n158_67610# XM2/a_n158_n86870# 9.28e-21
C6752 XM3/a_n158_n115914# m1_1634_n2388# 6.1e-20
C6753 XM1/a_n100_n35879# XM2/a_100_n189674# 1.45e-19
C6754 XM2/a_100_n176494# m1_1634_n2388# 0.017213f
C6755 XM2/a_n100_n150231# XM4/a_100_53990# 2.56e-20
C6756 XM1/a_n158_148026# XM2/a_n100_n5251# 7.26e-20
C6757 XM1/a_100_n160714# XM2/a_n158_n316202# 0.049874f
C6758 XM1/a_n158_41762# XM3/a_n100_93261# 1.94e-20
C6759 XM2/a_n158_n337290# XM3/a_n100_n131551# 1.45e-19
C6760 XM4/w_n358_n132787# XM2/a_n158_n245030# 0.104632f
C6761 XM1/a_n100_n132091# XM3/a_n100_n81823# 6.55e-19
C6762 XM1/a_n158_n124814# XM3/a_n100_n74571# 7.41e-21
C6763 XM1/a_n100_n27263# XM4/w_n358_n132787# 0.013602f
C6764 XM4/w_n358_n132787# XM3/a_n158_n21638# 0.032295f
C6765 XM4/a_n100_n8267# m1_1634_n2388# 0.072015f
C6766 XM1/a_n100_n53111# XM2/a_n158_n208126# 0.005074f
C6767 XM1/a_n158_n48706# XM3/a_n100_3129# 1.94e-20
C6768 XM1/a_n100_n15775# XM3/a_n158_36378# 2.85e-20
C6769 XM2/a_n158_n15698# XM1/a_n158_137974# 9.28e-21
C6770 XM1/a_100_36018# XM4/w_n358_n132787# 0.048442f
C6771 XM1/a_n100_n155067# XM2/a_100_n310930# 7.26e-20
C6772 XM4/a_n100_23849# m1_1634_n2388# 0.072015f
C6773 XM2/a_n100_n332115# XM3/a_n158_n125238# 0.005074f
C6774 XM4/w_n358_n132787# XM3/a_n100_n125335# 0.009106f
C6775 XM4/a_100_n110734# m1_1634_n2388# 6.1e-20
C6776 XM1/a_n158_n154970# XM3/a_n100_n103579# 2.18e-20
C6777 XM2/a_n100_n131779# XM3/a_n158_72638# 0.005074f
C6778 XM2/a_n158_n245030# XM3/a_n100_n38311# 7.26e-20
C6779 XM1/a_n100_n159375# m1_1634_n2388# 9.95e-20
C6780 XM2/a_n100_n173955# XM3/a_n158_30162# 0.005074f
C6781 XM4/w_n358_n132787# XM4/a_n100_118125# -0.004445f
C6782 XM1/a_100_n42962# XM3/a_n100_7273# 9.33e-21
C6783 XM2/a_n100_n115963# m1_1634_n2388# 7.61e-19
C6784 XM4/w_n358_n132787# XM3/a_n100_78757# 0.009186f
C6785 XM1/a_n100_12945# XM3/a_n100_63217# 6.65e-19
C6786 XM1/a_n100_51717# XM3/a_n158_103718# 2.85e-20
C6787 XM1/a_100_23094# XM3/a_n100_74613# 2.85e-20
C6788 XM4/w_n358_n132787# XM3/a_n158_n61006# 0.032295f
C6789 XM4/a_n100_n47635# m1_1634_n2388# 0.072015f
C6790 XM4/w_n358_n132787# XM2/a_100_n181766# 0.103342f
C6791 XM1/a_n158_104946# XM2/a_n158_n49966# 4.64e-21
C6792 XM1/a_100_33146# XM2/a_n158_n121138# 0.116862f
C6793 XM2/a_100_n300386# m1_1634_n2388# 0.023368f
C6794 XM1/a_n100_n51675# XM3/a_n158_118# 2.84e-20
C6795 XM4/w_n358_n132787# XM3/a_n100_23849# 0.009039f
C6796 XM1/a_n158_70482# XM3/a_n100_121233# 1.94e-20
C6797 XM1/a_n100_n129219# XM3/a_n100_n76643# 2.34e-19
C6798 XM1/a_n100_147929# XM2/a_100_n5154# 7.26e-20
C6799 XM2/a_n158_n276662# XM3/a_n158_n72402# 4.64e-21
C6800 XM1/a_100_n15678# XM2/a_n158_n168586# 0.049485f
C6801 XM3/a_n100_130557# XM4/a_n100_130557# 0.009521f
C6802 XM2/a_n158_n318838# XM3/a_n100_n113939# 1.45e-19
C6803 XM1/a_n100_n45931# XM4/w_n358_n132787# 0.013538f
C6804 XM1/a_n158_n96094# XM3/a_n100_n45563# 1.94e-20
C6805 XM1/a_n158_n80298# XM3/a_n100_n28987# 3.89e-20
C6806 XM1/a_100_n40090# XM4/w_n358_n132787# 0.049829f
C6807 XM1/a_n100_n4287# XM3/a_n158_46738# 2.85e-20
C6808 XM1/a_n158_118# XM3/a_n100_50785# 1.94e-20
C6809 XM2/a_n158_n92142# XM3/a_n100_112945# 1.45e-19
C6810 XM2/a_100_n274026# XM3/a_n158_n67222# 0.03858f
C6811 XM1/a_n100_n17211# XM3/a_n158_33270# 2.46e-20
C6812 XM2/a_n100_n279395# XM4/a_100_n72402# 2.56e-20
C6813 XM2/a_n158_n63146# XM4/w_n358_n132787# 0.105181f
C6814 XM4/w_n358_n132787# XM4/a_n100_78757# -0.004445f
C6815 XM1/a_n158_n17114# XM3/a_n100_35245# 8.22e-21
C6816 XM1/a_100_n123378# XM2/a_n158_n276662# 0.086094f
C6817 XM3/a_n100_n27951# m1_1634_n2388# 0.072015f
C6818 XM1/a_n100_132133# XM4/w_n358_n132787# 0.012279f
C6819 XM1/a_n100_n160811# XM2/a_100_n313566# 7.26e-20
C6820 XM1/a_n158_179618# XM2/a_n100_23745# 7.26e-20
C6821 XM1/a_n100_n31571# XM3/a_n158_20838# 2.85e-20
C6822 XM1/a_n158_n170766# XM2/a_n158_n324110# 4.64e-21
C6823 XM4/w_n358_n132787# XM3/a_n158_n100374# 0.032295f
C6824 XM4/a_n100_n87003# m1_1634_n2388# 0.072015f
C6825 XM2/a_n158_n226578# XM3/a_n100_n20699# 1.45e-19
C6826 XM3/a_n100_62181# m1_1634_n2388# 0.072015f
C6827 XM3/a_n100_33173# XM4/a_n100_33173# 0.009521f
C6828 XM4/w_n358_n132787# XM2/a_n100_n121235# 0.024813f
C6829 XM1/a_n100_133569# XM2/a_n158_n20970# 0.010147f
C6830 XM1/a_100_n147790# XM3/a_n158_n96230# 0.00544f
C6831 XM2/a_n100_n239855# m1_1634_n2388# 7.61e-19
C6832 XM1/a_100_n64502# XM3/a_n100_n12411# 2.85e-20
C6833 XM1/a_100_n60194# XM3/a_n158_n9206# 0.00544f
C6834 XM2/a_100_n107958# XM3/a_n100_96369# 0.005074f
C6835 XM4/w_n358_n132787# XM2/a_100_n305658# 0.1041f
C6836 XM1/a_100_n88914# XM2/a_100_n242394# 4.64e-21
C6837 XM1/a_n100_17253# XM2/a_n158_n136954# 0.010147f
C6838 XM2/a_n100_n221403# XM3/a_n158_n14386# 0.005074f
C6839 XM2/a_100_n150134# XM3/a_n100_53893# 0.005074f
C6840 XM1/a_n100_n146451# m1_1634_n2388# 9.15e-20
C6841 XM1/a_100_n139174# XM2/a_n158_n292478# 0.088042f
C6842 XM4/w_n358_n132787# XM3/a_n158_48810# 0.038462f
C6843 XM4/a_100_113042# m1_1634_n2388# 6.1e-20
C6844 XM1/a_n158_n21422# XM2/a_n100_n176591# 7.26e-20
C6845 XM1/a_100_14478# XM2/a_n158_n139590# 0.116862f
C6846 XM4/w_n358_n132787# XM4/a_n100_39389# -0.004445f
C6847 XM1/a_n158_n140610# XM3/a_n100_n90111# 1.94e-20
C6848 XM3/a_n100_n67319# m1_1634_n2388# 0.072015f
C6849 XM2/a_n158_n300386# XM3/a_n100_n96327# 7.26e-20
C6850 XM1/a_100_81970# XM2/a_100_n71054# 4.64e-21
C6851 XM1/a_100_50378# XM4/w_n358_n132787# 0.054609f
C6852 XM2/a_n100_n147595# XM3/a_n158_59170# 0.005074f
C6853 XM1/a_n100_n73215# XM2/a_n158_n226578# 0.005074f
C6854 XM4/a_n100_n126371# m1_1634_n2388# 0.072015f
C6855 XM1/a_n100_n76087# XM2/a_100_n231850# 7.26e-20
C6856 XM1/a_n100_129261# XM2/a_n158_n23606# 0.005074f
C6857 XM1/a_n100_119209# XM2/a_100_n34150# 7.26e-20
C6858 XM3/a_n100_n15519# XM4/a_n100_n15519# 0.009521f
C6859 XM1/a_100_5862# XM2/a_n100_n150231# 0.005074f
C6860 XM3/a_n100_113981# XM4/a_n100_113981# 0.009521f
C6861 XM1/a_100_44634# XM3/a_n100_96369# 2.85e-20
C6862 XM1/a_n100_n175171# XM4/w_n358_n132787# 0.01363f
C6863 XM2/a_100_n255574# XM3/a_n158_n49610# 0.077916f
C6864 XM1/a_100_123614# XM2/a_n158_n28878# 0.008981f
C6865 XM1/a_100_116434# XM2/a_100_n39422# 4.64e-21
C6866 XM1/a_n158_n18550# XM3/a_n100_33173# 1.94e-20
C6867 XM1/a_100_n166458# XM3/a_n100_n114975# 1.08e-19
C6868 XM2/a_100_n297750# XM3/a_n100_n91147# 0.005074f
C6869 XM1/a_n100_n35879# XM2/a_n158_n189674# 0.010147f
C6870 XM1/a_n158_119306# XM2/a_n158_n34150# 4.64e-21
C6871 XM1/a_100_87714# XM2/a_n100_n65879# 0.005074f
C6872 XM1/a_100_n134866# XM3/a_n158_n82762# 0.003891f
C6873 XM1/a_100_41762# XM3/a_n100_92225# 2.85e-20
C6874 XM1/a_100_n160714# XM2/a_n100_n316299# 0.005074f
C6875 XM4/w_n358_n132787# XM4/a_n100_n32095# -0.004445f
C6876 XM1/a_n100_112029# XM4/w_n358_n132787# 0.012279f
C6877 XM4/w_n358_n132787# XM2/a_n100_n245127# 0.024885f
C6878 XM3/a_n158_87142# m1_1634_n2388# 6.1e-20
C6879 XM1/a_n100_5765# XM4/w_n358_n132787# 0.013436f
C6880 XM3/a_n158_123402# m1_1634_n2388# 6.1e-20
C6881 XM4/a_100_73674# m1_1634_n2388# 6.1e-20
C6882 XM2/a_100_n136954# XM3/a_n100_68397# 0.010147f
C6883 XM1/a_n100_34485# XM3/a_n100_86009# 1.49e-19
C6884 XM2/a_n100_n147595# XM4/a_100_59170# 2.56e-20
C6885 XM3/a_n158_32234# m1_1634_n2388# 6.1e-20
C6886 XM3/a_n100_n106687# m1_1634_n2388# 0.072015f
C6887 XM2/a_100_n202854# XM3/a_n100_2093# 0.010147f
C6888 XM1/a_n100_n155067# XM2/a_n158_n310930# 0.005074f
C6889 XM1/a_n100_n57419# m1_1634_n2388# 4.56e-19
C6890 XM2/a_100_n179130# XM3/a_n100_25921# 0.010147f
C6891 XM1/a_n158_118# XM2/a_n158_n152770# 4.64e-21
C6892 XM2/a_100_n329382# XM3/a_n158_n125238# 0.014044f
C6893 XM1/a_100_113562# XM2/a_100_n42058# 4.64e-21
C6894 XM3/a_n100_n35203# XM4/a_n100_n35203# 0.009521f
C6895 XM1/a_n100_81873# XM4/w_n358_n132787# 0.012279f
C6896 XM1/a_n100_n48803# XM2/a_100_n202854# 1.45e-19
C6897 XM1/a_n100_107721# XM2/a_100_n47330# 7.26e-20
C6898 XM1/a_100_n163586# XM3/a_n158_n111770# 0.00544f
C6899 XM1/a_100_176746# XM2/a_100_23842# 4.64e-21
C6900 XM4/w_n358_n132787# XM3/a_n100_n12411# 0.009143f
C6901 XM1/a_100_112126# XM2/a_n158_n42058# 0.116862f
C6902 XM1/a_100_n11370# XM2/a_n158_n165950# 0.116862f
C6903 XM4/w_n358_n132787# XM4/a_n100_n71463# -0.004445f
C6904 XM3/a_n158_n42358# m1_1634_n2388# 6.1e-20
C6905 XM1/a_n158_66174# XM3/a_n100_118125# 1.94e-20
C6906 XM2/a_100_n113230# m1_1634_n2388# 0.017213f
C6907 XM1/a_n158_8734# XM3/a_n100_60109# 3.89e-20
C6908 XM4/w_n358_n132787# XM2/a_n158_n181766# 0.106257f
C6909 XM4/a_100_34306# m1_1634_n2388# 6.1e-20
C6910 XM2/a_100_n237122# XM3/a_n158_n31998# 0.077916f
C6911 XM1/a_n100_1457# XM3/a_n158_51918# 1.87e-20
C6912 XM1/a_n100_53153# m1_1634_n2388# 9.01e-20
C6913 XM2/a_100_n279298# XM3/a_n100_n73535# 0.010147f
C6914 XM1/a_n100_n17211# XM2/a_100_n171222# 1.45e-19
C6915 XM2/a_100_n123774# XM3/a_n100_82901# 0.005074f
C6916 XM1/a_100_n107582# XM3/a_n158_n56862# 0.004837f
C6917 XM1/a_n158_1554# XM3/a_n100_53893# 1.22e-20
C6918 XM1/a_100_15914# XM3/a_n100_67361# 4.58e-20
C6919 XM2/a_n100_n276759# XM3/a_n158_n72402# 0.005074f
C6920 XM1/a_n158_n37218# XM2/a_n158_n189674# 4.64e-21
C6921 XM1/a_100_n15678# XM2/a_n100_n168683# 0.005074f
C6922 XM4/w_n358_n132787# XM3/a_n158_121330# 0.032295f
C6923 XM1/a_n100_64641# m1_1634_n2388# 8.14e-20
C6924 XM1/a_100_n162150# XM3/a_n100_n111867# 2.35e-20
C6925 XM1/a_n100_156545# XM2/a_100_2754# 1.45e-19
C6926 XM3/a_n100_n54887# XM4/a_n100_n54887# 0.009521f
C6927 XM2/a_100_n165950# XM3/a_n100_40425# 0.005074f
C6928 XM3/a_n100_86009# XM4/a_n100_86009# 0.009521f
C6929 XM1/a_100_n4190# XM3/a_n100_47677# 2.85e-20
C6930 XM2/a_100_n92142# XM3/a_n158_114078# 0.077916f
C6931 XM4/a_n100_97405# m1_1634_n2388# 0.072015f
C6932 XM2/a_n158_n274026# XM3/a_n158_n67222# 4.64e-21
C6933 XM4/w_n358_n132787# XM3/a_n100_n51779# 0.008741f
C6934 XM4/a_100_n37178# m1_1634_n2388# 6.1e-20
C6935 XM1/a_100_n101838# XM3/a_n100_n50743# 2.85e-20
C6936 XM1/a_100_n94658# XM2/a_100_n250302# 4.64e-21
C6937 XM4/w_n358_n132787# XM4/a_n100_n110831# -0.004445f
C6938 XM3/a_n158_n81726# m1_1634_n2388# 6.1e-20
C6939 XM1/a_100_n123378# XM2/a_n100_n276759# 0.005074f
C6940 XM1/a_n100_n160811# XM2/a_n158_n313566# 0.005074f
C6941 XM3/a_n100_1057# m1_1634_n2388# 0.072015f
C6942 XM4/w_n358_n132787# XM1/a_100_178182# 0.048442f
C6943 XM1/a_n100_n51675# m1_1634_n2388# 1.29e-19
C6944 XM4/w_n358_n132787# XM4/a_n100_21# -0.004445f
C6945 XM4/w_n358_n132787# XM3/a_n100_97405# 0.009186f
C6946 XM1/a_n158_n170766# XM2/a_n100_n324207# 7.26e-20
C6947 XM1/a_n158_76226# XM2/a_n158_n78962# 4.64e-21
C6948 XM4/w_n358_n132787# XM2/a_100_n118502# 0.103341f
C6949 XM1/a_n100_n84703# XM3/a_n158_n34070# 2.85e-20
C6950 XM2/a_100_n237122# m1_1634_n2388# 0.025819f
C6951 XM4/w_n358_n132787# XM3/a_n100_42497# 0.008976f
C6952 XM2/a_n158_n107958# XM3/a_n100_96369# 7.26e-20
C6953 XM4/w_n358_n132787# XM2/a_n158_n305658# 0.101988f
C6954 XM1/a_100_n88914# XM2/a_n158_n242394# 0.105178f
C6955 XM3/a_n100_n74571# XM4/a_n100_n74571# 0.009521f
C6956 XM2/a_n100_n224039# XM4/a_100_n19566# 2.56e-20
C6957 XM2/a_100_n218670# XM3/a_n158_n14386# 0.027675f
C6958 XM2/a_n158_n150134# XM3/a_n100_53893# 7.26e-20
C6959 XM1/a_n158_n150662# XM2/a_n158_n305658# 4.64e-21
C6960 XM1/a_100_n139174# XM2/a_n100_n292575# 0.005074f
C6961 XM4/a_n100_58037# m1_1634_n2388# 0.072015f
C6962 XM4/w_n358_n132787# XM3/a_n100_n91147# 0.009084f
C6963 XM4/a_100_n76546# m1_1634_n2388# 6.1e-20
C6964 XM2/a_100_n260846# XM3/a_n100_n55923# 0.010147f
C6965 XM1/a_n100_94797# XM2/a_n158_n57874# 0.005074f
C6966 XM1/a_100_47506# XM3/a_n100_99477# 3.22e-20
C6967 XM1/a_n100_n172299# XM3/a_n158_n120058# 2.85e-20
C6968 XM1/a_n100_n96191# XM3/a_n100_n44527# 4.29e-19
C6969 XM1/a_n100_n76087# XM3/a_n158_n23710# 2.85e-20
C6970 XM2/a_n158_n15698# XM4/w_n358_n132787# 0.10321f
C6971 XM1/a_n158_57558# XM2/a_n100_n94875# 2.87e-20
C6972 XM3/a_n158_n121094# m1_1634_n2388# 6.1e-20
C6973 XM2/a_100_n144862# XM3/a_n158_59170# 0.003139f
C6974 XM1/a_100_10170# XM2/a_n100_n142323# 0.004998f
C6975 XM1/a_n100_n76087# XM2/a_n158_n231850# 0.005074f
C6976 XM1/a_100_5862# XM2/a_100_n147498# 4.64e-21
C6977 XM2/a_n158_118# XM4/w_n358_n132787# 0.103038f
C6978 XM3/a_n100_80829# m1_1634_n2388# 0.072015f
C6979 XM1/a_100_n111890# XM3/a_n100_n61103# 2.85e-20
C6980 XM2/a_n158_n297750# XM3/a_n100_n91147# 7.26e-20
C6981 XM4/w_n358_n132787# XM3/a_n158_n26818# 0.032295f
C6982 XM4/a_n100_n13447# m1_1634_n2388# 0.072015f
C6983 XM2/a_n100_n176591# m1_1634_n2388# 7.61e-19
C6984 XM3/a_n100_25921# m1_1634_n2388# 0.072015f
C6985 XM1/a_100_n160714# XM2/a_100_n313566# 4.64e-21
C6986 XM3/a_n100_n94255# XM4/a_n100_n94255# 0.009521f
C6987 XM4/w_n358_n132787# XM2/a_100_n242394# 0.105741f
C6988 XM1/a_n158_n14242# XM2/a_n158_n168586# 9.28e-21
C6989 XM1/a_n100_n117731# XM2/a_100_n271390# 1.45e-19
C6990 XM4/a_n100_18669# m1_1634_n2388# 0.072015f
C6991 XM3/a_n100_123305# m1_1634_n2388# 0.072015f
C6992 XM4/w_n358_n132787# XM3/a_n100_n130515# 0.009186f
C6993 XM4/a_100_n115914# m1_1634_n2388# 6.1e-20
C6994 XM2/a_n158_n136954# XM3/a_n100_68397# 1.45e-19
C6995 XM1/a_100_175310# XM2/a_n158_21206# 0.116862f
C6996 XM1/a_n100_54589# m1_1634_n2388# 1.07e-19
C6997 XM4/w_n358_n132787# XM3/a_n158_67458# 0.038462f
C6998 XM1/a_n100_83309# XM2/a_n158_n71054# 0.010147f
C6999 XM1/a_n100_n53111# XM2/a_100_n205490# 7.26e-20
C7000 XM1/a_100_118# XM2/a_100_n155406# 4.64e-21
C7001 XM2/a_n158_n202854# XM3/a_n100_2093# 1.45e-19
C7002 XM4/w_n358_n132787# XM3/a_n158_12550# 0.032295f
C7003 XM2/a_n158_n179130# XM3/a_n100_25921# 1.45e-19
C7004 XM1/a_n158_118# XM2/a_n100_n152867# 7.26e-20
C7005 XM4/w_n358_n132787# XM4/a_n100_112945# -0.004445f
C7006 XM2/a_n158_n329382# XM3/a_n158_n125238# 4.64e-21
C7007 XM2/a_100_n131682# XM3/a_n158_73674# 0.077916f
C7008 XM1/a_n100_n147887# XM3/a_n158_n97266# 2.85e-20
C7009 XM2/a_100_n242394# XM3/a_n100_n38311# 0.005074f
C7010 XM1/a_n100_n48803# XM2/a_n158_n202854# 0.010147f
C7011 XM1/a_n100_n173735# XM4/w_n358_n132787# 0.013471f
C7012 XM4/w_n358_n132787# XM3/a_n158_n66186# 0.032295f
C7013 XM4/a_n100_n52815# m1_1634_n2388# 0.072015f
C7014 XM2/a_100_n173858# XM3/a_n158_31198# 0.077916f
C7015 XM1/a_100_155206# XM2/a_n158_118# 0.088821f
C7016 XM1/a_n158_n8498# XM3/a_n100_42497# 1.94e-20
C7017 XM2/a_100_n326746# XM3/a_n158_n120058# 0.049874f
C7018 XM1/a_n158_n126250# XM3/a_n100_n74571# 4.81e-21
C7019 XM1/a_n158_100638# XM2/a_n158_n55238# 4.64e-21
C7020 XM2/a_n100_n332115# XM4/a_100_n125238# 2.56e-20
C7021 XM3/a_n100_n113939# XM4/a_n100_n113939# 0.009521f
C7022 XM1/a_100_n68810# XM3/a_n100_n16555# 0.001423f
C7023 XM1/a_100_n65938# XM3/a_n158_n14386# 0.00544f
C7024 XM1/a_n158_31710# XM2/a_n158_n123774# 4.64e-21
C7025 XM2/a_n100_n200315# XM4/a_100_4262# 2.56e-20
C7026 XM4/a_100_6334# m1_1634_n2388# 6.1e-20
C7027 XM4/w_n358_n132787# XM2/a_n100_n181863# 0.02519f
C7028 XM2/a_n100_n92239# XM4/a_100_112006# 2.56e-20
C7029 XM3/a_n100_53893# XM4/a_n100_53893# 0.009521f
C7030 XM2/a_n100_n300483# m1_1634_n2388# 0.001942f
C7031 XM1/a_100_1554# XM3/a_n100_52857# 5.71e-20
C7032 XM2/a_n158_n279298# XM3/a_n100_n73535# 1.45e-19
C7033 XM1/a_100_n54450# XM4/w_n358_n132787# 0.048442f
C7034 XM1/a_n158_n28602# XM3/a_n100_22813# 2.06e-20
C7035 XM1/a_n100_n17211# XM2/a_n158_n171222# 0.010147f
C7036 XM2/a_n158_n73690# XM3/a_n158_130654# 4.64e-21
C7037 XM2/a_n158_n123774# XM3/a_n100_82901# 7.26e-20
C7038 XM1/a_100_n131994# XM3/a_n100_n80787# 5.01e-19
C7039 XM1/a_100_n77426# XM3/a_n100_n26915# 2.85e-20
C7040 XM1/a_n158_n37218# XM2/a_n100_n189771# 7.26e-20
C7041 XM3/a_n158_50882# m1_1634_n2388# 6.1e-20
C7042 XM4/w_n358_n132787# XM3/a_n100_121233# 0.009186f
C7043 XM4/w_n358_n132787# XM4/a_n100_73577# -0.004445f
C7044 XM1/a_n100_n97627# XM2/a_100_n252938# 7.26e-20
C7045 XM2/a_n158_n165950# XM3/a_n100_40425# 7.26e-20
C7046 XM1/a_100_106382# XM2/a_n158_n47330# 0.116862f
C7047 XM3/a_n100_n33131# m1_1634_n2388# 0.072015f
C7048 XM2/a_100_n118502# XM3/a_n158_88178# 0.050653f
C7049 XM2/a_100_n92142# XM3/a_n100_113981# 0.010147f
C7050 XM4/w_n358_n132787# XM3/a_n158_n105554# 0.032295f
C7051 XM4/a_n100_n92183# m1_1634_n2388# 0.072015f
C7052 XM2/a_n100_n274123# XM3/a_n158_n67222# 0.005074f
C7053 XM1/a_100_97766# XM2/a_n158_n57874# 0.035075f
C7054 XM1/a_n100_n166555# XM3/a_n100_n114975# 5.67e-19
C7055 XM1/a_n158_n38654# XM3/a_n100_12453# 2.02e-20
C7056 XM1/a_n158_n104710# XM3/a_n100_n52815# 1.94e-20
C7057 XM1/a_100_n94658# XM2/a_n158_n250302# 0.034685f
C7058 XM2/a_100_n160678# XM3/a_n158_45702# 0.077916f
C7059 XM1/a_100_n86042# XM3/a_n100_n35203# 2.85e-20
C7060 XM1/a_n158_n63066# XM3/a_n100_n12411# 8.82e-21
C7061 XM4/w_n358_n132787# XM1/a_100_n162150# 0.048442f
C7062 XM1/a_n158_n134866# XM2/a_n158_n289842# 4.64e-21
C7063 XM1/a_n158_76226# XM2/a_n100_n79059# 7.26e-20
C7064 XM4/w_n358_n132787# XM2/a_n158_n118502# 0.107093f
C7065 XM1/a_n158_n177946# XM3/a_n100_n127407# 1.94e-20
C7066 XM4/a_100_107862# m1_1634_n2388# 6.1e-20
C7067 XM2/a_100_n308294# XM3/a_n158_n102446# 0.077916f
C7068 XM4/w_n358_n132787# XM2/a_n100_n305755# 0.025679f
C7069 XM4/w_n358_n132787# XM4/a_n100_34209# -0.004445f
C7070 XM1/a_100_n88914# XM2/a_n100_n242491# 0.005074f
C7071 XM2/a_n100_n31611# XM4/w_n358_n132787# 0.012195f
C7072 XM3/a_n100_n72499# m1_1634_n2388# 0.072015f
C7073 XM2/a_100_n197582# XM3/a_n100_7273# 0.010147f
C7074 XM2/a_n158_n218670# XM3/a_n158_n14386# 4.64e-21
C7075 XM1/a_100_47506# XM4/w_n358_n132787# 0.055071f
C7076 XM1/a_n158_n150662# XM2/a_n100_n305755# 7.26e-20
C7077 XM1/a_n158_13042# XM2/a_n158_n142226# 4.64e-21
C7078 XM2/a_n158_n260846# XM3/a_n100_n55923# 1.45e-19
C7079 XM1/a_n158_n21422# XM2/a_n158_n173858# 4.64e-21
C7080 XM1/a_n158_n94658# XM2/a_n158_n250302# 4.64e-21
C7081 XM1/a_100_n41526# XM4/w_n358_n132787# 0.053222f
C7082 XM1/a_100_92022# XM2/a_n100_n60607# 0.005074f
C7083 XM1/a_100_n123378# XM3/a_n100_n71463# 2.85e-20
C7084 XM1/a_100_n113326# XM3/a_n100_n62139# 5.4e-20
C7085 XM2/a_n100_n192407# XM3/a_n100_11417# 7.47e-19
C7086 XM1/a_n158_43198# XM3/a_n100_94297# 1.94e-20
C7087 XM2/a_n100_n221403# XM4/a_100_n14386# 2.56e-20
C7088 XM2/a_100_n216034# XM3/a_n158_n9206# 0.036243f
C7089 XM1/a_100_129358# XM2/a_n100_n23703# 0.005074f
C7090 XM2/a_n158_n144862# XM3/a_n158_59170# 4.64e-21
C7091 XM1/a_n158_71918# XM2/a_n158_n81598# 4.64e-21
C7092 XM1/a_100_126486# XM2/a_n100_n28975# 0.005074f
C7093 XM4/w_n358_n132787# XM4/a_n100_n37275# -0.004445f
C7094 XM1/a_n100_n83267# XM3/a_n158_n31998# 9.03e-21
C7095 XM3/a_n158_n8170# m1_1634_n2388# 6.1e-20
C7096 XM1/a_100_5862# XM2/a_n158_n147498# 0.093494f
C7097 XM4/w_n358_n132787# XM3/a_n158_118# 0.032295f
C7098 XM4/a_100_68494# m1_1634_n2388# 6.1e-20
C7099 XM1/a_100_n165022# XM3/a_n100_n112903# 2.85e-20
C7100 XM2/a_100_n173858# m1_1634_n2388# 0.025819f
C7101 XM4/w_n358_n132787# XM3/a_n100_61145# 0.008912f
C7102 XM1/a_n158_4426# XM2/a_n158_n150134# 9.28e-21
C7103 XM1/a_n100_n126347# XM3/a_n158_n74474# 2.85e-20
C7104 XM1/a_n100_n122039# XM3/a_n158_n71366# 2.85e-20
C7105 XM1/a_100_n120506# XM2/a_100_n274026# 4.64e-21
C7106 XM3/a_n100_n111867# m1_1634_n2388# 0.072015f
C7107 XM1/a_100_n160714# XM2/a_n158_n313566# 0.044032f
C7108 XM4/w_n358_n132787# XM2/a_n158_n242394# 0.101988f
C7109 XM1/a_n100_n117731# XM2/a_n158_n271390# 0.010147f
C7110 XM2/a_n100_15837# XM4/w_n358_n132787# 0.012765f
C7111 XM1/a_n100_n122039# m1_1634_n2388# 7.28e-20
C7112 XM1/a_100_n53014# XM2/a_100_n208126# 4.64e-21
C7113 XM2/a_n100_n73787# m1_1634_n2388# 3.8e-19
C7114 XM2/a_100_n289842# XM3/a_n158_n84834# 0.077916f
C7115 XM1/a_n100_n53111# XM2/a_n158_n205490# 0.005074f
C7116 XM4/a_n100_131593# m1_1634_n2388# 0.036019f
C7117 XM1/a_100_n180818# XM3/a_n100_n130515# 2.85e-20
C7118 XM1/a_100_n119070# XM3/a_n100_n67319# 2.85e-20
C7119 XM1/a_100_118# XM2/a_n158_n155406# 0.046369f
C7120 XM1/a_100_38890# XM3/a_n100_91189# 2.85e-20
C7121 XM2/a_100_n332018# XM3/a_n100_n126371# 0.010147f
C7122 XM1/a_100_n152098# XM4/w_n358_n132787# 0.049669f
C7123 XM4/w_n358_n132787# XM3/a_n100_n17591# 0.010106f
C7124 XM4/a_100_n2990# m1_1634_n2388# 6.1e-20
C7125 XM1/a_n100_n155067# XM2/a_100_n308294# 7.26e-20
C7126 XM2/a_n100_n329479# XM3/a_n158_n125238# 0.005074f
C7127 XM4/w_n358_n132787# XM4/a_n100_n76643# -0.004445f
C7128 XM3/a_n158_n47538# m1_1634_n2388# 6.1e-20
C7129 XM2/a_n158_n242394# XM3/a_n100_n38311# 7.26e-20
C7130 XM3/a_n100_21777# XM4/a_n100_21777# 0.009521f
C7131 XM4/a_100_29126# m1_1634_n2388# 6.1e-20
C7132 XM1/a_n100_n83267# m1_1634_n2388# 8.34e-20
C7133 XM2/a_100_n15698# XM1/a_n100_137877# 1.3e-19
C7134 XM3/a_n100_99477# m1_1634_n2388# 0.072015f
C7135 XM2/a_n158_n326746# XM3/a_n158_n120058# 4.64e-21
C7136 XM1/a_n100_n47367# XM4/w_n358_n132787# 0.013548f
C7137 XM1/a_n100_n146451# XM2/a_100_n300386# 1.45e-19
C7138 XM2/a_n100_n113327# m1_1634_n2388# 7.61e-19
C7139 XM1/a_n158_31710# XM2/a_n100_n123871# 7.26e-20
C7140 XM2/a_100_n239758# XM3/a_n100_n33131# 0.005074f
C7141 XM3/a_n100_44569# m1_1634_n2388# 0.072015f
C7142 XM1/a_100_110690# XM2/a_100_n44694# 4.64e-21
C7143 XM4/w_n358_n132787# XM2/a_100_n179130# 0.106377f
C7144 XM1/a_n158_155206# XM2/a_n100_21# 7.26e-20
C7145 XM2/a_100_n297750# m1_1634_n2388# 0.017213f
C7146 XM1/a_n158_70482# XM3/a_n100_122269# 1.94e-20
C7147 XM1/a_n158_109254# XM2/a_n158_n44694# 9.28e-21
C7148 XM2/a_n158_n73690# XM3/a_n100_130557# 7.26e-20
C7149 XM1/a_100_n27166# XM4/w_n358_n132787# 0.048442f
C7150 XM4/a_n100_92225# m1_1634_n2388# 0.072015f
C7151 XM4/w_n358_n132787# XM3/a_n158_86106# 0.037178f
C7152 XM4/w_n358_n132787# XM3/a_n100_n56959# 0.008831f
C7153 XM4/a_100_n42358# m1_1634_n2388# 6.1e-20
C7154 XM2/a_n100_n89603# XM4/a_100_117186# 2.56e-20
C7155 XM1/a_n158_7298# XM3/a_n100_59073# 1.94e-20
C7156 XM1/a_n100_n97627# XM2/a_n158_n252938# 0.005074f
C7157 XM1/a_n158_n88914# XM3/a_n158_n38214# 1.14e-21
C7158 XM2/a_n100_n166047# XM3/a_n100_40425# 0.001011f
C7159 XM4/w_n358_n132787# XM4/a_n100_n116011# -0.004445f
C7160 XM3/a_n158_n86906# m1_1634_n2388# 6.1e-20
C7161 XM4/w_n358_n132787# XM3/a_n158_31198# 0.032295f
C7162 XM2/a_n158_n118502# XM3/a_n158_88178# 4.64e-21
C7163 XM2/a_n158_n92142# XM3/a_n100_113981# 1.45e-19
C7164 XM2/a_100_n271390# XM3/a_n158_n67222# 0.016381f
C7165 XM2/a_n100_n276759# XM4/a_100_n72402# 2.56e-20
C7166 XM3/a_n100_2093# XM4/a_n100_2093# 0.009521f
C7167 XM1/a_100_n15678# XM3/a_n158_35342# 0.003891f
C7168 XM1/a_n158_61866# XM3/a_n100_112945# 1.94e-20
C7169 XM2/a_100_n313566# XM3/a_n100_n108759# 0.010147f
C7170 XM1/a_100_n94658# XM2/a_n100_n250399# 0.005074f
C7171 XM4/w_n358_n132787# XM3/a_n100_6237# 0.008456f
C7172 XM1/a_100_n35782# XM4/w_n358_n132787# 0.048442f
C7173 XM1/a_100_160950# XM2/a_100_5390# 4.64e-21
C7174 XM1/a_100_n116198# XM3/a_n158_n64114# 0.003891f
C7175 XM1/a_n100_n106243# XM3/a_n158_n55826# 5.8e-21
C7176 XM1/a_n158_n44398# XM2/a_n158_n200218# 4.64e-21
C7177 XM1/a_n158_n30038# XM3/a_n100_20741# 1.94e-20
C7178 XM1/a_n158_n134866# XM2/a_n100_n289939# 7.26e-20
C7179 XM1/a_100_n73118# XM3/a_n158_n22674# 0.001666f
C7180 XM2/a_100_n202854# XM3/a_n158_3226# 0.077916f
C7181 XM4/w_n358_n132787# XM2/a_n100_n118599# 0.025738f
C7182 XM2/a_n100_n237219# m1_1634_n2388# 7.61e-19
C7183 XM4/a_n100_52857# m1_1634_n2388# 0.072015f
C7184 XM1/a_100_23094# XM2/a_n158_n131682# 0.116862f
C7185 XM4/w_n358_n132787# XM3/a_n100_n96327# 0.009004f
C7186 XM4/a_100_n81726# m1_1634_n2388# 6.1e-20
C7187 XM4/w_n358_n132787# XM4/a_n100_6237# -0.004445f
C7188 XM1/a_n100_97669# XM2/a_n158_n57874# 0.005074f
C7189 XM4/w_n358_n132787# XM2/a_100_n303022# 0.103341f
C7190 XM2/a_100_n221306# XM3/a_n100_n15519# 0.010147f
C7191 XM2/a_n158_n197582# XM3/a_n100_7273# 1.45e-19
C7192 XM3/a_n158_69530# m1_1634_n2388# 6.1e-20
C7193 XM3/a_n158_n126274# m1_1634_n2388# 6.1e-20
C7194 XM1/a_n100_n101935# XM3/a_n100_n50743# 0.001106f
C7195 XM1/a_n100_152237# XM2/a_n158_n2518# 0.005074f
C7196 XM2/a_n100_n218767# XM3/a_n158_n14386# 0.005074f
C7197 XM1/a_n158_13042# XM2/a_n100_n142323# 7.26e-20
C7198 XM3/a_n158_14622# m1_1634_n2388# 6.1e-20
C7199 XM1/a_n158_n21422# XM2/a_n100_n173955# 7.26e-20
C7200 XM1/a_n100_94797# XM4/w_n358_n132787# 0.012279f
C7201 XM1/a_n158_n94658# XM2/a_n100_n250399# 7.26e-20
C7202 XM1/a_n100_n163683# XM3/a_n158_n112806# 2.85e-20
C7203 XM4/w_n358_n132787# XM3/a_n158_n31998# 0.032295f
C7204 XM4/a_n100_n18627# m1_1634_n2388# 0.072015f
C7205 XM2/a_n158_n216034# XM3/a_n158_n9206# 4.64e-21
C7206 XM1/a_n158_71918# XM2/a_n100_n81695# 6.58e-20
C7207 XM2/a_n100_n144959# XM3/a_n158_59170# 0.005074f
C7208 XM1/a_n158_n100402# XM3/a_n100_n49707# 1.94e-20
C7209 XM1/a_n100_n76087# XM2/a_100_n229214# 7.26e-20
C7210 XM1/a_n100_44537# XM3/a_n158_96466# 2.85e-20
C7211 XM1/a_100_5862# XM2/a_n100_n147595# 0.005074f
C7212 XM4/a_n100_13489# m1_1634_n2388# 0.072015f
C7213 XM4/a_100_n121094# m1_1634_n2388# 6.1e-20
C7214 XM2/a_100_n295114# XM3/a_n100_n91147# 0.005074f
C7215 XM1/a_100_n120506# XM2/a_n158_n274026# 0.109073f
C7216 XM1/a_100_84842# XM2/a_n158_n71054# 0.010149f
C7217 XM1/a_100_n160714# XM2/a_n100_n313663# 0.005074f
C7218 XM4/w_n358_n132787# XM2/a_n100_n242491# 0.024273f
C7219 XM3/a_n158_124438# m1_1634_n2388# 6.1e-20
C7220 XM4/w_n358_n132787# XM4/a_n100_107765# -0.004445f
C7221 XM1/a_100_n53014# XM2/a_n158_n208126# 0.086484f
C7222 XM3/a_n100_74613# XM4/a_n100_74613# 0.009521f
C7223 XM3/a_n158_2190# m1_1634_n2388# 6.1e-20
C7224 XM1/a_n158_n34346# XM3/a_n100_16597# 6.41e-21
C7225 XM1/a_100_113562# XM4/w_n358_n132787# 0.053546f
C7226 XM2/a_n100_n144959# XM4/a_100_59170# 2.56e-20
C7227 XM1/a_100_118# XM2/a_n100_n155503# 0.005074f
C7228 XM2/a_n100_n18431# XM1/a_n100_136441# 6.96e-19
C7229 XM2/a_100_n18334# XM1/a_100_136538# 4.64e-21
C7230 XM2/a_n158_n18334# XM1/a_n158_136538# 4.64e-21
C7231 XM2/a_n100_n21067# XM1/a_n100_135005# 0.003206f
C7232 XM2/a_n158_n332018# XM3/a_n100_n126371# 1.45e-19
C7233 XM4/w_n358_n132787# XM3/a_n158_n71366# 0.032295f
C7234 XM4/a_n100_n57995# m1_1634_n2388# 0.072015f
C7235 XM1/a_n100_n155067# XM2/a_n158_n308294# 0.005074f
C7236 XM1/a_100_n96094# XM3/a_n100_n45563# 2.85e-20
C7237 XM1/a_100_n54450# XM3/a_n100_n4123# 2.85e-20
C7238 XM4/w_n358_n132787# m1_1634_n2388# 30.779135f
C7239 XM1/a_n100_20125# XM3/a_n100_70469# 7.28e-19
C7240 XM1/a_100_25966# XM3/a_n158_77818# 0.004535f
C7241 XM1/a_n100_76129# XM3/a_n100_126413# 6.89e-19
C7242 XM2/a_n100_n326843# XM3/a_n158_n120058# 0.005074f
C7243 XM1/a_n100_n146451# XM2/a_n158_n300386# 0.010147f
C7244 XM2/a_100_n110594# m1_1634_n2388# 0.023368f
C7245 XM4/w_n358_n132787# XM3/a_n100_79793# 0.008905f
C7246 XM2/a_n158_n239758# XM3/a_n100_n33131# 7.26e-20
C7247 XM4/w_n358_n132787# XM2/a_n158_n179130# 0.101988f
C7248 XM4/w_n358_n132787# XM4/a_n100_68397# -0.004445f
C7249 XM1/a_n158_n97530# XM3/a_n100_n45563# 7.21e-21
C7250 XM1/a_n158_n28602# XM2/a_n158_n184402# 4.64e-21
C7251 XM3/a_n100_n38311# m1_1634_n2388# 0.072015f
C7252 XM1/a_100_n61630# XM3/a_n100_n11375# 1.52e-20
C7253 XM4/w_n358_n132787# XM3/a_n100_24885# 0.009186f
C7254 XM1/a_100_76226# XM3/a_n158_127546# 0.002344f
C7255 XM2/a_100_n121138# XM3/a_n100_82901# 0.005074f
C7256 XM1/a_100_n9934# XM3/a_n158_40522# 9.46e-19
C7257 XM1/a_100_2990# XM3/a_n158_53990# 0.00544f
C7258 XM4/w_n358_n132787# XM3/a_n158_122366# 0.03804f
C7259 XM4/w_n358_n132787# XM3/a_n158_n110734# 0.032295f
C7260 XM4/a_n100_n97363# m1_1634_n2388# 0.072015f
C7261 XM1/a_100_n129122# XM3/a_n158_n77582# 0.00544f
C7262 XM1/a_n100_169469# XM4/w_n358_n132787# 0.012074f
C7263 XM1/a_n158_158078# XM2/a_n100_2657# 7.26e-20
C7264 XM1/a_n100_n4287# XM3/a_n158_47774# 2.85e-20
C7265 XM1/a_n158_118# XM3/a_n100_51821# 5.41e-21
C7266 XM2/a_n100_n118599# XM3/a_n158_88178# 0.005074f
C7267 XM1/a_n100_n21519# m1_1634_n2388# 7.42e-20
C7268 XM2/a_n158_n271390# XM3/a_n158_n67222# 4.64e-21
C7269 XM1/a_n158_n67374# XM2/a_n158_n221306# 9.28e-21
C7270 XM4/w_n358_n132787# XM4/a_n100_n3087# -0.004445f
C7271 XM1/a_100_103510# XM2/a_100_n49966# 4.64e-21
C7272 XM2/a_n158_n60510# XM4/w_n358_n132787# 0.107093f
C7273 XM1/a_100_97766# XM4/w_n358_n132787# 0.053546f
C7274 XM2/a_n158_n313566# XM3/a_n100_n108759# 1.45e-19
C7275 XM1/a_100_n94658# XM2/a_100_n247666# 4.64e-21
C7276 XM1/a_100_n17114# XM4/w_n358_n132787# 0.048442f
C7277 XM4/a_100_102682# m1_1634_n2388# 6.1e-20
C7278 XM1/a_n158_n175074# XM3/a_n100_n124299# 1.94e-20
C7279 XM1/a_n100_n40187# XM4/w_n358_n132787# 0.015149f
C7280 XM1/a_n158_179618# XM2/a_n100_26381# 7.26e-20
C7281 XM1/a_n158_n103274# XM2/a_n158_n258210# 4.64e-21
C7282 XM1/a_n158_n44398# XM2/a_n100_n200315# 7.26e-20
C7283 XM4/w_n358_n132787# XM4/a_n100_29029# -0.004445f
C7284 XM1/a_n100_4329# m1_1634_n2388# 8.88e-20
C7285 XM2/a_n100_n274123# XM4/a_100_n67222# 2.56e-20
C7286 XM2/a_100_n268754# XM3/a_n158_n62042# 0.047538f
C7287 XM1/a_n158_76226# XM2/a_n158_n76326# 4.64e-21
C7288 XM3/a_n100_63217# m1_1634_n2388# 0.072015f
C7289 XM3/a_n100_n77679# m1_1634_n2388# 0.072015f
C7290 XM4/w_n358_n132787# XM2/a_100_n115866# 0.10657f
C7291 XM1/a_100_51814# XM4/w_n358_n132787# 0.048442f
C7292 XM2/a_100_n234486# m1_1634_n2388# 0.017213f
C7293 XM1/a_n100_n169427# XM4/w_n358_n132787# 0.012382f
C7294 XM1/a_n158_n27166# XM3/a_n100_23849# 1.94e-20
C7295 XM2/a_100_n107958# XM3/a_n100_97405# 0.010147f
C7296 XM4/w_n358_n132787# XM2/a_n158_n303022# 0.106161f
C7297 XM3/a_n100_n20699# XM4/a_n100_n20699# 0.009521f
C7298 XM1/a_n100_67513# XM4/w_n358_n132787# 0.013474f
C7299 XM2/a_n158_n221306# XM3/a_n100_n15519# 1.45e-19
C7300 XM1/a_100_94894# XM2/a_n100_n60607# 0.005074f
C7301 XM1/a_n100_n34443# XM3/a_n158_16694# 2.85e-20
C7302 XM2/a_100_n150134# XM3/a_n100_54929# 0.010147f
C7303 XM1/a_100_n160714# XM3/a_n100_n109795# 3.44e-19
C7304 XM1/a_100_n150662# XM3/a_n158_n98302# 3.95e-20
C7305 XM4/w_n358_n132787# XM3/a_n158_49846# 0.032295f
C7306 XM4/w_n358_n132787# XM4/a_n100_n42455# -0.004445f
C7307 XM3/a_n158_n13350# m1_1634_n2388# 6.1e-20
C7308 XM1/a_n158_n129122# XM2/a_n158_n284570# 4.64e-21
C7309 XM2/a_100_n192310# XM3/a_n100_12453# 0.007586f
C7310 XM1/a_n100_n173735# XM3/a_n100_n122227# 3.25e-20
C7311 XM2/a_n100_n216131# XM3/a_n158_n9206# 0.005074f
C7312 XM4/a_100_63314# m1_1634_n2388# 6.1e-20
C7313 XM1/a_n158_n123378# XM3/a_n100_n72499# 1.94e-20
C7314 XM1/a_n100_n76087# XM2/a_n158_n229214# 0.005074f
C7315 XM1/a_n100_172341# XM4/w_n358_n132787# 0.012279f
C7316 XM1/a_n100_80437# XM2/a_100_n73690# 1.45e-19
C7317 XM3/a_n100_n117047# m1_1634_n2388# 0.072015f
C7318 XM3/a_n100_42497# XM4/a_n100_42497# 0.009521f
C7319 XM1/a_100_116434# XM2/a_100_n36786# 4.64e-21
C7320 XM1/a_100_n143482# XM3/a_n100_n92183# 5.71e-20
C7321 XM2/a_n158_n295114# XM3/a_n100_n91147# 7.26e-20
C7322 XM1/a_100_n32910# XM2/a_n158_n187038# 0.116862f
C7323 XM3/a_n100_n40383# XM4/a_n100_n40383# 0.009521f
C7324 XM2/a_n100_n173955# m1_1634_n2388# 7.61e-19
C7325 XM1/a_100_41762# XM3/a_n100_93261# 2.85e-20
C7326 XM1/a_100_n120506# XM2/a_n100_n274123# 0.004269f
C7327 XM4/a_n100_126413# m1_1634_n2388# 0.072015f
C7328 XM1/a_100_n157842# XM2/a_100_n313566# 4.64e-21
C7329 XM1/a_n158_n98966# XM3/a_n100_n48671# 1.78e-20
C7330 XM4/w_n358_n132787# XM2/a_100_n239758# 0.103341f
C7331 XM2/a_100_n250302# XM3/a_n158_n44430# 0.077916f
C7332 XM4/w_n358_n132787# XM3/a_n100_n22771# 0.008054f
C7333 XM4/a_100_n8170# m1_1634_n2388# 6.1e-20
C7334 XM3/a_n158_88178# m1_1634_n2388# 6.1e-20
C7335 XM1/a_n100_146493# XM2/a_100_n7790# 1.45e-19
C7336 XM3/a_n100_124341# m1_1634_n2388# 0.072015f
C7337 XM1/a_n158_n176510# XM2/a_n158_n332018# 4.64e-21
C7338 XM2/a_100_n292478# XM3/a_n100_n85967# 0.005074f
C7339 XM1/a_n100_n68907# XM3/a_n158_n16458# 2.85e-20
C7340 XM1/a_100_n53014# XM2/a_n100_n208223# 0.005074f
C7341 XM2/a_100_n136954# XM3/a_n100_69433# 0.005074f
C7342 XM4/w_n358_n132787# XM4/a_n100_n81823# -0.004445f
C7343 XM3/a_n158_n52718# m1_1634_n2388# 6.1e-20
C7344 XM1/a_n100_34485# XM3/a_n100_87045# 4.42e-19
C7345 XM3/a_n158_33270# m1_1634_n2388# 6.1e-20
C7346 XM1/a_n158_n147790# XM3/a_n100_n96327# 2.75e-20
C7347 XM4/a_100_23946# m1_1634_n2388# 6.1e-20
C7348 XM1/a_100_118# XM2/a_100_n152770# 4.64e-21
C7349 XM3/a_n100_121233# XM4/a_n100_121233# 0.009521f
C7350 XM1/a_n158_34582# XM3/a_n100_84973# 1.94e-20
C7351 XM2/a_100_n179130# XM3/a_n100_26957# 0.010147f
C7352 XM1/a_100_n175074# XM3/a_n100_n124299# 2.85e-20
C7353 XM1/a_100_113562# XM2/a_100_n39422# 4.64e-21
C7354 XM1/a_n158_30274# XM3/a_n100_80829# 1.94e-20
C7355 XM2/a_n100_n142323# XM4/a_100_64350# 2.56e-20
C7356 XM1/a_n100_107721# XM2/a_100_n44694# 7.26e-20
C7357 XM2/a_100_n197582# XM3/a_n158_8406# 0.077916f
C7358 iout_n iout 0.028696f
C7359 XM1/a_n100_60333# XM3/a_n158_110970# 2.85e-20
C7360 XM1/a_n100_8637# XM3/a_n158_59170# 3.31e-19
C7361 XM3/a_n100_n60067# XM4/a_n100_n60067# 0.009521f
C7362 XM1/a_n100_n7159# XM4/w_n358_n132787# 0.012504f
C7363 XM1/a_n100_103413# XM4/w_n358_n132787# 0.012081f
C7364 XM2/a_100_n324110# XM3/a_n158_n120058# 0.005086f
C7365 XM1/a_n158_n142046# XM2/a_n158_n297750# 4.64e-21
C7366 XM1/a_n158_57558# XM3/a_n100_107765# 2e-22
C7367 XM4/a_n100_87045# m1_1634_n2388# 0.072015f
C7368 XM2/a_n100_n329479# XM4/a_100_n125238# 2.56e-20
C7369 XM1/a_100_173874# XM2/a_n100_18473# 0.005074f
C7370 XM1/a_n158_31710# XM2/a_n158_n121138# 4.64e-21
C7371 XM4/w_n358_n132787# XM3/a_n100_n62139# 0.009144f
C7372 XM1/a_n158_n100402# XM2/a_n158_n255574# 4.64e-21
C7373 XM4/a_100_n47538# m1_1634_n2388# 6.1e-20
C7374 XM4/w_n358_n132787# XM2/a_n100_n179227# 0.025223f
C7375 XM1/a_n100_n99063# XM2/a_100_n252938# 1.45e-19
C7376 XM1/a_n158_n28602# XM2/a_n100_n184499# 7.26e-20
C7377 XM4/w_n358_n132787# XM4/a_n100_n121191# -0.004445f
C7378 XM3/a_n158_n92086# m1_1634_n2388# 6.1e-20
C7379 XM2/a_n100_n297847# m1_1634_n2388# 7.61e-19
C7380 XM1/a_100_76226# XM3/a_n100_127449# 2.45e-19
C7381 XM1/a_n158_n83170# XM2/a_n158_n237122# 9.28e-21
C7382 XM2/a_n158_n121138# XM3/a_n100_82901# 7.26e-20
C7383 XM4/w_n358_n132787# XM3/a_n100_122269# 0.008387f
C7384 XM1/a_100_50378# XM3/a_n158_101646# 0.00544f
C7385 XM1/a_n100_n97627# XM2/a_100_n250302# 7.26e-20
C7386 XM2/a_100_n231850# XM3/a_n158_n26818# 0.077916f
C7387 XM1/a_n100_n28699# XM3/a_n158_21874# 2.85e-20
C7388 XM1/a_100_118# XM3/a_n100_50785# 2.85e-20
C7389 XM1/a_100_n97530# XM3/a_n100_n45563# 0.001324f
C7390 XM1/a_n100_n77523# XM3/a_n158_n25782# 1.37e-20
C7391 XM2/a_100_n274026# XM3/a_n100_n68355# 0.010147f
C7392 XM2/a_100_n115866# XM3/a_n158_88178# 0.004307f
C7393 XM2/a_100_n92142# XM3/a_n100_115017# 0.002941f
C7394 XM2/a_n100_n271487# XM3/a_n158_n67222# 0.005074f
C7395 XM1/a_n100_n67471# XM3/a_n158_n16458# 2.85e-20
C7396 XM3/a_n100_n79751# XM4/a_n100_n79751# 0.009521f
C7397 XM1/a_100_n94658# XM2/a_n158_n247666# 0.059221f
C7398 XM4/a_n100_47677# m1_1634_n2388# 0.072015f
C7399 XM4/w_n358_n132787# XM3/a_n100_n101507# 0.009186f
C7400 XM4/a_100_n86906# m1_1634_n2388# 6.1e-20
C7401 XM1/a_n158_n103274# XM2/a_n100_n258307# 7.26e-20
C7402 XM4/w_n358_n132787# XM3/a_n100_98441# 0.008464f
C7403 XM3/a_n100_104657# XM4/a_n100_104657# 0.009521f
C7404 XM1/a_n100_n120603# XM4/w_n358_n132787# 0.013776f
C7405 XM2/a_n158_n268754# XM3/a_n158_n62042# 4.64e-21
C7406 XM1/a_n158_76226# XM2/a_n100_n76423# 7.26e-20
C7407 XM3/a_n158_n131454# m1_1634_n2388# 6.1e-20
C7408 XM1/a_100_n147790# XM3/a_n100_n97363# 2.85e-20
C7409 XM4/w_n358_n132787# XM2/a_n158_n115866# 0.10297f
C7410 XM1/a_n158_n27166# XM2/a_n158_n181766# 9.28e-21
C7411 XM4/w_n358_n132787# XM3/a_n100_43533# 0.009186f
C7412 XM2/a_n158_n107958# XM3/a_n100_97405# 1.45e-19
C7413 XM4/w_n358_n132787# XM2/a_n100_n303119# 0.024812f
C7414 XM1/a_n100_97669# XM4/w_n358_n132787# 0.012279f
C7415 XM1/a_n158_n60194# XM2/a_n158_n216034# 4.64e-21
C7416 XM1/a_n100_159417# XM2/a_100_5390# 1.45e-19
C7417 XM1/a_n100_n142143# XM3/a_n158_n90014# 2.85e-20
C7418 XM1/a_100_169566# XM2/a_n158_15934# 0.116862f
C7419 XM3/a_n158_100610# m1_1634_n2388# 6.1e-20
C7420 XM4/w_n358_n132787# XM3/a_n158_n37178# 0.032295f
C7421 XM4/a_n100_n23807# m1_1634_n2388# 0.072015f
C7422 XM2/a_n158_n150134# XM3/a_n100_54929# 1.45e-19
C7423 XM1/a_n158_n150662# XM2/a_n100_n303119# 4.26e-20
C7424 XM1/a_n100_21# m1_1634_n2388# 1.3e-19
C7425 XM1/a_100_168130# XM2/a_n100_13201# 6.5e-19
C7426 XM1/a_n158_13042# XM2/a_n158_n139590# 4.64e-21
C7427 XM1/a_100_n121942# XM2/a_n158_n276662# 0.116862f
C7428 XM3/a_n100_10381# XM4/a_n100_10381# 0.009521f
C7429 XM1/a_100_n30038# XM2/a_n158_n184402# 0.116862f
C7430 XM1/a_100_89150# XM2/a_100_n65782# 4.64e-21
C7431 XM3/a_n100_95333# XM4/a_n100_95333# 0.009521f
C7432 XM1/a_100_n167894# XM3/a_n158_n116950# 7.57e-19
C7433 XM3/a_n100_n99435# XM4/a_n100_n99435# 0.009521f
C7434 XM1/a_n158_n129122# XM2/a_n100_n284667# 7.26e-20
C7435 XM1/a_n158_n94658# XM2/a_n158_n247666# 4.64e-21
C7436 XM2/a_n158_n192310# XM3/a_n100_12453# 1.21e-19
C7437 XM2/a_n158_n13062# XM4/w_n358_n132787# 0.107093f
C7438 XM2/a_100_n213398# XM3/a_n158_n9206# 0.018717f
C7439 XM1/a_n100_n55983# m1_1634_n2388# 1.07e-19
C7440 XM1/a_n158_155206# XM2/a_n158_2754# 4.64e-21
C7441 XM1/a_100_47506# XM2/a_100_n107958# 4.64e-21
C7442 XM4/a_100_n126274# m1_1634_n2388# 6.1e-20
C7443 XM2/a_n100_n218767# XM4/a_100_n14386# 2.56e-20
C7444 XM2/a_100_n144862# XM3/a_n158_60206# 0.077916f
C7445 XM1/a_100_166694# XM2/a_n158_13298# 0.096999f
C7446 XM1/a_n158_149462# XM2/a_n158_n5154# 9.28e-21
C7447 XM2/a_100_n255574# XM3/a_n100_n50743# 0.010147f
C7448 XM1/a_n158_126486# XM2/a_n158_n28878# 4.64e-21
C7449 XM2/a_100_n187038# XM3/a_n158_17730# 0.0748f
C7450 XM1/a_n100_61769# XM2/a_100_n92142# 1.45e-19
C7451 XM3/a_n100_81865# m1_1634_n2388# 0.072014f
C7452 XM1/a_100_n134866# XM3/a_n100_n83895# 2.85e-20
C7453 XM1/a_n100_n60291# m1_1634_n2388# 1.3e-19
C7454 XM4/w_n358_n132787# XM4/a_n100_102585# -0.004445f
C7455 XM1/a_100_n57322# XM3/a_n100_n5159# 2.85e-20
C7456 XM2/a_100_n171222# m1_1634_n2388# 0.017213f
C7457 XM3/a_n100_n4123# m1_1634_n2388# 0.072015f
C7458 XM1/a_n100_80437# XM3/a_n158_131690# 1.37e-20
C7459 XM1/a_100_n157842# XM2/a_n158_n313566# 0.026896f
C7460 XM3/a_n100_26957# m1_1634_n2388# 0.072015f
C7461 XM1/a_n158_37454# XM3/a_n100_88081# 1.94e-20
C7462 XM4/w_n358_n132787# XM2/a_n158_n239758# 0.104449f
C7463 XM4/w_n358_n132787# XM3/a_n158_n76546# 0.032295f
C7464 XM4/a_n100_n63175# m1_1634_n2388# 0.072015f
C7465 XM1/a_100_n22858# XM2/a_n158_n176494# 0.116862f
C7466 XM4/w_n358_n132787# XM3/a_n158_7370# 0.032295f
C7467 XM1/a_n158_n176510# XM2/a_n100_n332115# 7.26e-20
C7468 XM2/a_n158_n292478# XM3/a_n100_n85967# 7.26e-20
C7469 XM1/a_n100_n94755# XM3/a_n100_n44527# 2.08e-19
C7470 XM1/a_100_n78862# XM3/a_n100_n26915# 2.85e-20
C7471 XM1/a_n158_n65938# XM3/a_n100_n15519# 1.94e-20
C7472 XM1/a_100_n53014# XM2/a_100_n205490# 4.64e-21
C7473 XM4/w_n358_n132787# XM3/a_n158_68494# 0.032295f
C7474 XM2/a_n158_n136954# XM3/a_n100_69433# 7.26e-20
C7475 XM3/a_n100_n119119# XM4/a_n100_n119119# 0.009521f
C7476 XM2/a_n100_n189771# XM4/a_n100_16597# 1.28e-20
C7477 XM1/a_n158_n139174# XM2/a_n158_n295114# 4.64e-21
C7478 XM1/a_100_118# XM2/a_n158_n152770# 0.047538f
C7479 XM2/a_n158_29114# XM1/a_100_182490# 0.095052f
C7480 XM2/a_n100_26381# XM1/a_n100_182393# 3.73e-19
C7481 XM1/a_n158_n147790# XM2/a_n158_n303022# 4.64e-21
C7482 XM2/a_n158_n179130# XM3/a_n100_26957# 1.45e-19
C7483 XM1/a_100_80534# XM2/a_n158_n73690# 0.116862f
C7484 XM4/w_n358_n132787# XM3/a_n158_13586# 0.032295f
C7485 XM1/a_n100_n8595# XM4/w_n358_n132787# 0.012618f
C7486 XM1/a_100_n163586# XM3/a_n100_n112903# 2.85e-20
C7487 XM1/a_n158_n153534# XM3/a_n100_n101507# 1.94e-20
C7488 XM1/a_100_156642# XM4/w_n358_n132787# 0.048442f
C7489 XM2/a_100_n131682# XM3/a_n158_74710# 0.077916f
C7490 XM1/a_n100_22997# XM3/a_n158_73674# 2.85e-20
C7491 XM1/a_n158_n180818# XM3/a_n100_n129479# 3.89e-20
C7492 XM1/a_n100_n124911# XM3/a_n158_n72402# 2.58e-20
C7493 XM4/w_n358_n132787# XM4/a_n100_63217# -0.004445f
C7494 XM2/a_100_n173858# XM3/a_n158_32234# 0.077916f
C7495 XM1/a_n100_n12903# XM3/a_n158_39486# 2.85e-20
C7496 XM1/a_n158_n8498# XM3/a_n100_43533# 1.94e-20
C7497 XM1/a_n158_107818# XM2/a_n158_n47330# 4.64e-21
C7498 XM1/a_n100_n157939# XM2/a_100_n313566# 7.26e-20
C7499 XM3/a_n100_n43491# m1_1634_n2388# 0.072015f
C7500 XM2/a_n158_n324110# XM3/a_n158_n120058# 4.64e-21
C7501 XM1/a_n158_n142046# XM2/a_n100_n297847# 7.26e-20
C7502 XM1/a_n158_100638# XM2/a_n158_n52602# 4.64e-21
C7503 XM2/a_n100_n110691# m1_1634_n2388# 0.001261f
C7504 XM1/a_n100_33049# XM4/w_n358_n132787# 0.01363f
C7505 XM2/a_100_n237122# XM3/a_n100_n33131# 0.005074f
C7506 XM1/a_n158_31710# XM2/a_n100_n121235# 7.26e-20
C7507 XM4/w_n358_n132787# XM3/a_n158_n115914# 0.032295f
C7508 XM4/a_n100_n102543# m1_1634_n2388# 0.072015f
C7509 XM1/a_n158_n100402# XM2/a_n100_n255671# 7.26e-20
C7510 XM4/w_n358_n132787# XM2/a_100_n176494# 0.103341f
C7511 XM1/a_n100_n176607# XM3/a_n158_n124202# 2.85e-20
C7512 XM1/a_n100_n137835# m1_1634_n2388# 1.05e-19
C7513 XM1/a_n100_n99063# XM2/a_n158_n252938# 0.010147f
C7514 XM1/a_100_1554# XM3/a_n100_53893# 1.87e-20
C7515 XM2/a_100_n295114# m1_1634_n2388# 0.025819f
C7516 XM2/a_100_n321474# XM3/a_n158_n114878# 0.058832f
C7517 XM1/a_n100_109157# XM2/a_100_n44694# 1.45e-19
C7518 XM2/a_n158_n73690# XM3/a_n100_131593# 1.45e-19
C7519 XM2/a_n100_n326843# XM4/a_100_n120058# 2.56e-20
C7520 XM1/a_100_50378# XM3/a_n100_101549# 4.93e-20
C7521 XM4/w_n358_n132787# XM1/a_100_n133430# 0.048442f
C7522 XM4/w_n358_n132787# XM4/a_n100_n8267# -0.004445f
C7523 XM1/a_n158_n1318# XM3/a_n100_49749# 1.94e-20
C7524 XM3/a_n158_51918# m1_1634_n2388# 6.1e-20
C7525 XM2/a_n100_n86967# XM4/a_100_117186# 2.56e-20
C7526 XM1/a_n100_n97627# XM2/a_n158_n250302# 0.005074f
C7527 XM2/a_n100_n163411# XM3/a_n100_40425# 0.001628f
C7528 XM4/a_100_97502# m1_1634_n2388# 6.1e-20
C7529 XM1/a_100_n119070# XM4/w_n358_n132787# 0.053016f
C7530 XM1/a_n100_n136399# m1_1634_n2388# 3.35e-20
C7531 XM2/a_n158_n274026# XM3/a_n100_n68355# 1.45e-19
C7532 XM2/a_n158_n115866# XM3/a_n158_88178# 4.64e-21
C7533 XM4/w_n358_n132787# XM4/a_n100_23849# -0.004445f
C7534 XM2/a_n158_n92142# XM3/a_n100_115017# 3.46e-20
C7535 XM2/a_n100_n92239# XM3/a_n158_115114# 0.002941f
C7536 XM1/a_n158_n87478# XM3/a_n100_n35203# 1.8e-21
C7537 XM1/a_100_97766# XM2/a_n158_n55238# 0.058832f
C7538 XM3/a_n100_n82859# m1_1634_n2388# 0.072015f
C7539 XM1/a_100_n94658# XM2/a_n100_n247763# 0.005074f
C7540 XM1/a_n158_n40090# XM3/a_n100_10381# 1.94e-20
C7541 XM1/a_n158_n38654# XM3/a_n100_13489# 1.94e-20
C7542 XM1/a_n158_61866# XM3/a_n100_113981# 1.94e-20
C7543 XM1/a_n158_n44398# XM2/a_n158_n197582# 4.64e-21
C7544 XM1/a_100_74790# XM2/a_n158_n78962# 0.116862f
C7545 XM4/w_n358_n132787# XM1/a_n100_n159375# 0.013487f
C7546 XM1/a_n158_n134866# XM2/a_n100_n287303# 3.17e-20
C7547 XM2/a_n100_n268851# XM3/a_n158_n62042# 0.005074f
C7548 XM4/w_n358_n132787# XM2/a_n100_n115963# 0.026527f
C7549 XM2/a_n100_n234583# m1_1634_n2388# 7.61e-19
C7550 XM1/a_n100_n21519# XM2/a_100_n176494# 7.26e-20
C7551 XM3/a_n100_63217# XM4/a_n100_63217# 0.009521f
C7552 XM4/w_n358_n132787# XM4/a_n100_n47635# -0.004445f
C7553 XM1/a_n100_n61727# m1_1634_n2388# 8.14e-20
C7554 XM4/w_n358_n132787# XM2/a_100_n300386# 0.105949f
C7555 XM3/a_n158_n18530# m1_1634_n2388# 6.1e-20
C7556 XM1/a_100_126486# XM4/w_n358_n132787# 0.053546f
C7557 XM1/a_n158_n60194# XM2/a_n100_n216131# 7.26e-20
C7558 XM2/a_n100_n28975# XM4/w_n358_n132787# 0.012279f
C7559 XM4/a_100_58134# m1_1634_n2388# 6.1e-20
C7560 XM1/a_100_179618# XM4/w_n358_n132787# 0.053546f
C7561 XM2/a_100_n15698# XM1/a_100_139410# 4.64e-21
C7562 XM2/a_n158_n15698# XM1/a_n158_139410# 4.64e-21
C7563 XM3/a_n100_100513# m1_1634_n2388# 0.072015f
C7564 XM1/a_100_13042# XM2/a_100_n142226# 4.64e-21
C7565 XM1/a_n158_13042# XM2/a_n100_n139687# 7.26e-20
C7566 XM1/a_n100_n172299# XM3/a_n100_n121191# 3.25e-20
C7567 XM2/a_100_n303022# XM3/a_n158_n97266# 0.077916f
C7568 XM1/a_n100_n109115# XM3/a_n158_n56862# 2.85e-20
C7569 XM1/a_n100_n76087# XM3/a_n100_n24843# 6.89e-19
C7570 XM3/a_n100_n122227# m1_1634_n2388# 0.072015f
C7571 XM1/a_n100_149365# XM2/a_100_n5154# 1.45e-19
C7572 XM1/a_n100_8637# XM2/a_100_n144862# 7.26e-20
C7573 XM1/a_n158_n94658# XM2/a_n100_n247763# 7.26e-20
C7574 XM2/a_n100_n192407# XM3/a_n100_12453# 0.001572f
C7575 XM1/a_100_71918# XM2/a_100_n81598# 4.64e-21
C7576 XM1/a_n158_43198# XM3/a_n100_95333# 1.94e-20
C7577 XM2/a_n158_n213398# XM3/a_n158_n9206# 4.64e-21
C7578 XM1/a_100_47506# XM2/a_n158_n107958# 0.052211f
C7579 XM1/a_n158_n42962# XM3/a_n100_7273# 5.81e-21
C7580 XM1/a_n100_84745# XM4/w_n358_n132787# 0.012279f
C7581 XM2/a_n158_n255574# XM3/a_n100_n50743# 1.45e-19
C7582 XM1/a_100_126486# XM2/a_n100_n26339# 0.005074f
C7583 XM4/a_n100_121233# m1_1634_n2388# 0.072015f
C7584 XM1/a_n158_n166458# XM3/a_n100_n114975# 1.94e-20
C7585 XM4/w_n358_n132787# XM3/a_n100_n27951# 0.008957f
C7586 XM4/a_100_n13350# m1_1634_n2388# 6.1e-20
C7587 XM2/a_n158_n187038# XM3/a_n158_17730# 4.64e-21
C7588 XM2/a_n100_2657# XM4/w_n358_n132787# 0.012279f
C7589 XM1/a_n158_81970# XM2/a_n100_n73787# 7.26e-20
C7590 XM1/a_n100_61769# XM2/a_n158_n92142# 0.010147f
C7591 XM1/a_n158_38890# XM3/a_n100_89117# 4.21e-21
C7592 XM2/a_100_n210762# XM3/a_n158_n4026# 0.045201f
C7593 XM2/a_n100_n195043# XM4/a_100_11514# 1.58e-20
C7594 XM1/a_100_50378# XM2/a_100_n105322# 4.64e-21
C7595 XM2/a_n100_n216131# XM4/a_100_n9206# 2.56e-20
C7596 XM1/a_n158_158078# XM2/a_n158_5390# 4.64e-21
C7597 XM4/w_n358_n132787# XM3/a_n100_62181# 0.009186f
C7598 XM4/w_n358_n132787# XM4/a_n100_n87003# -0.004445f
C7599 XM3/a_n158_n57898# m1_1634_n2388# 6.1e-20
C7600 XM1/a_n100_80437# XM3/a_n100_131593# 6.5e-19
C7601 XM1/a_100_n157842# XM2/a_n100_n313663# 0.005074f
C7602 XM1/a_n158_n126250# XM2/a_n158_n281934# 4.64e-21
C7603 XM1/a_100_n140610# XM3/a_n100_n89075# 2.85e-20
C7604 XM4/w_n358_n132787# XM2/a_n100_n239855# 0.025065f
C7605 XM4/a_100_18766# m1_1634_n2388# 6.1e-20
C7606 XM2/a_n100_18473# XM4/w_n358_n132787# 0.012279f
C7607 XM3/a_n158_125474# m1_1634_n2388# 6.1e-20
C7608 XM1/a_n100_n97627# XM3/a_n158_n45466# 2.85e-20
C7609 XM1/a_n100_n83267# XM2/a_100_n237122# 1.45e-19
C7610 XM1/a_100_n53014# XM2/a_n158_n205490# 0.007423f
C7611 XM1/a_100_148026# XM2/a_n100_n7887# 0.005074f
C7612 XM1/a_n158_83406# XM2/a_n158_n71054# 9.28e-21
C7613 XM2/a_n100_n137051# XM3/a_n100_69433# 4.51e-19
C7614 XM1/a_n158_n139174# XM2/a_n100_n295211# 7.26e-20
C7615 XM1/a_n100_n146451# XM4/w_n358_n132787# 0.013449f
C7616 XM1/a_n100_n86139# m1_1634_n2388# 1.3e-19
C7617 XM1/a_100_118# XM2/a_n100_n152867# 0.005074f
C7618 XM1/a_n158_63302# XM3/a_n100_113981# 1.94e-20
C7619 XM1/a_n158_n147790# XM2/a_n100_n303119# 7.26e-20
C7620 XM2/a_n158_n10426# XM1/a_n100_143621# 0.010147f
C7621 XM2/a_n100_n10523# XM1/a_100_145154# 0.005074f
C7622 XM1/a_n158_152334# XM2/a_n100_n2615# 4.29e-20
C7623 XM1/a_100_109254# XM4/w_n358_n132787# 0.048442f
C7624 XM1/a_100_n25730# XM2/a_n100_n181863# 0.004352f
C7625 XM4/a_n100_81865# m1_1634_n2388# 0.072014f
C7626 XM1/a_n158_n139174# XM3/a_n100_n88039# 2.58e-20
C7627 XM1/a_100_n149226# XM2/a_n158_n303022# 0.116862f
C7628 XM2/a_100_n284570# XM3/a_n158_n79654# 0.077916f
C7629 XM4/w_n358_n132787# XM3/a_n100_n67319# 0.009186f
C7630 XM4/a_100_n52718# m1_1634_n2388# 6.1e-20
C7631 XM1/a_100_n12806# XM3/a_n158_38450# 0.00544f
C7632 XM1/a_100_n8498# XM3/a_n100_42497# 2.85e-20
C7633 XM1/a_100_155206# XM2/a_n100_2657# 0.005074f
C7634 XM2/a_100_n326746# XM3/a_n100_n121191# 0.010147f
C7635 XM1/a_100_163822# XM4/w_n358_n132787# 0.053546f
C7636 XM1/a_n158_110690# XM2/a_n100_n44791# 7.26e-20
C7637 XM4/w_n358_n132787# XM4/a_n100_n126371# -0.004445f
C7638 XM1/a_n100_n157939# XM2/a_n158_n313566# 0.005074f
C7639 XM3/a_n158_n97266# m1_1634_n2388# 6.1e-20
C7640 XM1/a_100_n65938# XM3/a_n100_n15519# 2.85e-20
C7641 XM2/a_n100_n324207# XM3/a_n158_n120058# 0.005074f
C7642 XM2/a_100_n107958# m1_1634_n2388# 0.017213f
C7643 XM2/a_n158_n237122# XM3/a_n100_n33131# 7.26e-20
C7644 XM3/a_n100_45605# m1_1634_n2388# 0.072015f
C7645 XM1/a_100_110690# XM2/a_100_n42058# 4.64e-21
C7646 XM1/a_100_10170# XM3/a_n158_62278# 0.005291f
C7647 XM1/a_100_n41526# XM3/a_n100_9345# 2.85e-20
C7648 XM4/w_n358_n132787# XM2/a_n158_n176494# 0.102824f
C7649 XM2/a_n100_n134415# XM4/a_n100_69433# 2.32e-20
C7650 XM1/a_100_n71682# XM4/w_n358_n132787# 0.050378f
C7651 XM1/a_n158_n28602# XM2/a_n158_n181766# 4.64e-21
C7652 XM1/a_100_n17114# XM2/a_n158_n171222# 0.116862f
C7653 XM1/a_100_150898# XM2/a_100_n2518# 4.64e-21
C7654 XM1/a_n100_n117731# XM3/a_n158_n67222# 2.85e-20
C7655 XM2/a_n158_n321474# XM3/a_n158_n114878# 4.64e-21
C7656 XM4/w_n358_n132787# XM3/a_n158_87142# 0.032295f
C7657 XM1/a_n100_7201# XM3/a_n158_58134# 2.85e-20
C7658 XM2/a_100_n234486# XM3/a_n100_n27951# 0.005074f
C7659 XM4/w_n358_n132787# XM3/a_n158_123402# 0.032295f
C7660 XM1/a_n100_77565# XM2/a_100_n76326# 1.45e-19
C7661 XM4/w_n358_n132787# XM3/a_n158_32234# 0.032295f
C7662 XM4/a_n100_42497# m1_1634_n2388# 0.072015f
C7663 XM4/w_n358_n132787# XM3/a_n100_n106687# 0.009042f
C7664 XM4/a_100_n92086# m1_1634_n2388# 6.1e-20
C7665 XM2/a_n100_n115963# XM3/a_n158_88178# 0.005074f
C7666 XM1/a_n100_153673# XM2/a_n158_118# 0.006883f
C7667 XM2/a_100_n89506# XM3/a_n158_115114# 0.06039f
C7668 XM2/a_n100_n92239# XM3/a_n100_115017# 0.002209f
C7669 XM1/a_n158_n84606# XM2/a_n158_n239758# 4.64e-21
C7670 XM1/a_n100_n57419# XM4/w_n358_n132787# 0.012983f
C7671 XM2/a_100_n208126# XM3/a_n100_n1015# 0.004917f
C7672 XM3/a_n100_31101# XM4/a_n100_31101# 0.009521f
C7673 XM2/a_n100_n84331# XM4/a_100_122366# 2.56e-20
C7674 XM1/a_n100_73257# XM2/a_100_n81598# 7.26e-20
C7675 XM1/a_n158_n30038# XM3/a_n100_21777# 1.94e-20
C7676 XM1/a_n158_n44398# XM2/a_n100_n197679# 7.26e-20
C7677 XM2/a_n100_n271487# XM4/a_100_n67222# 2.56e-20
C7678 XM2/a_100_n266118# XM3/a_n158_n62042# 0.007423f
C7679 XM4/w_n358_n132787# XM2/a_100_n113230# 0.103341f
C7680 XM2/a_100_n308294# XM3/a_n100_n103579# 0.005321f
C7681 XM4/w_n358_n132787# XM3/a_n158_n42358# 0.032295f
C7682 XM4/a_n100_n28987# m1_1634_n2388# 0.072015f
C7683 XM2/a_100_n231850# m1_1634_n2388# 0.025582f
C7684 XM1/a_n100_n21519# XM2/a_n158_n176494# 0.005074f
C7685 avdd XM4/w_n358_n132787# 0.003602f
C7686 XM1/a_100_n127686# XM3/a_n100_n76643# 2.85e-20
C7687 XM1/a_n100_155109# XM2/a_100_118# 7.26e-20
C7688 XM1/a_n100_97669# XM2/a_n158_n55238# 0.005074f
C7689 XM4/w_n358_n132787# XM2/a_n158_n300386# 0.107093f
C7690 XM1/a_n158_94894# XM2/a_n158_n60510# 4.64e-21
C7691 XM1/a_n100_53153# XM4/w_n358_n132787# 0.013458f
C7692 XM3/a_n158_70566# m1_1634_n2388# 6.1e-20
C7693 XM1/a_n158_166694# XM2/a_n100_10565# 4.86e-20
C7694 XM1/a_100_13042# XM2/a_n158_n142226# 0.071295f
C7695 XM1/a_n158_n124814# XM2/a_n158_n279298# 9.28e-21
C7696 XM1/a_n158_74790# XM2/a_n158_n78962# 9.28e-21
C7697 XM2/a_n100_n158139# XM4/a_100_46738# 5.27e-21
C7698 XM1/a_n100_64641# XM4/w_n358_n132787# 0.013401f
C7699 XM3/a_n158_15658# m1_1634_n2388# 6.1e-20
C7700 XM1/a_100_n31474# XM4/w_n358_n132787# 0.054609f
C7701 XM2/a_100_n216034# XM3/a_n100_n10339# 0.010147f
C7702 XM1/a_n158_87714# XM2/a_n100_n65879# 7.26e-20
C7703 XM1/a_n100_8637# XM2/a_n158_n144862# 0.005074f
C7704 XM1/a_n158_n129122# XM2/a_n158_n281934# 4.64e-21
C7705 XM1/a_n158_n57322# XM2/a_n100_n213495# 1.97e-20
C7706 XM1/a_100_71918# XM2/a_n158_n81598# 0.108683f
C7707 XM2/a_n100_n213495# XM3/a_n158_n9206# 0.005074f
C7708 XM1/a_100_172438# XM2/a_n158_18570# 0.116862f
C7709 XM4/w_n358_n132787# XM4/a_n100_97405# -0.004445f
C7710 XM1/a_100_47506# XM2/a_n100_n108055# 0.005074f
C7711 XM1/a_n100_n64599# XM2/a_100_n218670# 1.45e-19
C7712 XM4/w_n358_n132787# XM1/a_n100_143621# 0.012279f
C7713 XM3/a_n100_n9303# m1_1634_n2388# 0.072015f
C7714 XM1/a_100_122178# XM4/w_n358_n132787# 0.048442f
C7715 XM4/w_n358_n132787# XM3/a_n158_n81726# 0.032295f
C7716 XM4/a_n100_n68355# m1_1634_n2388# 0.072015f
C7717 XM2/a_n100_n187135# XM3/a_n158_17730# 6.5e-19
C7718 XM2/a_n158_n210762# XM3/a_n158_n4026# 4.64e-21
C7719 XM4/w_n358_n132787# XM3/a_n100_1057# 0.009182f
C7720 XM1/a_100_50378# XM2/a_n158_n105322# 0.029233f
C7721 XM1/a_n100_n116295# XM3/a_n158_n64114# 2.85e-20
C7722 XM1/a_n100_n86139# XM2/a_100_n239758# 1.45e-19
C7723 XM1/a_n100_n51675# XM4/w_n358_n132787# 0.013627f
C7724 XM2/a_n100_n171319# m1_1634_n2388# 7.61e-19
C7725 XM1/a_n158_n126250# XM2/a_n100_n282031# 7.26e-20
C7726 XM1/a_100_84842# XM2/a_n158_n68418# 0.083758f
C7727 XM1/a_100_n157842# XM2/a_100_n310930# 4.64e-21
C7728 XM4/w_n358_n132787# XM2/a_100_n237122# 0.10657f
C7729 XM1/a_n158_n159278# XM3/a_n100_n108759# 1.94e-20
C7730 XM4/w_n358_n132787# XM1/a_n100_178085# 0.012279f
C7731 XM3/a_n100_125377# m1_1634_n2388# 0.072015f
C7732 XM1/a_n158_n176510# XM2/a_n158_n329382# 4.64e-21
C7733 XM2/a_100_n289842# XM3/a_n100_n85967# 0.004513f
C7734 XM1/a_100_n113326# XM4/w_n358_n132787# 0.054609f
C7735 XM1/a_n100_n83267# XM2/a_n158_n237122# 0.010147f
C7736 XM1/a_100_n53014# XM2/a_n100_n205587# 0.005074f
C7737 XM4/a_100_131690# m1_1634_n2388# 3.05e-20
C7738 XM1/a_100_n121942# XM3/a_n100_n71463# 2.85e-20
C7739 XM1/a_n158_n34346# XM3/a_n100_17633# 1e-20
C7740 XM1/a_n158_n1318# XM2/a_n158_n155406# 9.28e-21
C7741 XM2/a_n100_n15795# XM1/a_n100_136441# 0.002019f
C7742 XM4/w_n358_n132787# XM4/a_n100_58037# -0.004445f
C7743 XM3/a_n100_n48671# m1_1634_n2388# 0.072015f
C7744 XM1/a_100_n4190# XM2/a_n158_n158042# 0.116862f
C7745 XM1/a_n100_n162247# XM2/a_100_n316202# 1.45e-19
C7746 XM1/a_n100_n152195# XM3/a_n158_n101410# 0.001493f
C7747 XM1/a_100_n54450# XM3/a_n100_n3087# 5.71e-20
C7748 XM4/a_100_118# m1_1634_n2388# 6.1e-20
C7749 XM1/a_n100_n43059# XM3/a_n100_7273# 8.85e-19
C7750 XM1/a_100_n25730# XM2/a_100_n179130# 4.64e-21
C7751 XM1/a_n158_113562# XM2/a_n100_n42155# 7.26e-20
C7752 XM1/a_100_n165022# XM2/a_n158_n318838# 0.116862f
C7753 XM1/a_n100_n30135# XM3/a_n158_20838# 2.85e-20
C7754 XM2/a_n100_n139687# XM4/a_100_64350# 9.75e-21
C7755 XM4/a_100_n130418# XM2/a_n100_n337387# 2.56e-20
C7756 XM4/w_n358_n132787# XM3/a_n158_n121094# 0.032295f
C7757 XM4/a_n100_n107723# m1_1634_n2388# 0.072015f
C7758 XM3/a_n100_n6195# XM4/a_n100_n6195# 0.009521f
C7759 XM4/w_n358_n132787# XM1/a_100_135102# 0.052325f
C7760 XM2/a_n158_n326746# XM3/a_n100_n121191# 1.45e-19
C7761 XM1/a_n158_n149226# XM3/a_n100_n98399# 1.94e-20
C7762 XM1/a_n100_n145015# m1_1634_n2388# 1.3e-19
C7763 XM1/a_100_n91786# XM3/a_n158_n40286# 0.001549f
C7764 XM1/a_100_n61630# XM2/a_n158_n216034# 0.116862f
C7765 XM1/a_n158_57558# XM3/a_n100_108801# 3.71e-20
C7766 XM1/a_n158_n142046# XM2/a_n158_n295114# 4.64e-21
C7767 XM4/w_n358_n132787# XM3/a_n100_80829# 0.008405f
C7768 XM1/a_n158_n100402# XM2/a_n158_n252938# 4.64e-21
C7769 XM4/w_n358_n132787# XM4/a_n100_n13447# -0.004445f
C7770 XM1/a_100_8734# XM3/a_n158_59170# 1.53e-19
C7771 XM4/w_n358_n132787# XM2/a_n100_n176591# 0.026356f
C7772 XM2/a_n100_n295211# m1_1634_n2388# 7.61e-19
C7773 XM1/a_n158_n28602# XM2/a_n100_n181863# 7.26e-20
C7774 XM4/w_n358_n132787# XM3/a_n100_25921# 0.008905f
C7775 XM1/a_100_76226# XM3/a_n100_128485# 2.85e-20
C7776 XM4/a_100_92322# m1_1634_n2388# 6.1e-20
C7777 XM2/a_n100_n321571# XM3/a_n158_n114878# 0.005074f
C7778 XM2/a_n158_n23606# XM1/a_100_132230# 0.015991f
C7779 XM2/a_100_n23606# XM1/a_n100_130697# 1.45e-19
C7780 XM1/a_n100_104849# XM2/a_n158_n49966# 0.005074f
C7781 XM3/a_n100_83937# XM4/a_n100_83937# 0.009521f
C7782 XM2/a_100_n121138# XM3/a_n100_83937# 0.010147f
C7783 XM2/a_n158_n234486# XM3/a_n100_n27951# 7.26e-20
C7784 XM4/w_n358_n132787# XM4/a_n100_18669# -0.004445f
C7785 XM4/w_n358_n132787# XM3/a_n100_123305# 0.009186f
C7786 XM1/a_n100_77565# XM2/a_n158_n76326# 0.010147f
C7787 XM3/a_n100_n88039# m1_1634_n2388# 0.072014f
C7788 XM2/a_100_n163314# XM3/a_n100_41461# 0.00864f
C7789 XM1/a_n100_54589# XM4/w_n358_n132787# 0.013511f
C7790 XM1/a_n158_n84606# XM2/a_n100_n239855# 7.26e-20
C7791 XM3/a_n100_n25879# XM4/a_n100_n25879# 0.009521f
C7792 XM1/a_n100_n17211# XM3/a_n158_35342# 1.29e-20
C7793 XM2/a_n158_n89506# XM3/a_n158_115114# 4.64e-21
C7794 XM2/a_100_n89506# XM3/a_n100_115017# 0.005074f
C7795 XM2/a_n158_n208126# XM3/a_n100_n1015# 6.66e-20
C7796 XM2/a_n158_n57874# XM4/w_n358_n132787# 0.107093f
C7797 XM1/a_100_n116198# XM3/a_n100_n65247# 2.85e-20
C7798 XM1/a_n158_n67374# XM3/a_n100_n16555# 1.94e-20
C7799 XM1/a_n100_73257# XM2/a_n158_n81598# 0.005074f
C7800 XM1/a_100_n131994# m1_1634_n2388# 0.002002f
C7801 XM4/w_n358_n132787# XM4/a_n100_n52815# -0.004445f
C7802 XM2/a_n158_n266118# XM3/a_n158_n62042# 4.64e-21
C7803 XM3/a_n158_n23710# m1_1634_n2388# 6.1e-20
C7804 XM1/a_n100_127825# XM4/w_n358_n132787# 0.012279f
C7805 XM1/a_100_21658# XM4/w_n358_n132787# 0.054609f
C7806 XM1/a_n100_n130655# XM3/a_n158_n79654# 2.85e-20
C7807 XM4/a_100_52954# m1_1634_n2388# 6.1e-20
C7808 XM1/a_100_163822# XM2/a_100_8026# 4.64e-21
C7809 XM1/a_100_70482# XM2/a_n158_n84234# 0.116862f
C7810 XM3/a_n100_64253# m1_1634_n2388# 0.072015f
C7811 XM1/a_n158_97766# XM2/a_n158_n57874# 4.64e-21
C7812 XM4/w_n358_n132787# XM2/a_n158_n113230# 0.101988f
C7813 XM2/a_n158_n308294# XM3/a_n100_n103579# 8.15e-20
C7814 XM2/a_n158_n231850# m1_1634_n2388# 2.36e-21
C7815 XM3/a_n100_9345# m1_1634_n2388# 0.072015f
C7816 XM1/a_n158_n27166# XM3/a_n100_24885# 1.94e-20
C7817 XM2/a_100_n107958# XM3/a_n100_98441# 0.005074f
C7818 XM3/a_n100_n127407# m1_1634_n2388# 0.072015f
C7819 XM4/w_n358_n132787# XM2/a_n100_n300483# 0.024572f
C7820 XM2/a_100_n263482# XM3/a_n158_n56862# 0.056495f
C7821 XM1/a_100_94894# XM2/a_n100_n57971# 0.005074f
C7822 XM2/a_n100_n268851# XM4/a_100_n62042# 2.56e-20
C7823 XM1/a_n158_n60194# XM2/a_n158_n213398# 4.64e-21
C7824 XM3/a_n158_101646# m1_1634_n2388# 6.1e-20
C7825 XM1/a_n100_n34443# XM3/a_n158_17730# 2.85e-20
C7826 XM1/a_n158_n19986# XM2/a_n158_n173858# 9.28e-21
C7827 XM1/a_100_13042# XM2/a_n100_n142323# 0.005074f
C7828 XM1/a_100_n166458# m1_1634_n2388# 6.08e-19
C7829 XM1/a_100_n133430# XM3/a_n100_n82859# 2.85e-20
C7830 XM4/a_n100_5201# m1_1634_n2388# 0.072015f
C7831 XM4/w_n358_n132787# XM3/a_n158_50882# 0.032295f
C7832 XM2/a_100_n150134# XM3/a_n100_55965# 0.010147f
C7833 XM1/a_n100_n170863# XM3/a_n158_n119022# 2.85e-20
C7834 XM3/a_n100_n45563# XM4/a_n100_n45563# 0.009521f
C7835 XM1/a_100_173874# XM4/w_n358_n132787# 0.053546f
C7836 XM1/a_n100_70385# XM2/a_100_n84234# 1.38e-19
C7837 XM4/a_n100_116053# m1_1634_n2388# 0.072015f
C7838 XM2/a_n158_n216034# XM3/a_n100_n10339# 1.45e-19
C7839 XM1/a_n100_8637# XM2/a_n100_n144959# 0.006262f
C7840 XM1/a_n158_n129122# XM2/a_n100_n282031# 7.26e-20
C7841 XM4/w_n358_n132787# XM3/a_n100_n33131# 0.008966f
C7842 XM4/a_100_n18530# m1_1634_n2388# 6.1e-20
C7843 XM2/a_100_n192310# XM3/a_n100_13489# 0.010147f
C7844 XM1/a_100_71918# XM2/a_n100_n81695# 0.004619f
C7845 XM1/a_100_47506# XM2/a_100_n105322# 4.64e-21
C7846 XM4/w_n358_n132787# XM4/a_n100_n92183# -0.004445f
C7847 XM1/a_100_n107582# XM2/a_100_n263482# 4.64e-21
C7848 XM1/a_n100_n64599# XM2/a_n158_n218670# 0.010147f
C7849 XM3/a_n158_n63078# m1_1634_n2388# 6.1e-20
C7850 XM1/a_100_n48706# XM2/a_n158_n202854# 0.116862f
C7851 XM4/a_100_13586# m1_1634_n2388# 6.1e-20
C7852 XM2/a_n100_n210859# XM3/a_n158_n4026# 0.005074f
C7853 XM1/a_100_50378# XM2/a_n100_n105419# 0.005074f
C7854 XM2/a_100_n337290# XM3/a_n158_n132490# 0.077904f
C7855 XM1/a_n158_n131994# XM3/a_n100_n80787# 2.89e-20
C7856 XM1/a_n100_n86139# XM2/a_n158_n239758# 0.010147f
C7857 XM2/a_100_n168586# m1_1634_n2388# 0.023368f
C7858 XM1/a_n100_n93319# XM3/a_n158_n41322# 2.85e-20
C7859 XM1/a_100_n80298# XM3/a_n100_n30023# 2.11e-20
C7860 XM1/a_100_n40090# XM3/a_n100_10381# 2.85e-20
C7861 XM1/a_100_n157842# XM2/a_n158_n310930# 0.067011f
C7862 XM4/w_n358_n132787# XM2/a_n158_n237122# 0.107093f
C7863 XM1/a_n100_n119167# m1_1634_n2388# 7.61e-20
C7864 XM3/a_n158_89214# m1_1634_n2388# 6.1e-20
C7865 XM1/a_n158_n176510# XM2/a_n100_n329479# 7.26e-20
C7866 XM3/a_n100_n65247# XM4/a_n100_n65247# 0.009521f
C7867 XM1/a_100_40326# XM2/a_100_n113230# 4.64e-21
C7868 XM2/a_n158_n289842# XM3/a_n100_n85967# 5.16e-20
C7869 XM1/a_n158_120742# XM2/a_n100_n34247# 6.88e-20
C7870 XM4/a_n100_76685# m1_1634_n2388# 0.072015f
C7871 XM1/a_n158_162386# XM2/a_n158_8026# 9.28e-21
C7872 XM1/a_n158_n139174# XM2/a_n158_n292478# 4.64e-21
C7873 XM4/w_n358_n132787# XM3/a_n100_n72499# 0.009147f
C7874 XM4/a_100_n57898# m1_1634_n2388# 6.1e-20
C7875 XM3/a_n158_34306# m1_1634_n2388# 6.1e-20
C7876 XM1/a_n158_34582# XM3/a_n100_86009# 2.58e-20
C7877 XM2/a_100_n245030# XM3/a_n158_n39250# 0.077916f
C7878 XM1/a_n100_n5723# XM2/a_100_n160678# 7.26e-20
C7879 XM1/a_n158_n147790# XM2/a_n158_n300386# 4.64e-21
C7880 XM2/a_100_n179130# XM3/a_n100_27993# 0.004675f
C7881 XM1/a_n158_20222# XM3/a_n100_70469# 8.22e-21
C7882 XM3/a_n158_n102446# m1_1634_n2388# 6.1e-20
C7883 XM2/a_100_n287206# XM3/a_n100_n80787# 0.005074f
C7884 XM1/a_n100_n162247# XM2/a_n158_n316202# 0.010147f
C7885 XM1/a_100_n25730# XM2/a_n158_n179130# 0.097389f
C7886 XM1/a_n158_30274# XM3/a_n100_81865# 1.94e-20
C7887 XM1/a_100_n25730# XM3/a_n100_24885# 2.85e-20
C7888 XM1/a_n100_60333# XM3/a_n100_111909# 7.98e-19
C7889 XM1/a_100_n88914# XM4/w_n358_n132787# 0.051632f
C7890 XM1/a_100_n22858# XM4/w_n358_n132787# 0.048442f
C7891 XM3/a_n100_51821# XM4/a_n100_51821# 0.009521f
C7892 XM1/a_n100_76129# XM3/a_n158_128582# 2.85e-20
C7893 XM1/a_n100_n183787# sw_b 8.1e-20
C7894 XM1/a_n100_n157939# XM2/a_100_n310930# 7.26e-20
C7895 XM1/a_100_n81734# XM3/a_n158_n29926# 0.00544f
C7896 XM4/w_n358_n132787# XM3/a_n158_n8170# 0.032295f
C7897 XM1/a_n158_n142046# XM2/a_n100_n295211# 7.26e-20
C7898 XM1/a_100_n45834# XM3/a_n100_6237# 2.85e-20
C7899 XM2/a_n100_n108055# m1_1634_n2388# 7.65e-19
C7900 XM1/a_n158_n100402# XM2/a_n100_n253035# 7.26e-20
C7901 XM1/a_100_173874# XM2/a_n100_21109# 0.005074f
C7902 XM2/a_n100_n137051# XM4/a_100_69530# 2.21e-20
C7903 XM1/a_n100_n106243# m1_1634_n2388# 7.61e-20
C7904 XM3/a_n100_n84931# XM4/a_n100_n84931# 0.009521f
C7905 XM4/w_n358_n132787# XM2/a_100_n173858# 0.10657f
C7906 XM3/a_n100_128485# XM4/a_n100_128485# 0.009521f
C7907 XM2/a_100_n292478# m1_1634_n2388# 0.017213f
C7908 XM4/a_n100_37317# m1_1634_n2388# 0.072015f
C7909 XM1/a_n100_1457# XM3/a_n158_53990# 1.87e-20
C7910 XM1/a_100_7298# XM3/a_n100_58037# 2.85e-20
C7911 XM2/a_n100_n324207# XM4/a_100_n120058# 2.56e-20
C7912 XM4/w_n358_n132787# XM3/a_n100_n111867# 0.009122f
C7913 XM4/a_100_n97266# m1_1634_n2388# 6.1e-20
C7914 XM1/a_100_158078# XM2/a_n100_2657# 0.005074f
C7915 XM2/a_n158_n121138# XM3/a_n100_83937# 1.45e-19
C7916 XM1/a_n100_n122039# XM4/w_n358_n132787# 0.013218f
C7917 XM1/a_n100_n54547# XM3/a_n100_n2051# 0.001249f
C7918 XM1/a_100_50378# XM3/a_n100_102585# 2.85e-20
C7919 XM1/a_n100_n179479# XM3/a_n158_n127310# 2.85e-20
C7920 XM1/a_100_n129122# XM3/a_n100_n78715# 2.85e-20
C7921 XM1/a_100_n88914# XM3/a_n100_n38311# 2.85e-20
C7922 XM2/a_n100_n73787# XM4/w_n358_n132787# 0.019008f
C7923 XM2/a_n158_5390# XM4/w_n358_n132787# 0.107093f
C7924 XM2/a_n158_n163314# XM3/a_n100_41461# 1.3e-19
C7925 XM1/a_100_118# XM3/a_n100_51821# 3.38e-19
C7926 XM4/w_n358_n132787# XM4/a_n100_131593# -3.9e-19
C7927 XM2/a_100_n115866# XM3/a_n158_89214# 0.077916f
C7928 XM1/a_100_100638# XM4/w_n358_n132787# 0.053546f
C7929 XM2/a_n100_n89603# XM3/a_n158_115114# 0.005074f
C7930 XM2/a_n158_n89506# XM3/a_n100_115017# 7.26e-20
C7931 XM2/a_n100_n208223# XM3/a_n100_n1015# 2.49e-19
C7932 XM1/a_n158_n179382# XM3/a_n100_n127407# 9.42e-21
C7933 XM1/a_n158_n156406# XM3/a_n100_n104615# 1.94e-20
C7934 XM2/a_100_n226578# XM3/a_n158_n21638# 0.077916f
C7935 XM4/w_n358_n132787# XM3/a_n158_n47538# 0.032295f
C7936 XM4/a_n100_n34167# m1_1634_n2388# 0.072015f
C7937 XM2/a_100_n158042# XM3/a_n158_46738# 0.075968f
C7938 XM2/a_100_n268754# XM3/a_n100_n63175# 0.010147f
C7939 XM1/a_n158_n117634# XM3/a_n100_n67319# 1.94e-20
C7940 XM1/a_n100_n83267# XM4/w_n358_n132787# 0.013411f
C7941 XM4/w_n358_n132787# XM3/a_n100_99477# 0.009163f
C7942 XM3/a_n100_n104615# XM4/a_n100_n104615# 0.009521f
C7943 XM2/a_n100_n266215# XM3/a_n158_n62042# 0.005074f
C7944 XM1/a_n158_93458# XM2/a_n158_n60510# 9.28e-21
C7945 XM1/a_n100_21561# XM2/a_100_n134318# 7.26e-20
C7946 XM1/a_n100_n155067# m1_1634_n2388# 8.07e-20
C7947 XM1/a_n100_126389# XM2/a_100_n28878# 7.26e-20
C7948 XM1/a_n100_n21519# XM2/a_100_n173858# 7.26e-20
C7949 XM4/w_n358_n132787# XM2/a_n100_n113327# 0.02579f
C7950 XM2/a_n100_n308391# XM3/a_n100_n103579# 0.005614f
C7951 XM2/a_n100_n231947# m1_1634_n2388# 7.8e-19
C7952 XM4/w_n358_n132787# XM3/a_n100_44569# 0.009026f
C7953 XM2/a_n100_n76423# XM4/a_n100_127449# 1.02e-20
C7954 XM1/a_100_n58758# XM4/w_n358_n132787# 0.048442f
C7955 XM2/a_n158_n107958# XM3/a_n100_98441# 7.26e-20
C7956 XM4/w_n358_n132787# XM2/a_100_n297750# 0.103341f
C7957 XM1/a_n100_n114859# XM3/a_n158_n64114# 2.85e-20
C7958 XM2/a_n158_n263482# XM3/a_n158_n56862# 4.64e-21
C7959 XM1/a_n158_n60194# XM2/a_n100_n213495# 7.26e-20
C7960 XM3/a_n100_101549# m1_1634_n2388# 0.072015f
C7961 XM1/a_100_n150662# XM3/a_n100_n99435# 3.43e-19
C7962 XM4/w_n358_n132787# XM4/a_n100_92225# -0.004445f
C7963 XM1/a_100_13042# XM2/a_100_n139590# 4.64e-21
C7964 XM2/a_n158_n150134# XM3/a_n100_55965# 1.45e-19
C7965 XM3/a_n100_n14483# m1_1634_n2388# 0.072015f
C7966 XM1/a_100_n53014# XM3/a_n100_n1015# 5.79e-20
C7967 XM1/a_n100_70385# XM2/a_n158_n84234# 0.009693f
C7968 XM3/a_n100_111909# XM4/a_n100_111909# 0.009521f
C7969 XM4/w_n358_n132787# XM3/a_n158_n86906# 0.032295f
C7970 XM4/a_n100_n73535# m1_1634_n2388# 0.072014f
C7971 XM1/a_n158_n57322# XM2/a_n158_n210762# 4.64e-21
C7972 XM2/a_n158_n192310# XM3/a_n100_13489# 1.45e-19
C7973 XM2/a_n158_n10426# XM4/w_n358_n132787# 0.107093f
C7974 XM1/a_100_47506# XM2/a_n158_n105322# 0.041696f
C7975 XM1/a_100_n130558# XM2/a_n158_n284570# 0.116862f
C7976 XM1/a_100_n107582# XM2/a_n158_n263482# 0.00976f
C7977 XM1/a_100_n103274# XM3/a_n158_n51682# 0.0031f
C7978 XM1/a_100_67610# XM2/a_n158_n86870# 0.116862f
C7979 XM2/a_100_n144862# XM3/a_n158_61242# 0.077916f
C7980 XM3/a_n100_n124299# XM4/a_n100_n124299# 0.009521f
C7981 XM1/a_100_8734# XM2/a_100_n144862# 4.64e-21
C7982 XM1/a_n158_126486# XM2/a_n158_n26242# 4.64e-21
C7983 XM3/a_n100_82901# m1_1634_n2388# 0.072015f
C7984 XM2/a_100_n187038# XM3/a_n158_18766# 0.077916f
C7985 XM1/a_n100_122081# XM2/a_n158_n31514# 0.010051f
C7986 XM2/a_100_n208126# XM3/a_n158_n4026# 0.00976f
C7987 XM1/a_100_50378# XM2/a_100_n102686# 4.64e-21
C7988 XM1/a_n100_7201# XM2/a_100_n147498# 7.56e-20
C7989 XM1/a_100_n64502# XM4/w_n358_n132787# 0.048442f
C7990 XM2/a_n100_n213495# XM4/a_100_n9206# 2.56e-20
C7991 XM4/a_100_126510# m1_1634_n2388# 6.1e-20
C7992 XM1/a_n158_n126250# XM2/a_n158_n279298# 4.64e-21
C7993 XM2/a_100_n250302# XM3/a_n100_n45563# 0.005805f
C7994 XM3/a_n100_n3087# m1_1634_n2388# 0.072015f
C7995 XM1/a_100_n157842# XM2/a_n100_n311027# 0.005074f
C7996 XM3/a_n100_27993# m1_1634_n2388# 0.072015f
C7997 XM1/a_n158_37454# XM3/a_n100_89117# 1.94e-20
C7998 XM4/w_n358_n132787# XM2/a_n100_n237219# 0.025738f
C7999 XM4/w_n358_n132787# XM4/a_n100_52857# -0.004445f
C8000 XM1/a_100_160950# XM2/a_n100_7929# 0.005074f
C8001 XM3/a_n158_126510# m1_1634_n2388# 6.1e-20
C8002 XM2/a_n100_n289939# XM3/a_n100_n85967# 8.7e-19
C8003 XM1/a_100_n130558# XM3/a_n100_n79751# 2.85e-20
C8004 XM3/a_n100_n53851# m1_1634_n2388# 0.072015f
C8005 XM1/a_100_40326# XM2/a_n158_n113230# 0.112578f
C8006 XM1/a_n100_n127783# XM2/a_100_n281934# 1.45e-19
C8007 XM4/w_n358_n132787# XM3/a_n158_69530# 0.033922f
C8008 XM2/a_n100_n134415# XM3/a_n100_69433# 0.002666f
C8009 XM4/w_n358_n132787# XM3/a_n158_n126274# 0.032295f
C8010 XM1/a_100_n167894# XM2/a_100_n321474# 4.64e-21
C8011 XM4/a_n100_n112903# m1_1634_n2388# 0.072015f
C8012 XM1/a_n158_n139174# XM2/a_n100_n292575# 7.26e-20
C8013 XM3/a_n100_19705# XM4/a_n100_19705# 0.009521f
C8014 XM1/a_n100_n96191# XM2/a_100_n250302# 1.45e-19
C8015 XM1/a_n100_n5723# XM2/a_n158_n160678# 0.005074f
C8016 XM1/a_n158_63302# XM3/a_n100_115017# 8.22e-21
C8017 XM1/a_n158_n147790# XM2/a_n100_n300483# 7.26e-20
C8018 XM4/w_n358_n132787# XM3/a_n158_14622# 0.038462f
C8019 XM2/a_n158_n179130# XM3/a_n100_27993# 5.76e-20
C8020 XM1/a_100_30274# XM3/a_n100_80829# 2.85e-20
C8021 XM2/a_n158_n287206# XM3/a_n100_n80787# 7.26e-20
C8022 XM1/a_100_n25730# XM2/a_n100_n179227# 0.005074f
C8023 XM1/a_n100_66077# m1_1634_n2388# 1.3e-19
C8024 XM1/a_n100_22997# XM3/a_n158_74710# 5.5e-21
C8025 XM4/w_n358_n132787# XM4/a_n100_n18627# -0.004445f
C8026 XM1/a_100_110690# XM4/w_n358_n132787# 0.053546f
C8027 XM1/a_n158_107818# XM2/a_n158_n44694# 4.64e-21
C8028 XM2/a_100_n173858# XM3/a_n158_33270# 0.007033f
C8029 XM4/a_100_87142# m1_1634_n2388# 6.1e-20
C8030 XM1/a_n100_n157939# XM2/a_n158_n310930# 0.005074f
C8031 XM2/a_100_n105322# m1_1634_n2388# 0.020206f
C8032 XM1/a_100_n84606# XM2/a_100_n239758# 4.64e-21
C8033 XM4/w_n358_n132787# XM4/a_n100_13489# -0.004445f
C8034 XM1/a_n158_n119070# XM3/a_n100_n67319# 1.94e-20
C8035 XM1/a_n158_n84606# XM3/a_n100_n33131# 2.5e-20
C8036 XM1/a_n100_n70343# XM3/a_n158_n19566# 3.22e-20
C8037 XM3/a_n100_n3087# XM4/a_n100_n3087# 0.009521f
C8038 XM1/a_n100_n166555# m1_1634_n2388# 1.34e-19
C8039 XM3/a_n100_n93219# m1_1634_n2388# 0.072015f
C8040 XM4/w_n358_n132787# XM2/a_n158_n173858# 0.107093f
C8041 XM4/w_n358_n132787# XM1/a_100_n183690# 0.048442f
C8042 XM1/a_n100_21# XM3/a_n158_50882# 2.85e-20
C8043 XM1/a_100_n163586# XM2/a_100_n318838# 4.64e-21
C8044 XM2/a_100_n231850# XM3/a_n100_n27951# 0.004998f
C8045 XM4/w_n358_n132787# XM3/a_n158_124438# 0.032295f
C8046 XM1/a_100_n177946# XM4/w_n358_n132787# 0.048442f
C8047 XM1/a_n158_n1318# XM3/a_n100_50785# 1.94e-20
C8048 XM3/a_n158_52954# m1_1634_n2388# 6.1e-20
C8049 XM4/w_n358_n132787# XM3/a_n158_2190# 0.032295f
C8050 XM1/a_100_n50142# XM3/a_n100_1057# 5.7e-20
C8051 XM2/a_n100_n163411# XM3/a_n100_41461# 0.001011f
C8052 XM2/a_n100_n321571# XM4/a_100_n114878# 2.56e-20
C8053 XM2/a_100_n316202# XM3/a_n158_n109698# 0.06779f
C8054 XM4/w_n358_n132787# XM4/a_n100_n57995# -0.004445f
C8055 XM1/a_n158_n84606# XM2/a_n158_n237122# 4.64e-21
C8056 XM3/a_n158_n28890# m1_1634_n2388# 6.1e-20
C8057 XM2/a_100_n89506# XM3/a_n158_116150# 0.077916f
C8058 XM2/a_100_n205490# XM3/a_n100_n1015# 0.005074f
C8059 XM4/a_100_47774# m1_1634_n2388# 6.1e-20
C8060 XM2/a_n100_n81695# XM4/a_100_122366# 1.61e-20
C8061 XM1/a_n158_n157842# XM3/a_n100_n105651# 1.94e-20
C8062 XM1/a_n158_n40090# XM3/a_n100_11417# 1.94e-20
C8063 XM2/a_n158_n158042# XM3/a_n158_46738# 4.64e-21
C8064 XM1/a_n100_73257# XM2/a_100_n78962# 1.37e-20
C8065 XM2/a_n158_n268754# XM3/a_n100_n63175# 1.45e-19
C8066 XM1/a_n100_38793# m1_1634_n2388# 4.34e-20
C8067 XM3/a_n100_n132587# m1_1634_n2388# 0.036019f
C8068 XM1/a_n100_21561# XM2/a_n158_n134318# 0.005074f
C8069 XM1/a_n100_n21519# XM2/a_n158_n173858# 0.005074f
C8070 XM4/w_n358_n132787# XM2/a_100_n110594# 0.106086f
C8071 XM1/a_n100_n165119# XM2/a_100_n318838# 1.45e-19
C8072 XM2/a_100_n229214# m1_1634_n2388# 0.017213f
C8073 XM1/a_100_17350# XM2/a_n158_n136954# 0.116862f
C8074 XM1/a_100_n114762# XM4/w_n358_n132787# 0.048442f
C8075 XM4/a_n100_110873# m1_1634_n2388# 0.072015f
C8076 XM2/a_n100_n108055# XM3/a_n100_98441# 3.11e-20
C8077 XM4/w_n358_n132787# XM2/a_n158_n297750# 0.107093f
C8078 XM2/a_n100_n263579# XM3/a_n158_n56862# 0.005074f
C8079 XM4/w_n358_n132787# XM3/a_n100_n38311# 0.009186f
C8080 XM4/a_100_n23710# m1_1634_n2388# 6.1e-20
C8081 XM2/a_n100_n26339# XM4/w_n358_n132787# 0.012279f
C8082 XM2/a_n100_n305755# XM3/a_n100_n98399# 0.002886f
C8083 XM1/a_n100_n33007# XM2/a_100_n187038# 1.45e-19
C8084 XM2/a_n158_n13062# XM1/a_n158_139410# 4.64e-21
C8085 XM2/a_100_n13062# XM1/a_100_139410# 4.64e-21
C8086 XM1/a_100_13042# XM2/a_n158_n139590# 0.022612f
C8087 XM4/w_n358_n132787# XM4/a_n100_n97363# -0.004445f
C8088 XM1/a_n100_n145015# XM2/a_100_n300386# 7.26e-20
C8089 XM1/a_n158_160950# XM2/a_n100_7929# 7.26e-20
C8090 XM3/a_n158_n68258# m1_1634_n2388# 6.1e-20
C8091 XM1/a_n100_70385# XM2/a_n100_n84331# 4.51e-19
C8092 XM1/a_n100_43101# XM3/a_n158_94394# 1.97e-21
C8093 XM1/a_n158_n57322# XM2/a_n100_n210859# 7.26e-20
C8094 XM1/a_n100_87617# XM2/a_n158_n65782# 0.005074f
C8095 XM1/a_100_155206# XM4/w_n358_n132787# 0.053546f
C8096 XM1/a_100_47506# XM2/a_n100_n105419# 0.005074f
C8097 XM1/a_100_n107582# XM2/a_n100_n263579# 0.005074f
C8098 XM1/a_n100_n21519# XM4/w_n358_n132787# 0.013373f
C8099 XM2/a_100_n297750# XM3/a_n158_n92086# 0.077916f
C8100 XM1/a_100_8734# XM2/a_n158_n144862# 0.116473f
C8101 XM1/a_n158_81970# XM2/a_n100_n71151# 7.26e-20
C8102 XM1/a_n158_n111890# XM2/a_n158_n266118# 9.28e-21
C8103 XM1/a_n100_150801# XM2/a_100_n5154# 3.76e-20
C8104 XM1/a_n158_38890# XM3/a_n100_90153# 3.89e-20
C8105 XM2/a_n158_n208126# XM3/a_n158_n4026# 4.64e-21
C8106 XM1/a_n100_4329# XM4/w_n358_n132787# 0.013436f
C8107 XM1/a_100_50378# XM2/a_n158_n102686# 0.064674f
C8108 XM1/a_n100_7201# XM2/a_n158_n147498# 0.005159f
C8109 XM2/a_n100_n337387# XM3/a_n158_n132490# 4.68e-21
C8110 XM1/a_100_n38654# XM4/w_n358_n132787# 0.048442f
C8111 XM2/a_n100_n168683# m1_1634_n2388# 0.002282f
C8112 XM3/a_n100_72541# XM4/a_n100_72541# 0.009521f
C8113 XM4/a_n100_71505# m1_1634_n2388# 0.072015f
C8114 XM4/w_n358_n132787# XM3/a_n100_63217# 0.009026f
C8115 XM1/a_n158_n126250# XM2/a_n100_n279395# 7.26e-20
C8116 XM2/a_n158_n250302# XM3/a_n100_n45563# 9.95e-20
C8117 XM4/w_n358_n132787# XM3/a_n100_n77679# 0.009068f
C8118 XM4/a_100_n63078# m1_1634_n2388# 6.1e-20
C8119 XM1/a_n100_n89011# XM3/a_n158_n38214# 6e-19
C8120 XM4/w_n358_n132787# XM2/a_100_n234486# 0.103341f
C8121 XM1/a_n100_38793# XM2/a_100_n115866# 1.09e-19
C8122 XM1/a_100_4426# XM2/a_n158_n150134# 0.116862f
C8123 XM1/a_n158_n169330# XM2/a_n158_n324110# 9.28e-21
C8124 XM1/a_n100_n60291# XM3/a_n158_n8170# 2.85e-20
C8125 XM2/a_n100_21109# XM4/w_n358_n132787# 0.012279f
C8126 XM3/a_n100_126413# m1_1634_n2388# 0.072015f
C8127 XM3/a_n158_n107626# m1_1634_n2388# 6.1e-20
C8128 XM1/a_100_40326# XM2/a_n100_n113327# 0.001105f
C8129 XM1/a_n100_n127783# XM2/a_n158_n281934# 0.010147f
C8130 XM2/a_n100_n210859# XM4/a_100_n4026# 2.56e-20
C8131 XM1/a_100_148026# XM2/a_n100_n5251# 0.005074f
C8132 XM1/a_n158_n75990# XM2/a_n158_n231850# 4.64e-21
C8133 XM1/a_n100_n68907# m1_1634_n2388# 9.25e-20
C8134 XM1/a_100_n167894# XM2/a_n158_n321474# 0.114915f
C8135 XM1/a_n100_n96191# XM2/a_n158_n250302# 0.010147f
C8136 XM1/a_n100_117773# XM2/a_n158_n36786# 0.010147f
C8137 XM1/a_100_n172202# XM4/w_n358_n132787# 0.048442f
C8138 XM2/a_n100_n179227# XM3/a_n100_27993# 6.21e-19
C8139 XM2/a_n100_n7887# XM1/a_100_145154# 0.005074f
C8140 XM4/w_n358_n132787# XM3/a_n158_n13350# 0.032295f
C8141 XM1/a_n100_155109# XM2/a_100_2754# 7.26e-20
C8142 XM4/a_100_n130418# XM2/a_n100_n334751# 2.56e-20
C8143 XM1/a_100_n8498# XM3/a_n100_43533# 2.85e-20
C8144 XM1/a_n158_80534# XM3/a_n100_131593# 1.94e-20
C8145 XM2/a_n100_n13159# XM1/a_100_142282# 0.005074f
C8146 XM2/a_n158_n13062# XM1/a_n100_140749# 0.010147f
C8147 XM1/a_n158_110690# XM2/a_n100_n42155# 7.26e-20
C8148 XM1/a_100_33146# XM4/w_n358_n132787# 0.048442f
C8149 XM2/a_n158_n173858# XM3/a_n158_33270# 4.64e-21
C8150 XM4/a_n100_32137# m1_1634_n2388# 0.072015f
C8151 XM2/a_n100_23745# XM1/a_100_179618# 0.005074f
C8152 XM1/a_n158_57558# XM3/a_n100_109837# 1.02e-20
C8153 avdd pbias 0.041634f
C8154 XM1/a_100_n170766# XM3/a_n100_n120155# 2.85e-20
C8155 XM4/w_n358_n132787# XM3/a_n100_n117047# 0.009186f
C8156 XM4/a_100_n102446# m1_1634_n2388# 6.1e-20
C8157 XM2/a_n158_n105322# m1_1634_n2388# 2.36e-21
C8158 XM1/a_100_18786# XM3/a_n100_69433# 0.001033f
C8159 XM2/a_100_n279298# XM3/a_n158_n74474# 0.077916f
C8160 XM1/a_100_n84606# XM2/a_n158_n239758# 0.082589f
C8161 XM3/a_n100_46641# m1_1634_n2388# 0.072015f
C8162 XM1/a_n100_n176607# XM3/a_n100_n125335# 3.25e-19
C8163 XM1/a_100_n109018# XM3/a_n100_n56959# 2.85e-20
C8164 XM2/a_100_n321474# XM3/a_n100_n116011# 0.010147f
C8165 XM1/a_100_n41526# XM3/a_n100_10381# 2.85e-20
C8166 XM4/w_n358_n132787# XM2/a_n100_n173955# 0.025738f
C8167 XM2/a_n100_n292575# m1_1634_n2388# 7.61e-19
C8168 XM1/a_100_63302# m1_1634_n2388# 7.88e-19
C8169 XM2/a_n100_n318935# XM3/a_n158_n114878# 0.004271f
C8170 XM4/w_n358_n132787# XM4/a_n100_126413# -0.004445f
C8171 XM4/w_n358_n132787# XM3/a_n158_88178# 0.038462f
C8172 XM1/a_n100_7201# XM3/a_n158_59170# 3.16e-19
C8173 XM1/a_100_n163586# XM2/a_n158_n318838# 0.072853f
C8174 XM2/a_n158_n231850# XM3/a_n100_n27951# 6.96e-20
C8175 XM4/w_n358_n132787# XM3/a_n100_124341# 0.00895f
C8176 XM4/w_n358_n132787# XM3/a_n158_n52718# 0.032295f
C8177 XM4/a_n100_n39347# m1_1634_n2388# 0.072015f
C8178 XM1/a_n100_163725# XM2/a_n158_8026# 0.005074f
C8179 XM4/w_n358_n132787# XM3/a_n158_33270# 0.038462f
C8180 XM2/a_n158_n316202# XM3/a_n158_n109698# 4.64e-21
C8181 XM1/a_100_100638# XM2/a_n158_n55238# 0.012096f
C8182 XM1/a_100_n91786# XM2/a_100_n247666# 4.64e-21
C8183 XM1/a_n158_n84606# XM2/a_n100_n237219# 7.26e-20
C8184 XM2/a_100_n229214# XM3/a_n100_n22771# 0.005074f
C8185 XM1/a_100_93458# XM2/a_n158_n60510# 0.116862f
C8186 XM2/a_100_n89506# XM3/a_n100_116053# 0.010147f
C8187 XM2/a_n158_n205490# XM3/a_n100_n1015# 7.26e-20
C8188 XM1/a_n100_170905# XM2/a_100_15934# 7.26e-20
C8189 XM1/a_n100_n67471# m1_1634_n2388# 1.3e-19
C8190 XM1/a_n158_89150# XM2/a_n158_n65782# 4.64e-21
C8191 XM2/a_n100_n158139# XM3/a_n158_46738# 4.08e-19
C8192 XM1/a_100_152334# XM2/a_n100_n2615# 0.001809f
C8193 XM1/a_n100_73257# XM2/a_n158_n78962# 4.8e-19
C8194 XM1/a_100_n180818# XM4/w_n358_n132787# 0.048442f
C8195 XM2/a_n100_n79059# XM4/a_100_127546# 2.56e-20
C8196 XM1/a_n158_n146354# XM3/a_n100_n95291# 1.94e-20
C8197 XM4/w_n358_n132787# XM2/a_n158_n110594# 0.106111f
C8198 XM4/w_n358_n132787# XM4/a_n100_87045# -0.004445f
C8199 XM1/a_n100_n165119# XM2/a_n158_n318838# 0.010147f
C8200 XM3/a_n100_n19663# m1_1634_n2388# 0.072015f
C8201 XM4/w_n358_n132787# XM2/a_n100_n297847# 0.025738f
C8202 XM1/a_n158_94894# XM2/a_n158_n57874# 4.64e-21
C8203 XM3/a_n158_71602# m1_1634_n2388# 6.1e-20
C8204 XM4/w_n358_n132787# XM3/a_n158_n92086# 0.032295f
C8205 XM4/a_n100_n78715# m1_1634_n2388# 0.072015f
C8206 XM2/a_n100_n266215# XM4/a_100_n62042# 2.56e-20
C8207 XM3/a_n158_102682# m1_1634_n2388# 6.1e-20
C8208 XM2/a_100_n303022# XM3/a_n100_n98399# 0.005074f
C8209 XM1/a_100_n100402# XM4/w_n358_n132787# 0.054609f
C8210 XM1/a_n100_n33007# XM2/a_n158_n187038# 0.010147f
C8211 XM1/a_n158_166694# XM2/a_n100_13201# 7.26e-20
C8212 XM1/a_100_13042# XM2/a_n100_n139687# 0.005074f
C8213 XM1/a_n100_n145015# XM2/a_n158_n300386# 0.005074f
C8214 XM1/a_n100_n109115# XM3/a_n100_n57995# 1.19e-19
C8215 XM1/a_n100_n96191# XM3/a_n158_n45466# 2.85e-20
C8216 XM3/a_n158_16694# m1_1634_n2388# 6.1e-20
C8217 XM3/a_n100_40425# XM4/a_n100_40425# 0.009521f
C8218 XM1/a_100_n107582# XM2/a_100_n260846# 4.64e-21
C8219 XM4/a_100_121330# m1_1634_n2388# 6.1e-20
C8220 XM1/a_n158_40326# XM3/a_n100_91189# 1.94e-20
C8221 XM1/a_n100_n45931# XM3/a_n158_5298# 2.08e-20
C8222 XM2/a_n100_n152867# XM4/a_100_51918# 2.56e-20
C8223 XM1/a_100_158078# XM2/a_n158_5390# 0.028064f
C8224 XM1/a_100_8734# XM2/a_n100_n144959# 8.54e-20
C8225 XM1/a_n100_n4287# m1_1634_n2388# 1.3e-19
C8226 XM2/a_100_n210762# XM3/a_n100_n5159# 0.010147f
C8227 XM1/a_n100_n25827# XM2/a_100_n181766# 4.56e-20
C8228 XM4/w_n358_n132787# XM4/a_n100_47677# -0.004445f
C8229 XM1/a_100_n44398# XM3/a_n158_6334# 0.003891f
C8230 XM3/a_n100_n59031# m1_1634_n2388# 0.072015f
C8231 XM2/a_n100_n208223# XM3/a_n158_n4026# 0.005074f
C8232 XM1/a_100_50378# XM2/a_n100_n102783# 0.005074f
C8233 XM1/a_100_40326# XM4/w_n358_n132787# 0.049726f
C8234 XM1/a_n100_7201# XM2/a_n100_n147595# 0.006262f
C8235 XM1/a_n100_n137835# XM3/a_n158_n86906# 2.85e-20
C8236 XM2/a_100_n165950# m1_1634_n2388# 0.017213f
C8237 XM2/a_n100_n250399# XM3/a_n100_n45563# 0.003389f
C8238 XM4/w_n358_n132787# XM3/a_n158_n131454# 0.032295f
C8239 XM4/a_n100_n118083# m1_1634_n2388# 0.072015f
C8240 XM3/a_n100_n11375# XM4/a_n100_n11375# 0.009521f
C8241 XM4/w_n358_n132787# XM2/a_n158_n234486# 0.107093f
C8242 XM1/a_n100_38793# XM2/a_n158_n115866# 0.006179f
C8243 XM1/a_100_119306# XM2/a_n158_n34150# 0.102841f
C8244 XM2/a_100_n134318# XM3/a_n100_70469# 0.009693f
C8245 XM1/a_n100_n178043# XM2/a_100_n332018# 1.45e-19
C8246 XM1/a_n158_n75990# XM2/a_n100_n231947# 7.26e-20
C8247 XM4/w_n358_n132787# XM3/a_n158_100610# 0.032295f
C8248 XM1/a_100_n167894# XM2/a_n100_n321571# 4.08e-19
C8249 XM4/w_n358_n132787# XM4/a_n100_n23807# -0.004445f
C8250 XM1/a_n100_n5723# XM2/a_100_n158042# 7.26e-20
C8251 XM1/a_n100_21# XM4/w_n358_n132787# 0.01363f
C8252 XM1/a_n100_107721# XM4/w_n358_n132787# 0.012279f
C8253 XM1/a_100_n173638# XM2/a_100_n329382# 4.64e-21
C8254 XM1/a_100_n106146# XM2/a_n158_n260846# 0.116862f
C8255 XM2/a_100_n176494# XM3/a_n100_27993# 0.005074f
C8256 XM4/a_100_81962# m1_1634_n2388# 6.1e-20
C8257 XM1/a_n158_113562# XM2/a_n100_n39519# 7.26e-20
C8258 XM1/a_100_n54450# XM3/a_n100_n2051# 1.09e-21
C8259 XM1/a_n100_n47367# XM3/a_n100_4165# 2.09e-19
C8260 XM1/a_n100_20125# XM3/a_n100_72541# 2.08e-19
C8261 XM1/a_n100_n55983# XM4/w_n358_n132787# 0.014293f
C8262 XM1/a_n100_n30135# XM3/a_n158_21874# 2.85e-20
C8263 XM1/a_n100_n120603# XM3/a_n158_n68258# 2.85e-20
C8264 XM1/a_100_n68810# XM3/a_n158_n17494# 0.001549f
C8265 XM1/a_100_20222# XM3/a_n100_70469# 1.29e-20
C8266 XM3/a_n100_n98399# m1_1634_n2388# 0.072015f
C8267 XM1/a_n158_n93222# XM2/a_n158_n247666# 9.28e-21
C8268 XM2/a_n100_n173955# XM3/a_n158_33270# 0.005074f
C8269 XM3/a_n100_n31059# XM4/a_n100_n31059# 0.009521f
C8270 XM2/a_n100_n105419# m1_1634_n2388# 0.001564f
C8271 XM4/w_n358_n132787# XM3/a_n100_81865# 0.009011f
C8272 XM1/a_n158_n106146# XM2/a_n158_n260846# 9.28e-21
C8273 XM1/a_100_n84606# XM2/a_n100_n239855# 0.005074f
C8274 XM1/a_n100_n60291# XM4/w_n358_n132787# 0.01363f
C8275 XM1/a_100_n47270# XM2/a_100_n202854# 4.64e-21
C8276 XM2/a_n158_n321474# XM3/a_n100_n116011# 1.45e-19
C8277 XM1/a_n158_n107582# XM3/a_n100_n55923# 1.94e-20
C8278 XM4/w_n358_n132787# XM3/a_n100_n4123# 0.009186f
C8279 XM4/w_n358_n132787# XM2/a_100_n171222# 0.103341f
C8280 XM2/a_100_n289842# m1_1634_n2388# 0.024149f
C8281 XM4/w_n358_n132787# XM3/a_n100_26957# 0.009186f
C8282 XM4/w_n358_n132787# XM4/a_n100_n63175# -0.004445f
C8283 XM1/a_100_n87478# XM3/a_n100_n35203# 0.001448f
C8284 XM2/a_n158_n20970# XM1/a_100_132230# 0.077916f
C8285 XM2/a_100_n121138# XM3/a_n100_84973# 0.010147f
C8286 XM1/a_100_n163586# XM2/a_n100_n318935# 0.005074f
C8287 XM3/a_n158_n34070# m1_1634_n2388# 6.1e-20
C8288 XM2/a_n100_n231947# XM3/a_n100_n27951# 1.24e-19
C8289 XM1/a_100_127922# XM4/w_n358_n132787# 0.048442f
C8290 XM1/a_100_30274# XM4/w_n358_n132787# 0.048442f
C8291 XM4/a_100_42594# m1_1634_n2388# 6.1e-20
C8292 XM1/a_n100_n166555# XM3/a_n158_n115914# 2.85e-20
C8293 XM2/a_100_n163314# XM3/a_n100_42497# 0.010147f
C8294 XM2/a_n100_n316299# XM3/a_n158_n109698# 0.005074f
C8295 XM1/a_n158_n104710# XM3/a_n158_n53754# 1.14e-21
C8296 XM1/a_100_n91786# XM2/a_n158_n247666# 0.011707f
C8297 XM2/a_n158_n229214# XM3/a_n100_n22771# 7.26e-20
C8298 XM2/a_n158_n89506# XM3/a_n100_116053# 1.45e-19
C8299 XM2/a_n158_n55238# XM4/w_n358_n132787# 0.107093f
C8300 XM3/a_n100_n50743# XM4/a_n100_n50743# 0.009521f
C8301 XM1/a_n100_73257# XM2/a_n100_n79059# 0.004047f
C8302 XM1/a_n100_162289# XM2/a_n158_8026# 0.010147f
C8303 XM4/a_n100_105693# m1_1634_n2388# 0.072015f
C8304 XM4/w_n358_n132787# XM3/a_n100_n43491# 0.009081f
C8305 XM4/a_100_n28890# m1_1634_n2388# 6.1e-20
C8306 XM1/a_n100_21561# XM2/a_100_n131682# 7.26e-20
C8307 XM3/a_n100_65289# m1_1634_n2388# 0.072015f
C8308 XM2/a_n100_n313663# XM4/a_n100_n109795# 3.39e-21
C8309 XM1/a_100_n44398# XM2/a_100_n200218# 4.64e-21
C8310 XM1/a_100_163822# XM2/a_100_10662# 4.64e-21
C8311 XM1/a_n158_n152098# XM3/a_n100_n100471# 1.94e-20
C8312 XM1/a_n158_97766# XM2/a_n158_n55238# 4.64e-21
C8313 XM4/w_n358_n132787# XM2/a_n100_n110691# 0.024134f
C8314 XM1/a_n158_n156406# XM2/a_n158_n310930# 9.28e-21
C8315 XM4/w_n358_n132787# XM4/a_n100_n102543# -0.004445f
C8316 XM2/a_n100_n229311# m1_1634_n2388# 7.61e-19
C8317 XM3/a_n100_7273# XM4/a_n100_7273# 0.009521f
C8318 XM3/a_n158_n73438# m1_1634_n2388# 6.1e-20
C8319 XM3/a_n100_10381# m1_1634_n2388# 0.072015f
C8320 XM1/a_n100_n137835# XM4/w_n358_n132787# 0.013537f
C8321 XM3/a_n100_93261# XM4/a_n100_93261# 0.009521f
C8322 XM4/w_n358_n132787# XM2/a_100_n295114# 0.10657f
C8323 XM3/a_n100_102585# m1_1634_n2388# 0.072015f
C8324 XM2/a_n158_n303022# XM3/a_n100_n98399# 7.26e-20
C8325 XM1/a_100_n123378# XM3/a_n158_n72402# 0.00544f
C8326 XM4/w_n358_n132787# XM3/a_n158_51918# 0.035059f
C8327 XM2/a_100_n150134# XM3/a_n100_57001# 0.004433f
C8328 XM4/a_n100_n131551# m1_1634_n2388# 0.072015f
C8329 XM2/a_100_n258210# XM3/a_n158_n51682# 0.065453f
C8330 XM1/a_n100_n35879# m1_1634_n2388# 7.88e-20
C8331 XM1/a_100_n146354# XM3/a_n100_n95291# 2.85e-20
C8332 XM4/w_n358_n132787# XM1/a_n100_n136399# 0.014176f
C8333 XM2/a_n100_n263579# XM4/a_100_n56862# 2.56e-20
C8334 XM1/a_100_n67374# XM3/a_n100_n15519# 2.85e-20
C8335 XM2/a_100_n192310# XM3/a_n100_14525# 0.005074f
C8336 XM1/a_n158_n21422# XM3/a_n100_29029# 1.94e-20
C8337 XM2/a_100_n300386# XM3/a_n100_n93219# 0.002238f
C8338 XM3/a_n100_n70427# XM4/a_n100_n70427# 0.009521f
C8339 XM1/a_100_n107582# XM2/a_n158_n260846# 0.084147f
C8340 XM4/a_n100_66325# m1_1634_n2388# 0.072015f
C8341 XM4/w_n358_n132787# XM3/a_n100_n82859# 0.009186f
C8342 XM4/a_100_n68258# m1_1634_n2388# 6.1e-20
C8343 XM2/a_n158_n210762# XM3/a_n100_n5159# 1.45e-19
C8344 XM1/a_n100_n25827# XM2/a_n158_n181766# 0.004352f
C8345 XM1/a_n158_n93222# XM3/a_n100_n41419# 1.94e-20
C8346 XM3/a_n158_n112806# m1_1634_n2388# 6.1e-20
C8347 XM1/a_n100_86181# XM2/a_n158_n68418# 0.010147f
C8348 XM1/a_n100_27305# XM3/a_n158_77818# 2.85e-20
C8349 XM1/a_100_n40090# XM3/a_n100_11417# 2.85e-20
C8350 XM1/a_n158_2990# XM2/a_n158_n152770# 4.64e-21
C8351 XM2/a_n100_n150231# XM4/a_100_57098# 1.71e-20
C8352 XM1/a_100_158078# XM4/w_n358_n132787# 0.053546f
C8353 XM4/w_n358_n132787# XM2/a_n100_n234583# 0.025738f
C8354 XM1/a_n100_38793# XM2/a_n100_n115963# 0.002599f
C8355 XM3/a_n158_90250# m1_1634_n2388# 6.1e-20
C8356 XM1/a_100_n149226# XM4/w_n358_n132787# 0.048442f
C8357 XM1/a_n100_n61727# XM4/w_n358_n132787# 0.013401f
C8358 XM1/a_100_n50142# XM4/w_n358_n132787# 0.054609f
C8359 XM3/a_n158_127546# m1_1634_n2388# 6.1e-20
C8360 XM2/a_100_n332018# XM3/a_n158_n127310# 0.068958f
C8361 XM1/a_n100_n160811# m1_1634_n2388# 1.3e-19
C8362 XM4/w_n358_n132787# XM3/a_n158_n18530# 0.032295f
C8363 XM4/a_n100_n5159# m1_1634_n2388# 0.072015f
C8364 XM1/a_n158_79098# XM2/a_n100_n73787# 7.26e-20
C8365 XM3/a_n100_4165# m1_1634_n2388# 0.072015f
C8366 XM2/a_n158_n134318# XM3/a_n100_70469# 1.38e-19
C8367 XM1/a_n100_n178043# XM2/a_n158_n332018# 0.010147f
C8368 XM2/a_n100_n247763# XM3/a_n100_n40383# 5.6e-19
C8369 XM3/a_n158_35342# m1_1634_n2388# 6.1e-20
C8370 XM4/w_n358_n132787# XM3/a_n100_100513# 0.009042f
C8371 XM1/a_n100_n142143# m1_1634_n2388# 1.3e-19
C8372 XM1/a_n158_n73118# XM2/a_n100_n229311# 7.48e-22
C8373 XM1/a_n100_n172299# XM2/a_100_n326746# 1.45e-19
C8374 XM3/a_n100_n90111# XM4/a_n100_n90111# 0.009521f
C8375 XM1/a_100_n34346# XM3/a_n100_16597# 0.001195f
C8376 XM1/a_n100_n5723# XM2/a_n158_n158042# 0.005074f
C8377 XM1/a_100_n173638# XM2/a_n158_n329382# 0.024949f
C8378 XM1/a_n100_n149323# XM2/a_100_n303022# 1.45e-19
C8379 XM4/a_n100_26957# m1_1634_n2388# 0.072015f
C8380 XM2/a_n158_n176494# XM3/a_n100_27993# 7.26e-20
C8381 XM1/a_n100_30177# XM3/a_n158_80926# 2.85e-20
C8382 XM1/a_n158_20222# XM3/a_n100_71505# 3.89e-20
C8383 XM1/a_n158_n9934# XM2/a_n100_n166047# 6.06e-20
C8384 XM4/w_n358_n132787# XM3/a_n100_n122227# 0.008296f
C8385 XM4/a_100_n107626# m1_1634_n2388# 6.1e-20
C8386 XM1/a_100_57558# m1_1634_n2388# 0.002487f
C8387 XM2/a_100_n129046# XM3/a_n158_75746# 0.077137f
C8388 XM1/a_100_n25730# XM3/a_n100_25921# 2.85e-20
C8389 XM1/a_100_51814# XM3/a_n100_102585# 2.85e-20
C8390 XM1/a_n100_n180915# XM3/a_n100_n128443# 9.37e-19
C8391 XM1/a_100_n91786# XM3/a_n100_n41419# 0.00117f
C8392 XM2/a_100_n239758# XM3/a_n158_n34070# 0.077916f
C8393 XM2/a_100_n171222# XM3/a_n158_33270# 0.047927f
C8394 XM2/a_100_n281934# XM3/a_n100_n75607# 0.005074f
C8395 XM4/w_n358_n132787# XM4/a_n100_121233# -0.004445f
C8396 XM1/a_n100_109157# XM4/w_n358_n132787# 0.012279f
C8397 XM2/a_100_n102686# m1_1634_n2388# 0.017213f
C8398 XM1/a_100_n84606# XM2/a_100_n237122# 4.64e-21
C8399 XM1/a_n100_100541# XM2/a_100_n55238# 7.26e-20
C8400 XM1/a_100_n47270# XM2/a_n158_n202854# 0.040527f
C8401 XM4/w_n358_n132787# XM3/a_n158_n57898# 0.032295f
C8402 XM4/a_n100_n44527# m1_1634_n2388# 0.072015f
C8403 XM4/w_n358_n132787# XM2/a_n158_n171222# 0.107093f
C8404 XM2/a_n158_n289842# m1_1634_n2388# 2.36e-21
C8405 XM1/a_100_7298# XM3/a_n100_59073# 2.85e-20
C8406 XM1/a_100_n37218# XM3/a_n158_14622# 0.00544f
C8407 XM1/a_n100_n182351# sw_b 0.003226f
C8408 XM2/a_n158_n121138# XM3/a_n100_84973# 1.45e-19
C8409 XM1/a_100_n163586# XM2/a_100_n316202# 4.64e-21
C8410 XM3/a_n100_n109795# XM4/a_n100_n109795# 0.009521f
C8411 XM1/a_n158_n68810# XM2/a_n158_n223942# 4.64e-21
C8412 XM4/w_n358_n132787# XM3/a_n158_125474# 0.038543f
C8413 XM2/a_n100_n71151# XM4/w_n358_n132787# 0.012279f
C8414 XM2/a_n158_n163314# XM3/a_n100_42497# 1.45e-19
C8415 XM1/a_n100_n159375# XM3/a_n158_n107626# 1.61e-20
C8416 XM1/a_n100_n175171# XM3/a_n158_n123166# 2.85e-20
C8417 XM2/a_n100_n318935# XM4/a_100_n114878# 1.5e-20
C8418 XM1/a_n100_n86139# XM4/w_n358_n132787# 0.01363f
C8419 XM2/a_100_n115866# XM3/a_n158_90250# 0.077916f
C8420 XM1/a_100_n91786# XM2/a_n100_n247763# 0.005074f
C8421 XM2/a_100_n89506# XM3/a_n158_117186# 0.049485f
C8422 XM4/w_n358_n132787# XM4/a_n100_81865# -0.004445f
C8423 XM1/a_n158_n30038# XM2/a_n158_n184402# 9.28e-21
C8424 XM2/a_100_n158042# XM3/a_n158_47774# 0.077916f
C8425 XM3/a_n100_61145# XM4/a_n100_61145# 0.009521f
C8426 XM3/a_n100_n24843# m1_1634_n2388# 0.072015f
C8427 XM2/a_100_21206# XM1/a_n100_176649# 7.26e-20
C8428 XM1/a_n100_n149323# m1_1634_n2388# 1.3e-19
C8429 XM4/w_n358_n132787# XM3/a_n158_n97266# 0.032295f
C8430 XM4/a_n100_n83895# m1_1634_n2388# 0.072015f
C8431 XM1/a_n100_126389# XM2/a_100_n26242# 7.26e-20
C8432 XM1/a_n100_21561# XM2/a_n158_n131682# 0.005074f
C8433 XM1/a_100_n44398# XM2/a_n158_n200218# 0.017549f
C8434 XM2/a_100_n221306# XM3/a_n158_n16458# 0.077916f
C8435 XM1/a_100_133666# XM2/a_n158_n20970# 0.116862f
C8436 XM4/w_n358_n132787# XM2/a_100_n107958# 0.103341f
C8437 XM1/a_n100_n178043# XM3/a_n100_n126371# 3.25e-19
C8438 XM1/a_n100_n150759# XM2/a_100_n305658# 7.26e-20
C8439 XM1/a_100_n93222# XM3/a_n100_n42455# 2.85e-20
C8440 XM2/a_100_n226578# m1_1634_n2388# 0.022835f
C8441 XM4/w_n358_n132787# XM3/a_n100_45605# 0.00823f
C8442 XM3/a_n100_n129479# XM4/a_n100_n129479# 0.009521f
C8443 XM2/a_100_n263482# XM3/a_n100_n57995# 0.010147f
C8444 XM2/a_n100_n105419# XM3/a_n100_98441# 0.004495f
C8445 XM1/a_n158_n169330# XM3/a_n100_n118083# 3.89e-20
C8446 XM4/w_n358_n132787# XM2/a_n158_n295114# 0.107093f
C8447 XM2/a_n100_n260943# XM3/a_n158_n56862# 0.004756f
C8448 XM1/a_n100_123517# XM2/a_n158_n31514# 0.005074f
C8449 XM4/a_100_5298# m1_1634_n2388# 6.1e-20
C8450 XM2/a_n100_n303119# XM3/a_n100_n98399# 4.1e-19
C8451 XM1/a_n100_n145015# XM2/a_100_n297750# 7.26e-20
C8452 XM1/a_100_n37218# XM4/w_n358_n132787# 0.054609f
C8453 XM4/a_100_116150# m1_1634_n2388# 6.1e-20
C8454 XM2/a_n158_n150134# XM3/a_n100_57001# 4.86e-20
C8455 XM1/a_n100_n1415# m1_1634_n2388# 8.88e-20
C8456 XM2/a_n158_n258210# XM3/a_n158_n51682# 4.64e-21
C8457 XM4/w_n358_n132787# XM4/a_n100_42497# -0.004445f
C8458 XM1/a_n158_n116198# XM3/a_n100_n64211# 4.21e-21
C8459 XM2/a_n158_n192310# XM3/a_n100_14525# 7.26e-20
C8460 XM2/a_n158_n7790# XM4/w_n358_n132787# 0.107093f
C8461 XM2/a_n158_n300386# XM3/a_n100_n93219# 2.87e-20
C8462 XM3/a_n100_n64211# m1_1634_n2388# 0.072014f
C8463 XM1/a_100_44634# XM4/w_n358_n132787# 0.054609f
C8464 XM1/a_100_n107582# XM2/a_n100_n260943# 0.005074f
C8465 XM2/a_100_n144862# XM3/a_n158_62278# 0.005865f
C8466 XM4/a_n100_n123263# m1_1634_n2388# 0.072015f
C8467 XM1/a_100_66174# XM2/a_100_n89506# 4.64e-21
C8468 XM1/a_n100_n25827# XM2/a_n100_n181863# 0.001118f
C8469 XM3/a_n100_83937# m1_1634_n2388# 0.072015f
C8470 XM1/a_n100_n162247# XM3/a_n100_n109795# 6.76e-19
C8471 XM1/a_n158_n54450# XM3/a_n100_n4123# 1.94e-20
C8472 XM2/a_100_n187038# XM3/a_n158_19802# 0.035075f
C8473 XM1/a_n158_n104710# XM2/a_n158_n258210# 4.64e-21
C8474 XM1/a_100_44634# XM2/a_100_n110594# 4.64e-21
C8475 XM3/a_n100_n2051# m1_1634_n2388# 0.072015f
C8476 XM2/a_n100_n166047# m1_1634_n2388# 0.001582f
C8477 XM1/a_n158_168130# XM2/a_n100_13201# 2.39e-20
C8478 XM3/a_n100_29029# m1_1634_n2388# 0.072015f
C8479 XM1/a_n158_2990# XM2/a_n100_n152867# 7.26e-20
C8480 XM4/w_n358_n132787# XM4/a_n100_n28987# -0.004445f
C8481 XM3/a_n100_119161# XM4/a_n100_119161# 0.009521f
C8482 XM4/w_n358_n132787# XM2/a_100_n231850# 0.106552f
C8483 XM2/a_100_n205490# XM3/a_n100_21# 0.010147f
C8484 XM3/a_n100_127449# m1_1634_n2388# 0.072015f
C8485 XM4/a_100_76782# m1_1634_n2388# 6.1e-20
C8486 XM2/a_n158_n332018# XM3/a_n158_n127310# 4.64e-21
C8487 XM2/a_n100_n208223# XM4/a_100_n4026# 2.56e-20
C8488 XM1/a_100_61866# XM2/a_n158_n92142# 0.116862f
C8489 XM2/a_n100_n134415# XM3/a_n100_70469# 4.51e-19
C8490 XM4/w_n358_n132787# XM3/a_n158_70566# 0.032295f
C8491 XM2/a_100_n245030# XM3/a_n100_n40383# 0.005074f
C8492 XM1/a_n158_n75990# XM2/a_n158_n229214# 4.64e-21
C8493 XM1/a_100_n84606# XM3/a_n100_n33131# 3.76e-20
C8494 XM1/a_n100_n172299# XM2/a_n158_n326746# 0.010147f
C8495 XM3/a_n100_n103579# m1_1634_n2388# 0.072015f
C8496 pbias XM4/w_n358_n132787# 0.003395f
C8497 XM1/a_100_n173638# XM2/a_n100_n329479# 0.005074f
C8498 XM1/a_n100_n149323# XM2/a_n158_n303022# 0.010147f
C8499 XM4/w_n358_n132787# XM3/a_n158_15658# 0.032295f
C8500 XM1/a_100_30274# XM3/a_n100_81865# 2.85e-20
C8501 XM2/a_n100_n284667# XM3/a_n100_n80787# 0.004878f
C8502 XM1/a_n100_n63163# XM2/a_100_n218670# 7.26e-20
C8503 XM2/a_n158_n129046# XM3/a_n158_75746# 4.64e-21
C8504 XM1/a_100_n81734# XM3/a_n100_n31059# 2.85e-20
C8505 XM2/a_n100_n94875# XM4/a_100_109934# 2.32e-20
C8506 XM4/w_n358_n132787# XM3/a_n100_n9303# 0.009109f
C8507 XM2/a_n158_n171222# XM3/a_n158_33270# 4.64e-21
C8508 XM1/a_100_153770# XM2/a_n158_118# 0.116862f
C8509 XM2/a_n158_n281934# XM3/a_n100_n75607# 7.26e-20
C8510 XM1/a_n100_n109115# XM2/a_100_n263482# 1.45e-19
C8511 XM4/w_n358_n132787# XM4/a_n100_n68355# -0.004445f
C8512 XM3/a_n158_n39250# m1_1634_n2388# 6.1e-20
C8513 XM1/a_100_n84606# XM2/a_n158_n237122# 0.011317f
C8514 XM1/a_100_n47270# XM2/a_n100_n202951# 0.005074f
C8515 XM4/a_100_37414# m1_1634_n2388# 6.1e-20
C8516 XM1/a_n158_n162150# XM3/a_n100_n111867# 1.54e-20
C8517 XM4/w_n358_n132787# XM2/a_n100_n171319# 0.025738f
C8518 XM1/a_100_107818# XM2/a_n100_n47427# 0.005074f
C8519 XM2/a_n100_n289939# m1_1634_n2388# 8.98e-19
C8520 XM1/a_n100_21# XM3/a_n158_51918# 2.85e-20
C8521 XM1/a_n100_n94755# XM2/a_100_n250302# 7.26e-20
C8522 XM1/a_100_n126250# XM3/a_n100_n75607# 9.77e-19
C8523 XM1/a_n100_n1415# XM3/a_n158_49846# 1.14e-20
C8524 XM1/a_100_n163586# XM2/a_n158_n316202# 0.021054f
C8525 XM1/a_n158_n68810# XM2/a_n100_n224039# 7.26e-20
C8526 XM3/a_n158_53990# m1_1634_n2388# 6.1e-20
C8527 XM4/w_n358_n132787# XM3/a_n100_125377# 0.009186f
C8528 XM3/a_n100_29029# XM4/a_n100_29029# 0.009521f
C8529 XM1/a_100_n160714# m1_1634_n2388# 0.002487f
C8530 XM4/a_n100_100513# m1_1634_n2388# 0.072015f
C8531 XM4/w_n358_n132787# XM3/a_n100_n48671# 0.00916f
C8532 XM1/a_100_n91786# XM2/a_100_n245030# 4.64e-21
C8533 XM4/a_100_n34070# m1_1634_n2388# 6.1e-20
C8534 XM2/a_100_n226578# XM3/a_n100_n22771# 2.49e-20
C8535 XM2/a_n158_n89506# XM3/a_n158_117186# 4.64e-21
C8536 XM2/a_100_n89506# XM3/a_n100_117089# 0.005074f
C8537 XM3/a_n100_102585# XM4/a_n100_102585# 0.009521f
C8538 XM4/w_n358_n132787# XM4/a_n100_n107723# -0.004445f
C8539 XM2/a_100_n310930# XM3/a_n158_n104518# 0.076747f
C8540 XM3/a_n158_n78618# m1_1634_n2388# 6.1e-20
C8541 XM1/a_100_54686# XM4/w_n358_n132787# 0.048442f
C8542 XM2/a_n100_n316299# XM4/a_100_n109698# 2.56e-20
C8543 XM4/w_n358_n132787# XM1/a_n100_n145015# 0.01363f
C8544 XM1/a_n100_89053# XM2/a_n158_n65782# 0.005074f
C8545 XM4/a_n100_n1015# m1_1634_n2388# 0.072015f
C8546 XM1/a_100_n44398# XM2/a_n100_n200315# 0.005074f
C8547 XM4/w_n358_n132787# XM2/a_n158_n107958# 0.107093f
C8548 XM1/a_n100_n150759# XM2/a_n158_n305658# 0.005074f
C8549 XM2/a_n158_n226578# m1_1634_n2388# 2.36e-21
C8550 XM1/a_n158_n70246# XM3/a_n100_n19663# 1.94e-20
C8551 XM2/a_n158_n263482# XM3/a_n100_n57995# 1.45e-19
C8552 XM1/a_n158_132230# XM2/a_n100_n23703# 7.26e-20
C8553 XM4/w_n358_n132787# XM2/a_n100_n295211# 0.025738f
C8554 XM2/a_n100_n23703# XM4/w_n358_n132787# 0.012279f
C8555 XM3/a_n158_103718# m1_1634_n2388# 6.1e-20
C8556 XM2/a_n100_n13159# XM1/a_n158_142282# 7.26e-20
C8557 XM1/a_100_51814# XM2/a_n158_n102686# 0.116862f
C8558 XM1/a_n100_n145015# XM2/a_n158_n297750# 0.005074f
C8559 XM4/a_n100_61145# m1_1634_n2388# 0.072015f
C8560 XM2/a_n100_n150231# XM3/a_n100_57001# 9.94e-19
C8561 XM1/a_n100_n173735# XM3/a_n158_n123166# 2.85e-20
C8562 XM4/w_n358_n132787# XM3/a_n100_n88039# 0.008979f
C8563 XM4/a_100_n73438# m1_1634_n2388# 6.1e-20
C8564 XM1/a_n100_n111987# XM2/a_100_n266118# 1.45e-19
C8565 XM1/a_n100_11509# XM2/a_100_n142226# 1.45e-19
C8566 XM1/a_n100_43101# XM3/a_n158_95430# 2.85e-20
C8567 XM2/a_n100_n258307# XM3/a_n158_n51682# 0.005074f
C8568 XM1/a_100_n103274# XM3/a_n100_n52815# 2.85e-20
C8569 XM1/a_100_n71682# XM3/a_n100_n19663# 2.85e-20
C8570 XM1/a_n158_n60194# XM3/a_n100_n8267# 1.94e-20
C8571 XM3/a_n158_n117986# m1_1634_n2388# 6.1e-20
C8572 XM2/a_n100_n300483# XM3/a_n100_n93219# 0.002708f
C8573 XM2/a_n158_n144862# XM3/a_n158_62278# 4.64e-21
C8574 XM1/a_100_66174# XM2/a_n158_n89506# 0.03118f
C8575 XM1/a_n100_n25827# XM2/a_100_n179130# 7.26e-20
C8576 XM1/a_100_n177946# XM3/a_n100_n127407# 2.85e-20
C8577 XM1/a_100_n131994# XM4/w_n358_n132787# 0.054925f
C8578 XM1/a_n100_n99063# XM3/a_n100_n46599# 8.33e-19
C8579 XM2/a_n158_n187038# XM3/a_n158_19802# 4.64e-21
C8580 XM1/a_n100_150801# XM2/a_100_n2518# 7.26e-20
C8581 XM1/a_n100_57461# m1_1634_n2388# 2.27e-20
C8582 XM1/a_n158_38890# XM3/a_n100_91189# 1.94e-20
C8583 XM1/a_n158_n104710# XM2/a_n100_n258307# 7.26e-20
C8584 XM4/w_n358_n132787# XM3/a_n158_n23710# 0.032295f
C8585 XM4/a_n100_n10339# m1_1634_n2388# 0.072015f
C8586 XM1/a_100_44634# XM2/a_n158_n110594# 0.075189f
C8587 XM2/a_n100_n255671# XM4/a_n100_n51779# 3.63e-20
C8588 XM2/a_100_n163314# m1_1634_n2388# 0.019664f
C8589 XM4/w_n358_n132787# XM3/a_n100_64253# 0.008358f
C8590 XM2/a_100_n292478# XM3/a_n158_n86906# 0.077916f
C8591 XM2/a_100_n334654# XM3/a_n100_n128443# 0.010051f
C8592 XM4/w_n358_n132787# XM2/a_n158_n231850# 0.107093f
C8593 XM2/a_n158_n205490# XM3/a_n100_21# 1.45e-19
C8594 XM1/a_n100_175213# XM2/a_100_21206# 1.45e-19
C8595 XM4/w_n358_n132787# XM3/a_n100_9345# 0.009173f
C8596 XM4/a_n100_21777# m1_1634_n2388# 0.072015f
C8597 XM2/a_n100_23745# XM4/w_n358_n132787# 0.012279f
C8598 XM2/a_n100_n332115# XM3/a_n158_n127310# 0.004978f
C8599 XM4/w_n358_n132787# XM3/a_n100_n127407# 0.008861f
C8600 XM4/a_100_n112806# m1_1634_n2388# 6.1e-20
C8601 XM1/a_100_n22858# XM3/a_n100_27993# 2.85e-20
C8602 XM2/a_n158_n245030# XM3/a_n100_n40383# 7.26e-20
C8603 XM1/a_n158_n75990# XM2/a_n100_n229311# 7.26e-20
C8604 XM1/a_n158_n73118# XM2/a_n158_n226578# 4.64e-21
C8605 XM4/w_n358_n132787# XM3/a_n158_101646# 0.038462f
C8606 iout VSUBS 0.164168f
C8607 iout_n VSUBS 0.134714f
C8608 sw_bn VSUBS 0.132254f
C8609 sw_b VSUBS 0.131112f
C8610 pcbias VSUBS 0.125664f
C8611 pbias VSUBS 0.127514f
C8612 avdd VSUBS 0.157659f
C8613 XM4/a_100_n132490# VSUBS 0.196066f
C8614 XM4/a_n100_n132587# VSUBS 0.260213f
C8615 XM4/a_100_n131454# VSUBS 0.190616f
C8616 XM4/a_n100_n131551# VSUBS 0.216482f
C8617 XM4/a_100_n130418# VSUBS 0.190616f
C8618 m1_1634_n2388# VSUBS 43.597813f
C8619 XM4/a_n100_n130515# VSUBS 0.216482f
C8620 XM4/a_100_n129382# VSUBS 0.190616f
C8621 XM4/a_n100_n129479# VSUBS 0.216482f
C8622 XM4/a_100_n128346# VSUBS 0.190616f
C8623 XM4/a_n100_n128443# VSUBS 0.216482f
C8624 XM4/a_100_n127310# VSUBS 0.190616f
C8625 XM4/a_n100_n127407# VSUBS 0.216482f
C8626 XM4/a_100_n126274# VSUBS 0.190616f
C8627 XM4/a_n100_n126371# VSUBS 0.216482f
C8628 XM4/a_100_n125238# VSUBS 0.190616f
C8629 XM4/a_n100_n125335# VSUBS 0.216482f
C8630 XM4/a_100_n124202# VSUBS 0.190616f
C8631 XM4/a_n100_n124299# VSUBS 0.216482f
C8632 XM4/a_100_n123166# VSUBS 0.190616f
C8633 XM4/a_n100_n123263# VSUBS 0.216482f
C8634 XM4/a_100_n122130# VSUBS 0.190616f
C8635 XM4/a_n100_n122227# VSUBS 0.216482f
C8636 XM4/a_100_n121094# VSUBS 0.190616f
C8637 XM4/a_n100_n121191# VSUBS 0.216482f
C8638 XM4/a_100_n120058# VSUBS 0.190616f
C8639 XM4/a_n100_n120155# VSUBS 0.216482f
C8640 XM4/a_100_n119022# VSUBS 0.190616f
C8641 XM4/a_n100_n119119# VSUBS 0.216482f
C8642 XM4/a_100_n117986# VSUBS 0.190616f
C8643 XM4/a_n100_n118083# VSUBS 0.216482f
C8644 XM4/a_100_n116950# VSUBS 0.190616f
C8645 XM4/a_n100_n117047# VSUBS 0.216482f
C8646 XM4/a_100_n115914# VSUBS 0.190616f
C8647 XM4/a_n100_n116011# VSUBS 0.216482f
C8648 XM4/a_100_n114878# VSUBS 0.190616f
C8649 XM4/a_n100_n114975# VSUBS 0.216482f
C8650 XM4/a_100_n113842# VSUBS 0.190616f
C8651 XM4/a_n100_n113939# VSUBS 0.216482f
C8652 XM4/a_100_n112806# VSUBS 0.190616f
C8653 XM4/a_n100_n112903# VSUBS 0.216482f
C8654 XM4/a_100_n111770# VSUBS 0.190616f
C8655 XM4/a_n100_n111867# VSUBS 0.216482f
C8656 XM4/a_100_n110734# VSUBS 0.190616f
C8657 XM4/a_n100_n110831# VSUBS 0.216482f
C8658 XM4/a_100_n109698# VSUBS 0.190616f
C8659 XM4/a_n100_n109795# VSUBS 0.216482f
C8660 XM4/a_100_n108662# VSUBS 0.190616f
C8661 XM4/a_n100_n108759# VSUBS 0.216482f
C8662 XM4/a_100_n107626# VSUBS 0.190616f
C8663 XM4/a_n100_n107723# VSUBS 0.216482f
C8664 XM4/a_100_n106590# VSUBS 0.190616f
C8665 XM4/a_n100_n106687# VSUBS 0.216482f
C8666 XM4/a_100_n105554# VSUBS 0.190616f
C8667 XM4/a_n100_n105651# VSUBS 0.216482f
C8668 XM4/a_100_n104518# VSUBS 0.190616f
C8669 XM4/a_n100_n104615# VSUBS 0.216482f
C8670 XM4/a_100_n103482# VSUBS 0.190616f
C8671 XM4/a_n100_n103579# VSUBS 0.216482f
C8672 XM4/a_100_n102446# VSUBS 0.190616f
C8673 XM4/a_n100_n102543# VSUBS 0.216482f
C8674 XM4/a_100_n101410# VSUBS 0.190616f
C8675 XM4/a_n100_n101507# VSUBS 0.216482f
C8676 XM4/a_100_n100374# VSUBS 0.190616f
C8677 XM4/a_n100_n100471# VSUBS 0.216482f
C8678 XM4/a_100_n99338# VSUBS 0.190616f
C8679 XM4/a_n100_n99435# VSUBS 0.216482f
C8680 XM4/a_100_n98302# VSUBS 0.190616f
C8681 XM4/a_n100_n98399# VSUBS 0.216482f
C8682 XM4/a_100_n97266# VSUBS 0.190616f
C8683 XM4/a_n100_n97363# VSUBS 0.216482f
C8684 XM4/a_100_n96230# VSUBS 0.190616f
C8685 XM4/a_n100_n96327# VSUBS 0.216482f
C8686 XM4/a_100_n95194# VSUBS 0.190616f
C8687 XM4/a_n100_n95291# VSUBS 0.216482f
C8688 XM4/a_100_n94158# VSUBS 0.190616f
C8689 XM4/a_n100_n94255# VSUBS 0.216482f
C8690 XM4/a_100_n93122# VSUBS 0.190616f
C8691 XM4/a_n100_n93219# VSUBS 0.216482f
C8692 XM4/a_100_n92086# VSUBS 0.190616f
C8693 XM4/a_n100_n92183# VSUBS 0.216482f
C8694 XM4/a_100_n91050# VSUBS 0.190616f
C8695 XM4/a_n100_n91147# VSUBS 0.216482f
C8696 XM4/a_100_n90014# VSUBS 0.190616f
C8697 XM4/a_n100_n90111# VSUBS 0.216482f
C8698 XM4/a_100_n88978# VSUBS 0.190616f
C8699 XM4/a_n100_n89075# VSUBS 0.216482f
C8700 XM4/a_100_n87942# VSUBS 0.190616f
C8701 XM4/a_n100_n88039# VSUBS 0.216482f
C8702 XM4/a_100_n86906# VSUBS 0.190616f
C8703 XM4/a_n100_n87003# VSUBS 0.216482f
C8704 XM4/a_100_n85870# VSUBS 0.190616f
C8705 XM4/a_n100_n85967# VSUBS 0.216482f
C8706 XM4/a_100_n84834# VSUBS 0.190616f
C8707 XM4/a_n100_n84931# VSUBS 0.216482f
C8708 XM4/a_100_n83798# VSUBS 0.190616f
C8709 XM4/a_n100_n83895# VSUBS 0.216482f
C8710 XM4/a_100_n82762# VSUBS 0.190616f
C8711 XM4/a_n100_n82859# VSUBS 0.216482f
C8712 XM4/a_100_n81726# VSUBS 0.190616f
C8713 XM4/a_n100_n81823# VSUBS 0.216482f
C8714 XM4/a_100_n80690# VSUBS 0.190616f
C8715 XM4/a_n100_n80787# VSUBS 0.216482f
C8716 XM4/a_100_n79654# VSUBS 0.190616f
C8717 XM4/a_n100_n79751# VSUBS 0.216482f
C8718 XM4/a_100_n78618# VSUBS 0.190616f
C8719 XM4/a_n100_n78715# VSUBS 0.216482f
C8720 XM4/a_100_n77582# VSUBS 0.190616f
C8721 XM4/a_n100_n77679# VSUBS 0.216482f
C8722 XM4/a_100_n76546# VSUBS 0.190616f
C8723 XM4/a_n100_n76643# VSUBS 0.216482f
C8724 XM4/a_100_n75510# VSUBS 0.190616f
C8725 XM4/a_n100_n75607# VSUBS 0.216482f
C8726 XM4/a_100_n74474# VSUBS 0.190616f
C8727 XM4/a_n100_n74571# VSUBS 0.216482f
C8728 XM4/a_100_n73438# VSUBS 0.190616f
C8729 XM4/a_n100_n73535# VSUBS 0.216482f
C8730 XM4/a_100_n72402# VSUBS 0.190616f
C8731 XM4/a_n100_n72499# VSUBS 0.216482f
C8732 XM4/a_100_n71366# VSUBS 0.190616f
C8733 XM4/a_n100_n71463# VSUBS 0.216482f
C8734 XM4/a_100_n70330# VSUBS 0.190616f
C8735 XM4/a_n100_n70427# VSUBS 0.216482f
C8736 XM4/a_100_n69294# VSUBS 0.190616f
C8737 XM4/a_n100_n69391# VSUBS 0.216482f
C8738 XM4/a_100_n68258# VSUBS 0.190616f
C8739 XM4/a_n100_n68355# VSUBS 0.216482f
C8740 XM4/a_100_n67222# VSUBS 0.190616f
C8741 XM4/a_n100_n67319# VSUBS 0.216482f
C8742 XM4/a_100_n66186# VSUBS 0.190616f
C8743 XM4/a_n100_n66283# VSUBS 0.216482f
C8744 XM4/a_100_n65150# VSUBS 0.190616f
C8745 XM4/a_n100_n65247# VSUBS 0.216482f
C8746 XM4/a_100_n64114# VSUBS 0.190616f
C8747 XM4/a_n100_n64211# VSUBS 0.216482f
C8748 XM4/a_100_n63078# VSUBS 0.190616f
C8749 XM4/a_n100_n63175# VSUBS 0.216482f
C8750 XM4/a_100_n62042# VSUBS 0.190616f
C8751 XM4/a_n100_n62139# VSUBS 0.216482f
C8752 XM4/a_100_n61006# VSUBS 0.190616f
C8753 XM4/a_n100_n61103# VSUBS 0.216482f
C8754 XM4/a_100_n59970# VSUBS 0.190616f
C8755 XM4/a_n100_n60067# VSUBS 0.216482f
C8756 XM4/a_100_n58934# VSUBS 0.190616f
C8757 XM4/a_n100_n59031# VSUBS 0.216482f
C8758 XM4/a_100_n57898# VSUBS 0.190616f
C8759 XM4/a_n100_n57995# VSUBS 0.216482f
C8760 XM4/a_100_n56862# VSUBS 0.190616f
C8761 XM4/a_n100_n56959# VSUBS 0.216482f
C8762 XM4/a_100_n55826# VSUBS 0.190616f
C8763 XM4/a_n100_n55923# VSUBS 0.216482f
C8764 XM4/a_100_n54790# VSUBS 0.190616f
C8765 XM4/a_n100_n54887# VSUBS 0.216482f
C8766 XM4/a_100_n53754# VSUBS 0.190616f
C8767 XM4/a_n100_n53851# VSUBS 0.216482f
C8768 XM4/a_100_n52718# VSUBS 0.190616f
C8769 XM4/a_n100_n52815# VSUBS 0.216482f
C8770 XM4/a_100_n51682# VSUBS 0.190616f
C8771 XM4/a_n100_n51779# VSUBS 0.216482f
C8772 XM4/a_100_n50646# VSUBS 0.190616f
C8773 XM4/a_n100_n50743# VSUBS 0.216482f
C8774 XM4/a_100_n49610# VSUBS 0.190616f
C8775 XM4/a_n100_n49707# VSUBS 0.216482f
C8776 XM4/a_100_n48574# VSUBS 0.190616f
C8777 XM4/a_n100_n48671# VSUBS 0.216482f
C8778 XM4/a_100_n47538# VSUBS 0.190616f
C8779 XM4/a_n100_n47635# VSUBS 0.216482f
C8780 XM4/a_100_n46502# VSUBS 0.190616f
C8781 XM4/a_n100_n46599# VSUBS 0.216482f
C8782 XM4/a_100_n45466# VSUBS 0.190616f
C8783 XM4/a_n100_n45563# VSUBS 0.216482f
C8784 XM4/a_100_n44430# VSUBS 0.190616f
C8785 XM4/a_n100_n44527# VSUBS 0.216482f
C8786 XM4/a_100_n43394# VSUBS 0.190616f
C8787 XM4/a_n100_n43491# VSUBS 0.216482f
C8788 XM4/a_100_n42358# VSUBS 0.190616f
C8789 XM4/a_n100_n42455# VSUBS 0.216482f
C8790 XM4/a_100_n41322# VSUBS 0.190616f
C8791 XM4/a_n100_n41419# VSUBS 0.216482f
C8792 XM4/a_100_n40286# VSUBS 0.190616f
C8793 XM4/a_n100_n40383# VSUBS 0.216482f
C8794 XM4/a_100_n39250# VSUBS 0.190616f
C8795 XM4/a_n100_n39347# VSUBS 0.216482f
C8796 XM4/a_100_n38214# VSUBS 0.190616f
C8797 XM4/a_n100_n38311# VSUBS 0.216482f
C8798 XM4/a_100_n37178# VSUBS 0.190616f
C8799 XM4/a_n100_n37275# VSUBS 0.216482f
C8800 XM4/a_100_n36142# VSUBS 0.190616f
C8801 XM4/a_n100_n36239# VSUBS 0.216482f
C8802 XM4/a_100_n35106# VSUBS 0.190616f
C8803 XM4/a_n100_n35203# VSUBS 0.216482f
C8804 XM4/a_100_n34070# VSUBS 0.190616f
C8805 XM4/a_n100_n34167# VSUBS 0.216482f
C8806 XM4/a_100_n33034# VSUBS 0.190616f
C8807 XM4/a_n100_n33131# VSUBS 0.216482f
C8808 XM4/a_100_n31998# VSUBS 0.190616f
C8809 XM4/a_n100_n32095# VSUBS 0.216482f
C8810 XM4/a_100_n30962# VSUBS 0.190616f
C8811 XM4/a_n100_n31059# VSUBS 0.216482f
C8812 XM4/a_100_n29926# VSUBS 0.190616f
C8813 XM4/a_n100_n30023# VSUBS 0.216482f
C8814 XM4/a_100_n28890# VSUBS 0.190616f
C8815 XM4/a_n100_n28987# VSUBS 0.216482f
C8816 XM4/a_100_n27854# VSUBS 0.190616f
C8817 XM4/a_n100_n27951# VSUBS 0.216482f
C8818 XM4/a_100_n26818# VSUBS 0.190616f
C8819 XM4/a_n100_n26915# VSUBS 0.216482f
C8820 XM4/a_100_n25782# VSUBS 0.190616f
C8821 XM4/a_n100_n25879# VSUBS 0.216482f
C8822 XM4/a_100_n24746# VSUBS 0.190616f
C8823 XM4/a_n100_n24843# VSUBS 0.216482f
C8824 XM4/a_100_n23710# VSUBS 0.190616f
C8825 XM4/a_n100_n23807# VSUBS 0.216482f
C8826 XM4/a_100_n22674# VSUBS 0.190616f
C8827 XM4/a_n100_n22771# VSUBS 0.216482f
C8828 XM4/a_100_n21638# VSUBS 0.190616f
C8829 XM4/a_n100_n21735# VSUBS 0.216482f
C8830 XM4/a_100_n20602# VSUBS 0.190616f
C8831 XM4/a_n100_n20699# VSUBS 0.216482f
C8832 XM4/a_100_n19566# VSUBS 0.190616f
C8833 XM4/a_n100_n19663# VSUBS 0.216482f
C8834 XM4/a_100_n18530# VSUBS 0.190616f
C8835 XM4/a_n100_n18627# VSUBS 0.216482f
C8836 XM4/a_100_n17494# VSUBS 0.190616f
C8837 XM4/a_n100_n17591# VSUBS 0.216482f
C8838 XM4/a_100_n16458# VSUBS 0.190616f
C8839 XM4/a_n100_n16555# VSUBS 0.216482f
C8840 XM4/a_100_n15422# VSUBS 0.190616f
C8841 XM4/a_n100_n15519# VSUBS 0.216482f
C8842 XM4/a_100_n14386# VSUBS 0.190616f
C8843 XM4/a_n100_n14483# VSUBS 0.216482f
C8844 XM4/a_100_n13350# VSUBS 0.190616f
C8845 XM4/a_n100_n13447# VSUBS 0.216482f
C8846 XM4/a_100_n12314# VSUBS 0.190616f
C8847 XM4/a_n100_n12411# VSUBS 0.216482f
C8848 XM4/a_100_n11278# VSUBS 0.190616f
C8849 XM4/a_n100_n11375# VSUBS 0.216482f
C8850 XM4/a_100_n10242# VSUBS 0.190616f
C8851 XM4/a_n100_n10339# VSUBS 0.216482f
C8852 XM4/a_100_n9206# VSUBS 0.190616f
C8853 XM4/a_n100_n9303# VSUBS 0.216482f
C8854 XM4/a_100_n8170# VSUBS 0.190616f
C8855 XM4/a_n100_n8267# VSUBS 0.216482f
C8856 XM4/a_100_n7134# VSUBS 0.190616f
C8857 XM4/a_n100_n7231# VSUBS 0.216482f
C8858 XM4/a_100_n6098# VSUBS 0.190616f
C8859 XM4/a_n100_n6195# VSUBS 0.216482f
C8860 XM4/a_100_n5062# VSUBS 0.190616f
C8861 XM4/a_n100_n5159# VSUBS 0.216482f
C8862 XM4/a_100_n4026# VSUBS 0.190616f
C8863 XM4/a_n100_n4123# VSUBS 0.216482f
C8864 XM4/a_100_n2990# VSUBS 0.190616f
C8865 XM4/a_n100_n3087# VSUBS 0.216482f
C8866 XM4/a_100_n1954# VSUBS 0.190616f
C8867 XM4/a_n100_n2051# VSUBS 0.216482f
C8868 XM4/a_100_n918# VSUBS 0.190616f
C8869 XM4/a_n100_n1015# VSUBS 0.216482f
C8870 XM4/a_100_118# VSUBS 0.190616f
C8871 XM4/a_n100_21# VSUBS 0.216482f
C8872 XM4/a_100_1154# VSUBS 0.190616f
C8873 XM4/a_n100_1057# VSUBS 0.216482f
C8874 XM4/a_100_2190# VSUBS 0.190616f
C8875 XM4/a_n100_2093# VSUBS 0.216482f
C8876 XM4/a_100_3226# VSUBS 0.190616f
C8877 XM4/a_n100_3129# VSUBS 0.216482f
C8878 XM4/a_100_4262# VSUBS 0.190616f
C8879 XM4/a_n100_4165# VSUBS 0.216482f
C8880 XM4/a_100_5298# VSUBS 0.190616f
C8881 XM4/a_n100_5201# VSUBS 0.216482f
C8882 XM4/a_100_6334# VSUBS 0.190616f
C8883 XM4/a_n100_6237# VSUBS 0.216482f
C8884 XM4/a_100_7370# VSUBS 0.190616f
C8885 XM4/a_n100_7273# VSUBS 0.216482f
C8886 XM4/a_100_8406# VSUBS 0.190616f
C8887 XM4/a_n100_8309# VSUBS 0.216482f
C8888 XM4/a_100_9442# VSUBS 0.190616f
C8889 XM4/a_n100_9345# VSUBS 0.216482f
C8890 XM4/a_100_10478# VSUBS 0.190616f
C8891 XM4/a_n100_10381# VSUBS 0.216482f
C8892 XM4/a_100_11514# VSUBS 0.190616f
C8893 XM4/a_n100_11417# VSUBS 0.216482f
C8894 XM4/a_100_12550# VSUBS 0.190616f
C8895 XM4/a_n100_12453# VSUBS 0.216482f
C8896 XM4/a_100_13586# VSUBS 0.190616f
C8897 XM4/a_n100_13489# VSUBS 0.216482f
C8898 XM4/a_100_14622# VSUBS 0.190616f
C8899 XM4/a_n100_14525# VSUBS 0.216482f
C8900 XM4/a_100_15658# VSUBS 0.190616f
C8901 XM4/a_n100_15561# VSUBS 0.216482f
C8902 XM4/a_100_16694# VSUBS 0.190616f
C8903 XM4/a_n100_16597# VSUBS 0.216482f
C8904 XM4/a_100_17730# VSUBS 0.190616f
C8905 XM4/a_n100_17633# VSUBS 0.216482f
C8906 XM4/a_100_18766# VSUBS 0.190616f
C8907 XM4/a_n100_18669# VSUBS 0.216482f
C8908 XM4/a_100_19802# VSUBS 0.190616f
C8909 XM4/a_n100_19705# VSUBS 0.216482f
C8910 XM4/a_100_20838# VSUBS 0.190616f
C8911 XM4/a_n100_20741# VSUBS 0.216482f
C8912 XM4/a_100_21874# VSUBS 0.190616f
C8913 XM4/a_n100_21777# VSUBS 0.216482f
C8914 XM4/a_100_22910# VSUBS 0.190616f
C8915 XM4/a_n100_22813# VSUBS 0.216482f
C8916 XM4/a_100_23946# VSUBS 0.190616f
C8917 XM4/a_n100_23849# VSUBS 0.216482f
C8918 XM4/a_100_24982# VSUBS 0.190616f
C8919 XM4/a_n100_24885# VSUBS 0.216482f
C8920 XM4/a_100_26018# VSUBS 0.190616f
C8921 XM4/a_n100_25921# VSUBS 0.216482f
C8922 XM4/a_100_27054# VSUBS 0.190616f
C8923 XM4/a_n100_26957# VSUBS 0.216482f
C8924 XM4/a_100_28090# VSUBS 0.190616f
C8925 XM4/a_n100_27993# VSUBS 0.216482f
C8926 XM4/a_100_29126# VSUBS 0.190616f
C8927 XM4/a_n100_29029# VSUBS 0.216482f
C8928 XM4/a_100_30162# VSUBS 0.190616f
C8929 XM4/a_n100_30065# VSUBS 0.216482f
C8930 XM4/a_100_31198# VSUBS 0.190616f
C8931 XM4/a_n100_31101# VSUBS 0.216482f
C8932 XM4/a_100_32234# VSUBS 0.190616f
C8933 XM4/a_n100_32137# VSUBS 0.216482f
C8934 XM4/a_100_33270# VSUBS 0.190616f
C8935 XM4/a_n100_33173# VSUBS 0.216482f
C8936 XM4/a_100_34306# VSUBS 0.190616f
C8937 XM4/a_n100_34209# VSUBS 0.216482f
C8938 XM4/a_100_35342# VSUBS 0.190616f
C8939 XM4/a_n100_35245# VSUBS 0.216482f
C8940 XM4/a_100_36378# VSUBS 0.190616f
C8941 XM4/a_n100_36281# VSUBS 0.216482f
C8942 XM4/a_100_37414# VSUBS 0.190616f
C8943 XM4/a_n100_37317# VSUBS 0.216482f
C8944 XM4/a_100_38450# VSUBS 0.190616f
C8945 XM4/a_n100_38353# VSUBS 0.216482f
C8946 XM4/a_100_39486# VSUBS 0.190616f
C8947 XM4/a_n100_39389# VSUBS 0.216482f
C8948 XM4/a_100_40522# VSUBS 0.190616f
C8949 XM4/a_n100_40425# VSUBS 0.216482f
C8950 XM4/a_100_41558# VSUBS 0.190616f
C8951 XM4/a_n100_41461# VSUBS 0.216482f
C8952 XM4/a_100_42594# VSUBS 0.190616f
C8953 XM4/a_n100_42497# VSUBS 0.216482f
C8954 XM4/a_100_43630# VSUBS 0.190616f
C8955 XM4/a_n100_43533# VSUBS 0.216482f
C8956 XM4/a_100_44666# VSUBS 0.190616f
C8957 XM4/a_n100_44569# VSUBS 0.216482f
C8958 XM4/a_100_45702# VSUBS 0.190616f
C8959 XM4/a_n100_45605# VSUBS 0.216482f
C8960 XM4/a_100_46738# VSUBS 0.190616f
C8961 XM4/a_n100_46641# VSUBS 0.216482f
C8962 XM4/a_100_47774# VSUBS 0.190616f
C8963 XM4/a_n100_47677# VSUBS 0.216482f
C8964 XM4/a_100_48810# VSUBS 0.190616f
C8965 XM4/a_n100_48713# VSUBS 0.216482f
C8966 XM4/a_100_49846# VSUBS 0.190616f
C8967 XM4/a_n100_49749# VSUBS 0.216482f
C8968 XM4/a_100_50882# VSUBS 0.190616f
C8969 XM4/a_n100_50785# VSUBS 0.216482f
C8970 XM4/a_100_51918# VSUBS 0.190616f
C8971 XM4/a_n100_51821# VSUBS 0.216482f
C8972 XM4/a_100_52954# VSUBS 0.190616f
C8973 XM4/a_n100_52857# VSUBS 0.216482f
C8974 XM4/a_100_53990# VSUBS 0.190616f
C8975 XM4/a_n100_53893# VSUBS 0.216482f
C8976 XM4/a_100_55026# VSUBS 0.190616f
C8977 XM4/a_n100_54929# VSUBS 0.216482f
C8978 XM4/a_100_56062# VSUBS 0.190616f
C8979 XM4/a_n100_55965# VSUBS 0.216482f
C8980 XM4/a_100_57098# VSUBS 0.190616f
C8981 XM4/a_n100_57001# VSUBS 0.216482f
C8982 XM4/a_100_58134# VSUBS 0.190616f
C8983 XM4/a_n100_58037# VSUBS 0.216482f
C8984 XM4/a_100_59170# VSUBS 0.190616f
C8985 XM4/a_n100_59073# VSUBS 0.216482f
C8986 XM4/a_100_60206# VSUBS 0.190616f
C8987 XM4/a_n100_60109# VSUBS 0.216482f
C8988 XM4/a_100_61242# VSUBS 0.190616f
C8989 XM4/a_n100_61145# VSUBS 0.216482f
C8990 XM4/a_100_62278# VSUBS 0.190616f
C8991 XM4/a_n100_62181# VSUBS 0.216482f
C8992 XM4/a_100_63314# VSUBS 0.190616f
C8993 XM4/a_n100_63217# VSUBS 0.216482f
C8994 XM4/a_100_64350# VSUBS 0.190616f
C8995 XM4/a_n100_64253# VSUBS 0.216482f
C8996 XM4/a_100_65386# VSUBS 0.190616f
C8997 XM4/a_n100_65289# VSUBS 0.216482f
C8998 XM4/a_100_66422# VSUBS 0.190616f
C8999 XM4/a_n100_66325# VSUBS 0.216482f
C9000 XM4/a_100_67458# VSUBS 0.190616f
C9001 XM4/a_n100_67361# VSUBS 0.216482f
C9002 XM4/a_100_68494# VSUBS 0.190616f
C9003 XM4/a_n100_68397# VSUBS 0.216482f
C9004 XM4/a_100_69530# VSUBS 0.190616f
C9005 XM4/a_n100_69433# VSUBS 0.216482f
C9006 XM4/a_100_70566# VSUBS 0.190616f
C9007 XM4/a_n100_70469# VSUBS 0.216482f
C9008 XM4/a_100_71602# VSUBS 0.190616f
C9009 XM4/a_n100_71505# VSUBS 0.216482f
C9010 XM4/a_100_72638# VSUBS 0.190616f
C9011 XM4/a_n100_72541# VSUBS 0.216482f
C9012 XM4/a_100_73674# VSUBS 0.190616f
C9013 XM4/a_n100_73577# VSUBS 0.216482f
C9014 XM4/a_100_74710# VSUBS 0.190616f
C9015 XM4/a_n100_74613# VSUBS 0.216482f
C9016 XM4/a_100_75746# VSUBS 0.190616f
C9017 XM4/a_n100_75649# VSUBS 0.216482f
C9018 XM4/a_100_76782# VSUBS 0.190616f
C9019 XM4/a_n100_76685# VSUBS 0.216482f
C9020 XM4/a_100_77818# VSUBS 0.190616f
C9021 XM4/a_n100_77721# VSUBS 0.216482f
C9022 XM4/a_100_78854# VSUBS 0.190616f
C9023 XM4/a_n100_78757# VSUBS 0.216482f
C9024 XM4/a_100_79890# VSUBS 0.190616f
C9025 XM4/a_n100_79793# VSUBS 0.216482f
C9026 XM4/a_100_80926# VSUBS 0.190616f
C9027 XM4/a_n100_80829# VSUBS 0.216482f
C9028 XM4/a_100_81962# VSUBS 0.190616f
C9029 XM4/a_n100_81865# VSUBS 0.216482f
C9030 XM4/a_100_82998# VSUBS 0.190616f
C9031 XM4/a_n100_82901# VSUBS 0.216482f
C9032 XM4/a_100_84034# VSUBS 0.190616f
C9033 XM4/a_n100_83937# VSUBS 0.216482f
C9034 XM4/a_100_85070# VSUBS 0.190616f
C9035 XM4/a_n100_84973# VSUBS 0.216482f
C9036 XM4/a_100_86106# VSUBS 0.190616f
C9037 XM4/a_n100_86009# VSUBS 0.216482f
C9038 XM4/a_100_87142# VSUBS 0.190616f
C9039 XM4/a_n100_87045# VSUBS 0.216482f
C9040 XM4/a_100_88178# VSUBS 0.190616f
C9041 XM4/a_n100_88081# VSUBS 0.216482f
C9042 XM4/a_100_89214# VSUBS 0.190616f
C9043 XM4/a_n100_89117# VSUBS 0.216482f
C9044 XM4/a_100_90250# VSUBS 0.190616f
C9045 XM4/a_n100_90153# VSUBS 0.216482f
C9046 XM4/a_100_91286# VSUBS 0.190616f
C9047 XM4/a_n100_91189# VSUBS 0.216482f
C9048 XM4/a_100_92322# VSUBS 0.190616f
C9049 XM4/a_n100_92225# VSUBS 0.216482f
C9050 XM4/a_100_93358# VSUBS 0.190616f
C9051 XM4/a_n100_93261# VSUBS 0.216482f
C9052 XM4/a_100_94394# VSUBS 0.190616f
C9053 XM4/a_n100_94297# VSUBS 0.216482f
C9054 XM4/a_100_95430# VSUBS 0.190616f
C9055 XM4/a_n100_95333# VSUBS 0.216482f
C9056 XM4/a_100_96466# VSUBS 0.190616f
C9057 XM4/a_n100_96369# VSUBS 0.216482f
C9058 XM4/a_100_97502# VSUBS 0.190616f
C9059 XM4/a_n100_97405# VSUBS 0.216482f
C9060 XM4/a_100_98538# VSUBS 0.190616f
C9061 XM4/a_n100_98441# VSUBS 0.216482f
C9062 XM4/a_100_99574# VSUBS 0.190616f
C9063 XM4/a_n100_99477# VSUBS 0.216482f
C9064 XM4/a_100_100610# VSUBS 0.190616f
C9065 XM4/a_n100_100513# VSUBS 0.216482f
C9066 XM4/a_100_101646# VSUBS 0.190616f
C9067 XM4/a_n100_101549# VSUBS 0.216482f
C9068 XM4/a_100_102682# VSUBS 0.190616f
C9069 XM4/a_n100_102585# VSUBS 0.216482f
C9070 XM4/a_100_103718# VSUBS 0.190616f
C9071 XM4/a_n100_103621# VSUBS 0.216482f
C9072 XM4/a_100_104754# VSUBS 0.190616f
C9073 XM4/a_n100_104657# VSUBS 0.216482f
C9074 XM4/a_100_105790# VSUBS 0.190616f
C9075 XM4/a_n100_105693# VSUBS 0.216482f
C9076 XM4/a_100_106826# VSUBS 0.190616f
C9077 XM4/a_n100_106729# VSUBS 0.216482f
C9078 XM4/a_100_107862# VSUBS 0.190616f
C9079 XM4/a_n100_107765# VSUBS 0.216482f
C9080 XM4/a_100_108898# VSUBS 0.190616f
C9081 XM4/a_n100_108801# VSUBS 0.216482f
C9082 XM4/a_100_109934# VSUBS 0.190616f
C9083 XM4/a_n100_109837# VSUBS 0.216482f
C9084 XM4/a_100_110970# VSUBS 0.190616f
C9085 XM4/a_n100_110873# VSUBS 0.216482f
C9086 XM4/a_100_112006# VSUBS 0.190616f
C9087 XM4/a_n100_111909# VSUBS 0.216482f
C9088 XM4/a_100_113042# VSUBS 0.190616f
C9089 XM4/a_n100_112945# VSUBS 0.216482f
C9090 XM4/a_100_114078# VSUBS 0.190616f
C9091 XM4/a_n100_113981# VSUBS 0.216482f
C9092 XM4/a_100_115114# VSUBS 0.190616f
C9093 XM4/a_n100_115017# VSUBS 0.216482f
C9094 XM4/a_100_116150# VSUBS 0.190616f
C9095 XM4/a_n100_116053# VSUBS 0.216482f
C9096 XM4/a_100_117186# VSUBS 0.190616f
C9097 XM4/a_n100_117089# VSUBS 0.216482f
C9098 XM4/a_100_118222# VSUBS 0.190616f
C9099 XM4/a_n100_118125# VSUBS 0.216482f
C9100 XM4/a_100_119258# VSUBS 0.190616f
C9101 XM4/a_n100_119161# VSUBS 0.216482f
C9102 XM4/a_100_120294# VSUBS 0.190616f
C9103 XM4/a_n100_120197# VSUBS 0.216482f
C9104 XM4/a_100_121330# VSUBS 0.190616f
C9105 XM4/a_n100_121233# VSUBS 0.216482f
C9106 XM4/a_100_122366# VSUBS 0.190616f
C9107 XM4/a_n100_122269# VSUBS 0.216482f
C9108 XM4/a_100_123402# VSUBS 0.190616f
C9109 XM4/a_n100_123305# VSUBS 0.216482f
C9110 XM4/a_100_124438# VSUBS 0.190616f
C9111 XM4/a_n100_124341# VSUBS 0.216482f
C9112 XM4/a_100_125474# VSUBS 0.190616f
C9113 XM4/a_n100_125377# VSUBS 0.216482f
C9114 XM4/a_100_126510# VSUBS 0.190616f
C9115 XM4/a_n100_126413# VSUBS 0.216482f
C9116 XM4/a_100_127546# VSUBS 0.190616f
C9117 XM4/a_n100_127449# VSUBS 0.216482f
C9118 XM4/a_100_128582# VSUBS 0.190616f
C9119 XM4/a_n100_128485# VSUBS 0.216482f
C9120 XM4/a_100_129618# VSUBS 0.190616f
C9121 XM4/a_n100_129521# VSUBS 0.216482f
C9122 XM4/a_100_130654# VSUBS 0.190616f
C9123 XM4/a_n100_130557# VSUBS 0.216482f
C9124 XM4/a_100_131690# VSUBS 0.196066f
C9125 XM4/a_n100_131593# VSUBS 0.260213f
C9126 XM3/a_n158_n132490# VSUBS 0.196066f
C9127 XM3/a_n100_n132587# VSUBS 0.260213f
C9128 XM3/a_n158_n131454# VSUBS 0.190616f
C9129 XM3/a_n100_n131551# VSUBS 0.216482f
C9130 XM3/a_n158_n130418# VSUBS 0.190616f
C9131 XM3/a_n100_n130515# VSUBS 0.216482f
C9132 XM3/a_n158_n129382# VSUBS 0.190616f
C9133 XM3/a_n100_n129479# VSUBS 0.216482f
C9134 XM3/a_n158_n128346# VSUBS 0.190616f
C9135 XM3/a_n100_n128443# VSUBS 0.216482f
C9136 XM3/a_n158_n127310# VSUBS 0.190616f
C9137 XM3/a_n100_n127407# VSUBS 0.216482f
C9138 XM3/a_n158_n126274# VSUBS 0.190616f
C9139 XM3/a_n100_n126371# VSUBS 0.216482f
C9140 XM3/a_n158_n125238# VSUBS 0.190616f
C9141 XM3/a_n100_n125335# VSUBS 0.216482f
C9142 XM3/a_n158_n124202# VSUBS 0.190616f
C9143 XM3/a_n100_n124299# VSUBS 0.216482f
C9144 XM3/a_n158_n123166# VSUBS 0.190616f
C9145 XM3/a_n100_n123263# VSUBS 0.216482f
C9146 XM3/a_n158_n122130# VSUBS 0.190616f
C9147 XM3/a_n100_n122227# VSUBS 0.216482f
C9148 XM3/a_n158_n121094# VSUBS 0.190616f
C9149 XM3/a_n100_n121191# VSUBS 0.216482f
C9150 XM3/a_n158_n120058# VSUBS 0.190616f
C9151 XM3/a_n100_n120155# VSUBS 0.216482f
C9152 XM3/a_n158_n119022# VSUBS 0.190616f
C9153 XM3/a_n100_n119119# VSUBS 0.216482f
C9154 XM3/a_n158_n117986# VSUBS 0.190616f
C9155 XM3/a_n100_n118083# VSUBS 0.216482f
C9156 XM3/a_n158_n116950# VSUBS 0.190616f
C9157 XM3/a_n100_n117047# VSUBS 0.216482f
C9158 XM3/a_n158_n115914# VSUBS 0.190616f
C9159 XM3/a_n100_n116011# VSUBS 0.216482f
C9160 XM3/a_n158_n114878# VSUBS 0.190616f
C9161 XM3/a_n100_n114975# VSUBS 0.216482f
C9162 XM3/a_n158_n113842# VSUBS 0.190616f
C9163 XM3/a_n100_n113939# VSUBS 0.216482f
C9164 XM3/a_n158_n112806# VSUBS 0.190616f
C9165 XM3/a_n100_n112903# VSUBS 0.216482f
C9166 XM3/a_n158_n111770# VSUBS 0.190616f
C9167 XM3/a_n100_n111867# VSUBS 0.216482f
C9168 XM3/a_n158_n110734# VSUBS 0.190616f
C9169 XM3/a_n100_n110831# VSUBS 0.216482f
C9170 XM3/a_n158_n109698# VSUBS 0.190616f
C9171 XM3/a_n100_n109795# VSUBS 0.216482f
C9172 XM3/a_n158_n108662# VSUBS 0.190616f
C9173 XM3/a_n100_n108759# VSUBS 0.216482f
C9174 XM3/a_n158_n107626# VSUBS 0.190616f
C9175 XM3/a_n100_n107723# VSUBS 0.216482f
C9176 XM3/a_n158_n106590# VSUBS 0.190616f
C9177 XM3/a_n100_n106687# VSUBS 0.216482f
C9178 XM3/a_n158_n105554# VSUBS 0.190616f
C9179 XM3/a_n100_n105651# VSUBS 0.216482f
C9180 XM3/a_n158_n104518# VSUBS 0.190616f
C9181 XM3/a_n100_n104615# VSUBS 0.216482f
C9182 XM3/a_n158_n103482# VSUBS 0.190616f
C9183 XM3/a_n100_n103579# VSUBS 0.216482f
C9184 XM3/a_n158_n102446# VSUBS 0.190616f
C9185 XM3/a_n100_n102543# VSUBS 0.216482f
C9186 XM3/a_n158_n101410# VSUBS 0.190616f
C9187 XM3/a_n100_n101507# VSUBS 0.216482f
C9188 XM3/a_n158_n100374# VSUBS 0.190616f
C9189 XM3/a_n100_n100471# VSUBS 0.216482f
C9190 XM3/a_n158_n99338# VSUBS 0.190616f
C9191 XM3/a_n100_n99435# VSUBS 0.216482f
C9192 XM3/a_n158_n98302# VSUBS 0.190616f
C9193 XM3/a_n100_n98399# VSUBS 0.216482f
C9194 XM3/a_n158_n97266# VSUBS 0.190616f
C9195 XM3/a_n100_n97363# VSUBS 0.216482f
C9196 XM3/a_n158_n96230# VSUBS 0.190616f
C9197 XM3/a_n100_n96327# VSUBS 0.216482f
C9198 XM3/a_n158_n95194# VSUBS 0.190616f
C9199 XM3/a_n100_n95291# VSUBS 0.216482f
C9200 XM3/a_n158_n94158# VSUBS 0.190616f
C9201 XM3/a_n100_n94255# VSUBS 0.216482f
C9202 XM3/a_n158_n93122# VSUBS 0.190616f
C9203 XM3/a_n100_n93219# VSUBS 0.216482f
C9204 XM3/a_n158_n92086# VSUBS 0.190616f
C9205 XM3/a_n100_n92183# VSUBS 0.216482f
C9206 XM3/a_n158_n91050# VSUBS 0.190616f
C9207 XM3/a_n100_n91147# VSUBS 0.216482f
C9208 XM3/a_n158_n90014# VSUBS 0.190616f
C9209 XM3/a_n100_n90111# VSUBS 0.216482f
C9210 XM3/a_n158_n88978# VSUBS 0.190616f
C9211 XM3/a_n100_n89075# VSUBS 0.216482f
C9212 XM3/a_n158_n87942# VSUBS 0.190616f
C9213 XM3/a_n100_n88039# VSUBS 0.216482f
C9214 XM3/a_n158_n86906# VSUBS 0.190616f
C9215 XM3/a_n100_n87003# VSUBS 0.216482f
C9216 XM3/a_n158_n85870# VSUBS 0.190616f
C9217 XM3/a_n100_n85967# VSUBS 0.216482f
C9218 XM3/a_n158_n84834# VSUBS 0.190616f
C9219 XM3/a_n100_n84931# VSUBS 0.216482f
C9220 XM3/a_n158_n83798# VSUBS 0.190616f
C9221 XM3/a_n100_n83895# VSUBS 0.216482f
C9222 XM3/a_n158_n82762# VSUBS 0.190616f
C9223 XM3/a_n100_n82859# VSUBS 0.216482f
C9224 XM3/a_n158_n81726# VSUBS 0.190616f
C9225 XM3/a_n100_n81823# VSUBS 0.216482f
C9226 XM3/a_n158_n80690# VSUBS 0.190616f
C9227 XM3/a_n100_n80787# VSUBS 0.216482f
C9228 XM3/a_n158_n79654# VSUBS 0.190616f
C9229 XM3/a_n100_n79751# VSUBS 0.216482f
C9230 XM3/a_n158_n78618# VSUBS 0.190616f
C9231 XM3/a_n100_n78715# VSUBS 0.216482f
C9232 XM3/a_n158_n77582# VSUBS 0.190616f
C9233 XM3/a_n100_n77679# VSUBS 0.216482f
C9234 XM3/a_n158_n76546# VSUBS 0.190616f
C9235 XM3/a_n100_n76643# VSUBS 0.216482f
C9236 XM3/a_n158_n75510# VSUBS 0.190616f
C9237 XM3/a_n100_n75607# VSUBS 0.216482f
C9238 XM3/a_n158_n74474# VSUBS 0.190616f
C9239 XM3/a_n100_n74571# VSUBS 0.216482f
C9240 XM3/a_n158_n73438# VSUBS 0.190616f
C9241 XM3/a_n100_n73535# VSUBS 0.216482f
C9242 XM3/a_n158_n72402# VSUBS 0.190616f
C9243 XM3/a_n100_n72499# VSUBS 0.216482f
C9244 XM3/a_n158_n71366# VSUBS 0.190616f
C9245 XM3/a_n100_n71463# VSUBS 0.216482f
C9246 XM3/a_n158_n70330# VSUBS 0.190616f
C9247 XM3/a_n100_n70427# VSUBS 0.216482f
C9248 XM3/a_n158_n69294# VSUBS 0.190616f
C9249 XM3/a_n100_n69391# VSUBS 0.216482f
C9250 XM3/a_n158_n68258# VSUBS 0.190616f
C9251 XM3/a_n100_n68355# VSUBS 0.216482f
C9252 XM3/a_n158_n67222# VSUBS 0.190616f
C9253 XM3/a_n100_n67319# VSUBS 0.216482f
C9254 XM3/a_n158_n66186# VSUBS 0.190616f
C9255 XM3/a_n100_n66283# VSUBS 0.216482f
C9256 XM3/a_n158_n65150# VSUBS 0.190616f
C9257 XM3/a_n100_n65247# VSUBS 0.216482f
C9258 XM3/a_n158_n64114# VSUBS 0.190616f
C9259 XM3/a_n100_n64211# VSUBS 0.216482f
C9260 XM3/a_n158_n63078# VSUBS 0.190616f
C9261 XM3/a_n100_n63175# VSUBS 0.216482f
C9262 XM3/a_n158_n62042# VSUBS 0.190616f
C9263 XM3/a_n100_n62139# VSUBS 0.216482f
C9264 XM3/a_n158_n61006# VSUBS 0.190616f
C9265 XM3/a_n100_n61103# VSUBS 0.216482f
C9266 XM3/a_n158_n59970# VSUBS 0.190616f
C9267 XM3/a_n100_n60067# VSUBS 0.216482f
C9268 XM3/a_n158_n58934# VSUBS 0.190616f
C9269 XM3/a_n100_n59031# VSUBS 0.216482f
C9270 XM3/a_n158_n57898# VSUBS 0.190616f
C9271 XM3/a_n100_n57995# VSUBS 0.216482f
C9272 XM3/a_n158_n56862# VSUBS 0.190616f
C9273 XM3/a_n100_n56959# VSUBS 0.216482f
C9274 XM3/a_n158_n55826# VSUBS 0.190616f
C9275 XM3/a_n100_n55923# VSUBS 0.216482f
C9276 XM3/a_n158_n54790# VSUBS 0.190616f
C9277 XM3/a_n100_n54887# VSUBS 0.216482f
C9278 XM3/a_n158_n53754# VSUBS 0.190616f
C9279 XM3/a_n100_n53851# VSUBS 0.216482f
C9280 XM3/a_n158_n52718# VSUBS 0.190616f
C9281 XM3/a_n100_n52815# VSUBS 0.216482f
C9282 XM3/a_n158_n51682# VSUBS 0.190616f
C9283 XM3/a_n100_n51779# VSUBS 0.216482f
C9284 XM3/a_n158_n50646# VSUBS 0.190616f
C9285 XM3/a_n100_n50743# VSUBS 0.216482f
C9286 XM3/a_n158_n49610# VSUBS 0.190616f
C9287 XM3/a_n100_n49707# VSUBS 0.216482f
C9288 XM3/a_n158_n48574# VSUBS 0.190616f
C9289 XM3/a_n100_n48671# VSUBS 0.216482f
C9290 XM3/a_n158_n47538# VSUBS 0.190616f
C9291 XM3/a_n100_n47635# VSUBS 0.216482f
C9292 XM3/a_n158_n46502# VSUBS 0.190616f
C9293 XM3/a_n100_n46599# VSUBS 0.216482f
C9294 XM3/a_n158_n45466# VSUBS 0.190616f
C9295 XM3/a_n100_n45563# VSUBS 0.216482f
C9296 XM3/a_n158_n44430# VSUBS 0.190616f
C9297 XM3/a_n100_n44527# VSUBS 0.216482f
C9298 XM3/a_n158_n43394# VSUBS 0.190616f
C9299 XM3/a_n100_n43491# VSUBS 0.216482f
C9300 XM3/a_n158_n42358# VSUBS 0.190616f
C9301 XM3/a_n100_n42455# VSUBS 0.216482f
C9302 XM3/a_n158_n41322# VSUBS 0.190616f
C9303 XM3/a_n100_n41419# VSUBS 0.216482f
C9304 XM3/a_n158_n40286# VSUBS 0.190616f
C9305 XM3/a_n100_n40383# VSUBS 0.216482f
C9306 XM3/a_n158_n39250# VSUBS 0.190616f
C9307 XM3/a_n100_n39347# VSUBS 0.216482f
C9308 XM3/a_n158_n38214# VSUBS 0.190616f
C9309 XM3/a_n100_n38311# VSUBS 0.216482f
C9310 XM3/a_n158_n37178# VSUBS 0.190616f
C9311 XM3/a_n100_n37275# VSUBS 0.216482f
C9312 XM3/a_n158_n36142# VSUBS 0.190616f
C9313 XM3/a_n100_n36239# VSUBS 0.216482f
C9314 XM3/a_n158_n35106# VSUBS 0.190616f
C9315 XM3/a_n100_n35203# VSUBS 0.216482f
C9316 XM3/a_n158_n34070# VSUBS 0.190616f
C9317 XM3/a_n100_n34167# VSUBS 0.216482f
C9318 XM3/a_n158_n33034# VSUBS 0.190616f
C9319 XM3/a_n100_n33131# VSUBS 0.216482f
C9320 XM3/a_n158_n31998# VSUBS 0.190616f
C9321 XM3/a_n100_n32095# VSUBS 0.216482f
C9322 XM3/a_n158_n30962# VSUBS 0.190616f
C9323 XM3/a_n100_n31059# VSUBS 0.216482f
C9324 XM3/a_n158_n29926# VSUBS 0.190616f
C9325 XM3/a_n100_n30023# VSUBS 0.216482f
C9326 XM3/a_n158_n28890# VSUBS 0.190616f
C9327 XM3/a_n100_n28987# VSUBS 0.216482f
C9328 XM3/a_n158_n27854# VSUBS 0.190616f
C9329 XM3/a_n100_n27951# VSUBS 0.216482f
C9330 XM3/a_n158_n26818# VSUBS 0.190616f
C9331 XM3/a_n100_n26915# VSUBS 0.216482f
C9332 XM3/a_n158_n25782# VSUBS 0.190616f
C9333 XM3/a_n100_n25879# VSUBS 0.216482f
C9334 XM3/a_n158_n24746# VSUBS 0.190616f
C9335 XM3/a_n100_n24843# VSUBS 0.216482f
C9336 XM3/a_n158_n23710# VSUBS 0.190616f
C9337 XM3/a_n100_n23807# VSUBS 0.216482f
C9338 XM3/a_n158_n22674# VSUBS 0.190616f
C9339 XM3/a_n100_n22771# VSUBS 0.216482f
C9340 XM3/a_n158_n21638# VSUBS 0.190616f
C9341 XM3/a_n100_n21735# VSUBS 0.216482f
C9342 XM3/a_n158_n20602# VSUBS 0.190616f
C9343 XM3/a_n100_n20699# VSUBS 0.216482f
C9344 XM3/a_n158_n19566# VSUBS 0.190616f
C9345 XM3/a_n100_n19663# VSUBS 0.216482f
C9346 XM3/a_n158_n18530# VSUBS 0.190616f
C9347 XM3/a_n100_n18627# VSUBS 0.216482f
C9348 XM3/a_n158_n17494# VSUBS 0.190616f
C9349 XM3/a_n100_n17591# VSUBS 0.216482f
C9350 XM3/a_n158_n16458# VSUBS 0.190616f
C9351 XM3/a_n100_n16555# VSUBS 0.216482f
C9352 XM3/a_n158_n15422# VSUBS 0.190616f
C9353 XM3/a_n100_n15519# VSUBS 0.216482f
C9354 XM3/a_n158_n14386# VSUBS 0.190616f
C9355 XM3/a_n100_n14483# VSUBS 0.216482f
C9356 XM3/a_n158_n13350# VSUBS 0.190616f
C9357 XM3/a_n100_n13447# VSUBS 0.216482f
C9358 XM3/a_n158_n12314# VSUBS 0.190616f
C9359 XM3/a_n100_n12411# VSUBS 0.216482f
C9360 XM3/a_n158_n11278# VSUBS 0.190616f
C9361 XM3/a_n100_n11375# VSUBS 0.216482f
C9362 XM3/a_n158_n10242# VSUBS 0.190616f
C9363 XM3/a_n100_n10339# VSUBS 0.216482f
C9364 XM3/a_n158_n9206# VSUBS 0.190616f
C9365 XM3/a_n100_n9303# VSUBS 0.216482f
C9366 XM3/a_n158_n8170# VSUBS 0.190616f
C9367 XM3/a_n100_n8267# VSUBS 0.216482f
C9368 XM3/a_n158_n7134# VSUBS 0.190616f
C9369 XM3/a_n100_n7231# VSUBS 0.216482f
C9370 XM3/a_n158_n6098# VSUBS 0.190616f
C9371 XM3/a_n100_n6195# VSUBS 0.216482f
C9372 XM3/a_n158_n5062# VSUBS 0.190616f
C9373 XM3/a_n100_n5159# VSUBS 0.216482f
C9374 XM3/a_n158_n4026# VSUBS 0.190616f
C9375 XM3/a_n100_n4123# VSUBS 0.216482f
C9376 XM3/a_n158_n2990# VSUBS 0.190616f
C9377 XM3/a_n100_n3087# VSUBS 0.216482f
C9378 XM3/a_n158_n1954# VSUBS 0.190616f
C9379 XM3/a_n100_n2051# VSUBS 0.216482f
C9380 XM3/a_n158_n918# VSUBS 0.190616f
C9381 XM3/a_n100_n1015# VSUBS 0.216482f
C9382 XM3/a_n158_118# VSUBS 0.190616f
C9383 XM3/a_n100_21# VSUBS 0.216482f
C9384 XM3/a_n158_1154# VSUBS 0.190616f
C9385 XM3/a_n100_1057# VSUBS 0.216482f
C9386 XM3/a_n158_2190# VSUBS 0.190616f
C9387 XM3/a_n100_2093# VSUBS 0.216482f
C9388 XM3/a_n158_3226# VSUBS 0.190616f
C9389 XM3/a_n100_3129# VSUBS 0.216482f
C9390 XM3/a_n158_4262# VSUBS 0.190616f
C9391 XM3/a_n100_4165# VSUBS 0.216482f
C9392 XM3/a_n158_5298# VSUBS 0.190616f
C9393 XM3/a_n100_5201# VSUBS 0.216482f
C9394 XM3/a_n158_6334# VSUBS 0.190616f
C9395 XM3/a_n100_6237# VSUBS 0.216482f
C9396 XM3/a_n158_7370# VSUBS 0.190616f
C9397 XM3/a_n100_7273# VSUBS 0.216482f
C9398 XM3/a_n158_8406# VSUBS 0.190616f
C9399 XM3/a_n100_8309# VSUBS 0.216482f
C9400 XM3/a_n158_9442# VSUBS 0.190616f
C9401 XM3/a_n100_9345# VSUBS 0.216482f
C9402 XM3/a_n158_10478# VSUBS 0.190616f
C9403 XM3/a_n100_10381# VSUBS 0.216482f
C9404 XM3/a_n158_11514# VSUBS 0.190616f
C9405 XM3/a_n100_11417# VSUBS 0.216482f
C9406 XM3/a_n158_12550# VSUBS 0.190616f
C9407 XM3/a_n100_12453# VSUBS 0.216482f
C9408 XM3/a_n158_13586# VSUBS 0.190616f
C9409 XM3/a_n100_13489# VSUBS 0.216482f
C9410 XM3/a_n158_14622# VSUBS 0.190616f
C9411 XM3/a_n100_14525# VSUBS 0.216482f
C9412 XM3/a_n158_15658# VSUBS 0.190616f
C9413 XM3/a_n100_15561# VSUBS 0.216482f
C9414 XM3/a_n158_16694# VSUBS 0.190616f
C9415 XM3/a_n100_16597# VSUBS 0.216482f
C9416 XM3/a_n158_17730# VSUBS 0.190616f
C9417 XM3/a_n100_17633# VSUBS 0.216482f
C9418 XM3/a_n158_18766# VSUBS 0.190616f
C9419 XM3/a_n100_18669# VSUBS 0.216482f
C9420 XM3/a_n158_19802# VSUBS 0.190616f
C9421 XM3/a_n100_19705# VSUBS 0.216482f
C9422 XM3/a_n158_20838# VSUBS 0.190616f
C9423 XM3/a_n100_20741# VSUBS 0.216482f
C9424 XM3/a_n158_21874# VSUBS 0.190616f
C9425 XM3/a_n100_21777# VSUBS 0.216482f
C9426 XM3/a_n158_22910# VSUBS 0.190616f
C9427 XM3/a_n100_22813# VSUBS 0.216482f
C9428 XM3/a_n158_23946# VSUBS 0.190616f
C9429 XM3/a_n100_23849# VSUBS 0.216482f
C9430 XM3/a_n158_24982# VSUBS 0.190616f
C9431 XM3/a_n100_24885# VSUBS 0.216482f
C9432 XM3/a_n158_26018# VSUBS 0.190616f
C9433 XM3/a_n100_25921# VSUBS 0.216482f
C9434 XM3/a_n158_27054# VSUBS 0.190616f
C9435 XM3/a_n100_26957# VSUBS 0.216482f
C9436 XM3/a_n158_28090# VSUBS 0.190616f
C9437 XM3/a_n100_27993# VSUBS 0.216482f
C9438 XM3/a_n158_29126# VSUBS 0.190616f
C9439 XM3/a_n100_29029# VSUBS 0.216482f
C9440 XM3/a_n158_30162# VSUBS 0.190616f
C9441 XM3/a_n100_30065# VSUBS 0.216482f
C9442 XM3/a_n158_31198# VSUBS 0.190616f
C9443 XM3/a_n100_31101# VSUBS 0.216482f
C9444 XM3/a_n158_32234# VSUBS 0.190616f
C9445 XM3/a_n100_32137# VSUBS 0.216482f
C9446 XM3/a_n158_33270# VSUBS 0.190616f
C9447 XM3/a_n100_33173# VSUBS 0.216482f
C9448 XM3/a_n158_34306# VSUBS 0.190616f
C9449 XM3/a_n100_34209# VSUBS 0.216482f
C9450 XM3/a_n158_35342# VSUBS 0.190616f
C9451 XM3/a_n100_35245# VSUBS 0.216482f
C9452 XM3/a_n158_36378# VSUBS 0.190616f
C9453 XM3/a_n100_36281# VSUBS 0.216482f
C9454 XM3/a_n158_37414# VSUBS 0.190616f
C9455 XM3/a_n100_37317# VSUBS 0.216482f
C9456 XM3/a_n158_38450# VSUBS 0.190616f
C9457 XM3/a_n100_38353# VSUBS 0.216482f
C9458 XM3/a_n158_39486# VSUBS 0.190616f
C9459 XM3/a_n100_39389# VSUBS 0.216482f
C9460 XM3/a_n158_40522# VSUBS 0.190616f
C9461 XM3/a_n100_40425# VSUBS 0.216482f
C9462 XM3/a_n158_41558# VSUBS 0.190616f
C9463 XM3/a_n100_41461# VSUBS 0.216482f
C9464 XM3/a_n158_42594# VSUBS 0.190616f
C9465 XM3/a_n100_42497# VSUBS 0.216482f
C9466 XM3/a_n158_43630# VSUBS 0.190616f
C9467 XM3/a_n100_43533# VSUBS 0.216482f
C9468 XM3/a_n158_44666# VSUBS 0.190616f
C9469 XM3/a_n100_44569# VSUBS 0.216482f
C9470 XM3/a_n158_45702# VSUBS 0.190616f
C9471 XM3/a_n100_45605# VSUBS 0.216482f
C9472 XM3/a_n158_46738# VSUBS 0.190616f
C9473 XM3/a_n100_46641# VSUBS 0.216482f
C9474 XM3/a_n158_47774# VSUBS 0.190616f
C9475 XM3/a_n100_47677# VSUBS 0.216482f
C9476 XM3/a_n158_48810# VSUBS 0.190616f
C9477 XM3/a_n100_48713# VSUBS 0.216482f
C9478 XM3/a_n158_49846# VSUBS 0.190616f
C9479 XM3/a_n100_49749# VSUBS 0.216482f
C9480 XM3/a_n158_50882# VSUBS 0.190616f
C9481 XM3/a_n100_50785# VSUBS 0.216482f
C9482 XM3/a_n158_51918# VSUBS 0.190616f
C9483 XM3/a_n100_51821# VSUBS 0.216482f
C9484 XM3/a_n158_52954# VSUBS 0.190616f
C9485 XM3/a_n100_52857# VSUBS 0.216482f
C9486 XM3/a_n158_53990# VSUBS 0.190616f
C9487 XM3/a_n100_53893# VSUBS 0.216482f
C9488 XM3/a_n158_55026# VSUBS 0.190616f
C9489 XM3/a_n100_54929# VSUBS 0.216482f
C9490 XM3/a_n158_56062# VSUBS 0.190616f
C9491 XM3/a_n100_55965# VSUBS 0.216482f
C9492 XM3/a_n158_57098# VSUBS 0.190616f
C9493 XM3/a_n100_57001# VSUBS 0.216482f
C9494 XM3/a_n158_58134# VSUBS 0.190616f
C9495 XM3/a_n100_58037# VSUBS 0.216482f
C9496 XM3/a_n158_59170# VSUBS 0.190616f
C9497 XM3/a_n100_59073# VSUBS 0.216482f
C9498 XM3/a_n158_60206# VSUBS 0.190616f
C9499 XM3/a_n100_60109# VSUBS 0.216482f
C9500 XM3/a_n158_61242# VSUBS 0.190616f
C9501 XM3/a_n100_61145# VSUBS 0.216482f
C9502 XM3/a_n158_62278# VSUBS 0.190616f
C9503 XM3/a_n100_62181# VSUBS 0.216482f
C9504 XM3/a_n158_63314# VSUBS 0.190616f
C9505 XM3/a_n100_63217# VSUBS 0.216482f
C9506 XM3/a_n158_64350# VSUBS 0.190616f
C9507 XM3/a_n100_64253# VSUBS 0.216482f
C9508 XM3/a_n158_65386# VSUBS 0.190616f
C9509 XM3/a_n100_65289# VSUBS 0.216482f
C9510 XM3/a_n158_66422# VSUBS 0.190616f
C9511 XM3/a_n100_66325# VSUBS 0.216482f
C9512 XM3/a_n158_67458# VSUBS 0.190616f
C9513 XM3/a_n100_67361# VSUBS 0.216482f
C9514 XM3/a_n158_68494# VSUBS 0.190616f
C9515 XM3/a_n100_68397# VSUBS 0.216482f
C9516 XM3/a_n158_69530# VSUBS 0.190616f
C9517 XM3/a_n100_69433# VSUBS 0.216482f
C9518 XM3/a_n158_70566# VSUBS 0.190616f
C9519 XM3/a_n100_70469# VSUBS 0.216482f
C9520 XM3/a_n158_71602# VSUBS 0.190616f
C9521 XM3/a_n100_71505# VSUBS 0.216482f
C9522 XM3/a_n158_72638# VSUBS 0.190616f
C9523 XM3/a_n100_72541# VSUBS 0.216482f
C9524 XM3/a_n158_73674# VSUBS 0.190616f
C9525 XM3/a_n100_73577# VSUBS 0.216482f
C9526 XM3/a_n158_74710# VSUBS 0.190616f
C9527 XM3/a_n100_74613# VSUBS 0.216482f
C9528 XM3/a_n158_75746# VSUBS 0.190616f
C9529 XM3/a_n100_75649# VSUBS 0.216482f
C9530 XM3/a_n158_76782# VSUBS 0.190616f
C9531 XM3/a_n100_76685# VSUBS 0.216482f
C9532 XM3/a_n158_77818# VSUBS 0.190616f
C9533 XM3/a_n100_77721# VSUBS 0.216482f
C9534 XM3/a_n158_78854# VSUBS 0.190616f
C9535 XM3/a_n100_78757# VSUBS 0.216482f
C9536 XM3/a_n158_79890# VSUBS 0.190616f
C9537 XM3/a_n100_79793# VSUBS 0.216482f
C9538 XM3/a_n158_80926# VSUBS 0.190616f
C9539 XM3/a_n100_80829# VSUBS 0.216482f
C9540 XM3/a_n158_81962# VSUBS 0.190616f
C9541 XM3/a_n100_81865# VSUBS 0.216482f
C9542 XM3/a_n158_82998# VSUBS 0.190616f
C9543 XM3/a_n100_82901# VSUBS 0.216482f
C9544 XM3/a_n158_84034# VSUBS 0.190616f
C9545 XM3/a_n100_83937# VSUBS 0.216482f
C9546 XM3/a_n158_85070# VSUBS 0.190616f
C9547 XM3/a_n100_84973# VSUBS 0.216482f
C9548 XM3/a_n158_86106# VSUBS 0.190616f
C9549 XM3/a_n100_86009# VSUBS 0.216482f
C9550 XM3/a_n158_87142# VSUBS 0.190616f
C9551 XM3/a_n100_87045# VSUBS 0.216482f
C9552 XM3/a_n158_88178# VSUBS 0.190616f
C9553 XM3/a_n100_88081# VSUBS 0.216482f
C9554 XM3/a_n158_89214# VSUBS 0.190616f
C9555 XM3/a_n100_89117# VSUBS 0.216482f
C9556 XM3/a_n158_90250# VSUBS 0.190616f
C9557 XM3/a_n100_90153# VSUBS 0.216482f
C9558 XM3/a_n158_91286# VSUBS 0.190616f
C9559 XM3/a_n100_91189# VSUBS 0.216482f
C9560 XM3/a_n158_92322# VSUBS 0.190616f
C9561 XM3/a_n100_92225# VSUBS 0.216482f
C9562 XM3/a_n158_93358# VSUBS 0.190616f
C9563 XM3/a_n100_93261# VSUBS 0.216482f
C9564 XM3/a_n158_94394# VSUBS 0.190616f
C9565 XM3/a_n100_94297# VSUBS 0.216482f
C9566 XM3/a_n158_95430# VSUBS 0.190616f
C9567 XM3/a_n100_95333# VSUBS 0.216482f
C9568 XM3/a_n158_96466# VSUBS 0.190616f
C9569 XM3/a_n100_96369# VSUBS 0.216482f
C9570 XM3/a_n158_97502# VSUBS 0.190616f
C9571 XM3/a_n100_97405# VSUBS 0.216482f
C9572 XM3/a_n158_98538# VSUBS 0.190616f
C9573 XM3/a_n100_98441# VSUBS 0.216482f
C9574 XM3/a_n158_99574# VSUBS 0.190616f
C9575 XM3/a_n100_99477# VSUBS 0.216482f
C9576 XM3/a_n158_100610# VSUBS 0.190616f
C9577 XM3/a_n100_100513# VSUBS 0.216482f
C9578 XM3/a_n158_101646# VSUBS 0.190616f
C9579 XM3/a_n100_101549# VSUBS 0.216482f
C9580 XM3/a_n158_102682# VSUBS 0.190616f
C9581 XM3/a_n100_102585# VSUBS 0.216482f
C9582 XM3/a_n158_103718# VSUBS 0.190616f
C9583 XM3/a_n100_103621# VSUBS 0.216482f
C9584 XM3/a_n158_104754# VSUBS 0.190616f
C9585 XM3/a_n100_104657# VSUBS 0.216482f
C9586 XM3/a_n158_105790# VSUBS 0.190616f
C9587 XM3/a_n100_105693# VSUBS 0.216482f
C9588 XM3/a_n158_106826# VSUBS 0.190616f
C9589 XM3/a_n100_106729# VSUBS 0.216482f
C9590 XM3/a_n158_107862# VSUBS 0.190616f
C9591 XM3/a_n100_107765# VSUBS 0.216482f
C9592 XM3/a_n158_108898# VSUBS 0.190616f
C9593 XM3/a_n100_108801# VSUBS 0.216482f
C9594 XM3/a_n158_109934# VSUBS 0.190616f
C9595 XM3/a_n100_109837# VSUBS 0.216482f
C9596 XM3/a_n158_110970# VSUBS 0.190616f
C9597 XM3/a_n100_110873# VSUBS 0.216482f
C9598 XM3/a_n158_112006# VSUBS 0.190616f
C9599 XM3/a_n100_111909# VSUBS 0.216482f
C9600 XM3/a_n158_113042# VSUBS 0.190616f
C9601 XM3/a_n100_112945# VSUBS 0.216482f
C9602 XM3/a_n158_114078# VSUBS 0.190616f
C9603 XM3/a_n100_113981# VSUBS 0.216482f
C9604 XM3/a_n158_115114# VSUBS 0.190616f
C9605 XM3/a_n100_115017# VSUBS 0.216482f
C9606 XM3/a_n158_116150# VSUBS 0.190616f
C9607 XM3/a_n100_116053# VSUBS 0.216482f
C9608 XM3/a_n158_117186# VSUBS 0.190616f
C9609 XM3/a_n100_117089# VSUBS 0.216482f
C9610 XM3/a_n158_118222# VSUBS 0.190616f
C9611 XM3/a_n100_118125# VSUBS 0.216482f
C9612 XM3/a_n158_119258# VSUBS 0.190616f
C9613 XM3/a_n100_119161# VSUBS 0.216482f
C9614 XM3/a_n158_120294# VSUBS 0.190616f
C9615 XM3/a_n100_120197# VSUBS 0.216482f
C9616 XM3/a_n158_121330# VSUBS 0.190616f
C9617 XM3/a_n100_121233# VSUBS 0.216482f
C9618 XM3/a_n158_122366# VSUBS 0.190616f
C9619 XM3/a_n100_122269# VSUBS 0.216482f
C9620 XM3/a_n158_123402# VSUBS 0.190616f
C9621 XM3/a_n100_123305# VSUBS 0.216482f
C9622 XM3/a_n158_124438# VSUBS 0.190616f
C9623 XM3/a_n100_124341# VSUBS 0.216482f
C9624 XM3/a_n158_125474# VSUBS 0.190616f
C9625 XM3/a_n100_125377# VSUBS 0.216482f
C9626 XM3/a_n158_126510# VSUBS 0.190616f
C9627 XM3/a_n100_126413# VSUBS 0.216482f
C9628 XM3/a_n158_127546# VSUBS 0.190616f
C9629 XM3/a_n100_127449# VSUBS 0.216482f
C9630 XM3/a_n158_128582# VSUBS 0.190616f
C9631 XM3/a_n100_128485# VSUBS 0.216482f
C9632 XM3/a_n158_129618# VSUBS 0.190616f
C9633 XM3/a_n100_129521# VSUBS 0.216482f
C9634 XM3/a_n158_130654# VSUBS 0.190616f
C9635 XM3/a_n100_130557# VSUBS 0.216482f
C9636 XM3/a_n158_131690# VSUBS 0.196066f
C9637 XM3/a_n100_131593# VSUBS 0.260213f
C9638 XM2/a_100_n337290# VSUBS 0.58217f
C9639 XM2/a_n158_n337290# VSUBS 0.58217f
C9640 XM2/a_n100_n337387# VSUBS 0.291162f
C9641 XM2/a_100_n334654# VSUBS 0.576721f
C9642 XM2/a_n158_n334654# VSUBS 0.576721f
C9643 XM2/a_n100_n334751# VSUBS 0.247431f
C9644 XM2/a_100_n332018# VSUBS 0.576721f
C9645 XM2/a_n158_n332018# VSUBS 0.576721f
C9646 XM2/a_n100_n332115# VSUBS 0.247431f
C9647 XM2/a_100_n329382# VSUBS 0.576721f
C9648 XM2/a_n158_n329382# VSUBS 0.576721f
C9649 XM2/a_n100_n329479# VSUBS 0.247431f
C9650 XM2/a_100_n326746# VSUBS 0.576721f
C9651 XM2/a_n158_n326746# VSUBS 0.576721f
C9652 XM2/a_n100_n326843# VSUBS 0.247431f
C9653 XM2/a_100_n324110# VSUBS 0.576721f
C9654 XM2/a_n158_n324110# VSUBS 0.576721f
C9655 XM2/a_n100_n324207# VSUBS 0.247431f
C9656 XM2/a_100_n321474# VSUBS 0.576721f
C9657 XM2/a_n158_n321474# VSUBS 0.576721f
C9658 XM2/a_n100_n321571# VSUBS 0.247431f
C9659 XM2/a_100_n318838# VSUBS 0.576721f
C9660 XM2/a_n158_n318838# VSUBS 0.576721f
C9661 XM2/a_n100_n318935# VSUBS 0.247431f
C9662 XM2/a_100_n316202# VSUBS 0.576721f
C9663 XM2/a_n158_n316202# VSUBS 0.576721f
C9664 XM2/a_n100_n316299# VSUBS 0.247431f
C9665 XM2/a_100_n313566# VSUBS 0.576721f
C9666 XM2/a_n158_n313566# VSUBS 0.576721f
C9667 XM2/a_n100_n313663# VSUBS 0.247431f
C9668 XM2/a_100_n310930# VSUBS 0.576721f
C9669 XM2/a_n158_n310930# VSUBS 0.576721f
C9670 XM2/a_n100_n311027# VSUBS 0.247431f
C9671 XM2/a_100_n308294# VSUBS 0.576721f
C9672 XM2/a_n158_n308294# VSUBS 0.576721f
C9673 XM2/a_n100_n308391# VSUBS 0.247431f
C9674 XM2/a_100_n305658# VSUBS 0.576721f
C9675 XM2/a_n158_n305658# VSUBS 0.576721f
C9676 XM2/a_n100_n305755# VSUBS 0.247431f
C9677 XM2/a_100_n303022# VSUBS 0.576721f
C9678 XM2/a_n158_n303022# VSUBS 0.576721f
C9679 XM2/a_n100_n303119# VSUBS 0.247431f
C9680 XM2/a_100_n300386# VSUBS 0.576721f
C9681 XM2/a_n158_n300386# VSUBS 0.576721f
C9682 XM2/a_n100_n300483# VSUBS 0.247431f
C9683 XM2/a_100_n297750# VSUBS 0.576721f
C9684 XM2/a_n158_n297750# VSUBS 0.576721f
C9685 XM2/a_n100_n297847# VSUBS 0.247431f
C9686 XM2/a_100_n295114# VSUBS 0.576721f
C9687 XM2/a_n158_n295114# VSUBS 0.576721f
C9688 XM2/a_n100_n295211# VSUBS 0.247431f
C9689 XM2/a_100_n292478# VSUBS 0.576721f
C9690 XM2/a_n158_n292478# VSUBS 0.576721f
C9691 XM2/a_n100_n292575# VSUBS 0.247431f
C9692 XM2/a_100_n289842# VSUBS 0.576721f
C9693 XM2/a_n158_n289842# VSUBS 0.576721f
C9694 XM2/a_n100_n289939# VSUBS 0.247431f
C9695 XM2/a_100_n287206# VSUBS 0.576721f
C9696 XM2/a_n158_n287206# VSUBS 0.576721f
C9697 XM2/a_n100_n287303# VSUBS 0.247431f
C9698 XM2/a_100_n284570# VSUBS 0.576721f
C9699 XM2/a_n158_n284570# VSUBS 0.576721f
C9700 XM2/a_n100_n284667# VSUBS 0.247431f
C9701 XM2/a_100_n281934# VSUBS 0.576721f
C9702 XM2/a_n158_n281934# VSUBS 0.576721f
C9703 XM2/a_n100_n282031# VSUBS 0.247431f
C9704 XM2/a_100_n279298# VSUBS 0.576721f
C9705 XM2/a_n158_n279298# VSUBS 0.576721f
C9706 XM2/a_n100_n279395# VSUBS 0.247431f
C9707 XM2/a_100_n276662# VSUBS 0.576721f
C9708 XM2/a_n158_n276662# VSUBS 0.576721f
C9709 XM2/a_n100_n276759# VSUBS 0.247431f
C9710 XM2/a_100_n274026# VSUBS 0.576721f
C9711 XM2/a_n158_n274026# VSUBS 0.576721f
C9712 XM2/a_n100_n274123# VSUBS 0.247431f
C9713 XM2/a_100_n271390# VSUBS 0.576721f
C9714 XM2/a_n158_n271390# VSUBS 0.576721f
C9715 XM2/a_n100_n271487# VSUBS 0.247431f
C9716 XM2/a_100_n268754# VSUBS 0.576721f
C9717 XM2/a_n158_n268754# VSUBS 0.576721f
C9718 XM2/a_n100_n268851# VSUBS 0.247431f
C9719 XM2/a_100_n266118# VSUBS 0.576721f
C9720 XM2/a_n158_n266118# VSUBS 0.576721f
C9721 XM2/a_n100_n266215# VSUBS 0.247431f
C9722 XM2/a_100_n263482# VSUBS 0.576721f
C9723 XM2/a_n158_n263482# VSUBS 0.576721f
C9724 XM2/a_n100_n263579# VSUBS 0.247431f
C9725 XM2/a_100_n260846# VSUBS 0.576721f
C9726 XM2/a_n158_n260846# VSUBS 0.576721f
C9727 XM2/a_n100_n260943# VSUBS 0.247431f
C9728 XM2/a_100_n258210# VSUBS 0.576721f
C9729 XM2/a_n158_n258210# VSUBS 0.576721f
C9730 XM2/a_n100_n258307# VSUBS 0.247431f
C9731 XM2/a_100_n255574# VSUBS 0.576721f
C9732 XM2/a_n158_n255574# VSUBS 0.576721f
C9733 XM2/a_n100_n255671# VSUBS 0.247431f
C9734 XM2/a_100_n252938# VSUBS 0.576721f
C9735 XM2/a_n158_n252938# VSUBS 0.576721f
C9736 XM2/a_n100_n253035# VSUBS 0.247431f
C9737 XM2/a_100_n250302# VSUBS 0.576721f
C9738 XM2/a_n158_n250302# VSUBS 0.576721f
C9739 XM2/a_n100_n250399# VSUBS 0.247431f
C9740 XM2/a_100_n247666# VSUBS 0.576721f
C9741 XM2/a_n158_n247666# VSUBS 0.576721f
C9742 XM2/a_n100_n247763# VSUBS 0.247431f
C9743 XM2/a_100_n245030# VSUBS 0.576721f
C9744 XM2/a_n158_n245030# VSUBS 0.576721f
C9745 XM2/a_n100_n245127# VSUBS 0.247431f
C9746 XM2/a_100_n242394# VSUBS 0.576721f
C9747 XM2/a_n158_n242394# VSUBS 0.576721f
C9748 XM2/a_n100_n242491# VSUBS 0.247431f
C9749 XM2/a_100_n239758# VSUBS 0.576721f
C9750 XM2/a_n158_n239758# VSUBS 0.576721f
C9751 XM2/a_n100_n239855# VSUBS 0.247431f
C9752 XM2/a_100_n237122# VSUBS 0.576721f
C9753 XM2/a_n158_n237122# VSUBS 0.576721f
C9754 XM2/a_n100_n237219# VSUBS 0.247431f
C9755 XM2/a_100_n234486# VSUBS 0.576721f
C9756 XM2/a_n158_n234486# VSUBS 0.576721f
C9757 XM2/a_n100_n234583# VSUBS 0.247431f
C9758 XM2/a_100_n231850# VSUBS 0.576721f
C9759 XM2/a_n158_n231850# VSUBS 0.576721f
C9760 XM2/a_n100_n231947# VSUBS 0.247431f
C9761 XM2/a_100_n229214# VSUBS 0.576721f
C9762 XM2/a_n158_n229214# VSUBS 0.576721f
C9763 XM2/a_n100_n229311# VSUBS 0.247431f
C9764 XM2/a_100_n226578# VSUBS 0.576721f
C9765 XM2/a_n158_n226578# VSUBS 0.576721f
C9766 XM2/a_n100_n226675# VSUBS 0.247431f
C9767 XM2/a_100_n223942# VSUBS 0.576721f
C9768 XM2/a_n158_n223942# VSUBS 0.576721f
C9769 XM2/a_n100_n224039# VSUBS 0.247431f
C9770 XM2/a_100_n221306# VSUBS 0.576721f
C9771 XM2/a_n158_n221306# VSUBS 0.576721f
C9772 XM2/a_n100_n221403# VSUBS 0.247431f
C9773 XM2/a_100_n218670# VSUBS 0.576721f
C9774 XM2/a_n158_n218670# VSUBS 0.576721f
C9775 XM2/a_n100_n218767# VSUBS 0.247431f
C9776 XM2/a_100_n216034# VSUBS 0.576721f
C9777 XM2/a_n158_n216034# VSUBS 0.576721f
C9778 XM2/a_n100_n216131# VSUBS 0.247431f
C9779 XM2/a_100_n213398# VSUBS 0.576721f
C9780 XM2/a_n158_n213398# VSUBS 0.576721f
C9781 XM2/a_n100_n213495# VSUBS 0.247431f
C9782 XM2/a_100_n210762# VSUBS 0.576721f
C9783 XM2/a_n158_n210762# VSUBS 0.576721f
C9784 XM2/a_n100_n210859# VSUBS 0.247431f
C9785 XM2/a_100_n208126# VSUBS 0.576721f
C9786 XM2/a_n158_n208126# VSUBS 0.576721f
C9787 XM2/a_n100_n208223# VSUBS 0.247431f
C9788 XM2/a_100_n205490# VSUBS 0.576721f
C9789 XM2/a_n158_n205490# VSUBS 0.576721f
C9790 XM2/a_n100_n205587# VSUBS 0.247431f
C9791 XM2/a_100_n202854# VSUBS 0.576721f
C9792 XM2/a_n158_n202854# VSUBS 0.576721f
C9793 XM2/a_n100_n202951# VSUBS 0.247431f
C9794 XM2/a_100_n200218# VSUBS 0.576721f
C9795 XM2/a_n158_n200218# VSUBS 0.576721f
C9796 XM2/a_n100_n200315# VSUBS 0.247431f
C9797 XM2/a_100_n197582# VSUBS 0.576721f
C9798 XM2/a_n158_n197582# VSUBS 0.576721f
C9799 XM2/a_n100_n197679# VSUBS 0.247431f
C9800 XM2/a_100_n194946# VSUBS 0.576721f
C9801 XM2/a_n158_n194946# VSUBS 0.576721f
C9802 XM2/a_n100_n195043# VSUBS 0.247431f
C9803 XM2/a_100_n192310# VSUBS 0.576721f
C9804 XM2/a_n158_n192310# VSUBS 0.576721f
C9805 XM2/a_n100_n192407# VSUBS 0.247431f
C9806 XM2/a_100_n189674# VSUBS 0.576721f
C9807 XM2/a_n158_n189674# VSUBS 0.576721f
C9808 XM2/a_n100_n189771# VSUBS 0.247431f
C9809 XM2/a_100_n187038# VSUBS 0.576721f
C9810 XM2/a_n158_n187038# VSUBS 0.576721f
C9811 XM2/a_n100_n187135# VSUBS 0.247431f
C9812 XM2/a_100_n184402# VSUBS 0.576721f
C9813 XM2/a_n158_n184402# VSUBS 0.576721f
C9814 XM2/a_n100_n184499# VSUBS 0.247431f
C9815 XM2/a_100_n181766# VSUBS 0.576721f
C9816 XM2/a_n158_n181766# VSUBS 0.576721f
C9817 XM2/a_n100_n181863# VSUBS 0.247431f
C9818 XM2/a_100_n179130# VSUBS 0.576721f
C9819 XM2/a_n158_n179130# VSUBS 0.576721f
C9820 XM2/a_n100_n179227# VSUBS 0.247431f
C9821 XM2/a_100_n176494# VSUBS 0.576721f
C9822 XM2/a_n158_n176494# VSUBS 0.576721f
C9823 XM2/a_n100_n176591# VSUBS 0.247431f
C9824 XM2/a_100_n173858# VSUBS 0.576721f
C9825 XM2/a_n158_n173858# VSUBS 0.576721f
C9826 XM2/a_n100_n173955# VSUBS 0.247431f
C9827 XM2/a_100_n171222# VSUBS 0.576721f
C9828 XM2/a_n158_n171222# VSUBS 0.576721f
C9829 XM2/a_n100_n171319# VSUBS 0.247431f
C9830 XM2/a_100_n168586# VSUBS 0.576721f
C9831 XM2/a_n158_n168586# VSUBS 0.576721f
C9832 XM2/a_n100_n168683# VSUBS 0.247431f
C9833 XM2/a_100_n165950# VSUBS 0.576721f
C9834 XM2/a_n158_n165950# VSUBS 0.576721f
C9835 XM2/a_n100_n166047# VSUBS 0.247431f
C9836 XM2/a_100_n163314# VSUBS 0.576721f
C9837 XM2/a_n158_n163314# VSUBS 0.576721f
C9838 XM2/a_n100_n163411# VSUBS 0.247431f
C9839 XM2/a_100_n160678# VSUBS 0.576721f
C9840 XM2/a_n158_n160678# VSUBS 0.576721f
C9841 XM2/a_n100_n160775# VSUBS 0.247431f
C9842 XM2/a_100_n158042# VSUBS 0.576721f
C9843 XM2/a_n158_n158042# VSUBS 0.576721f
C9844 XM2/a_n100_n158139# VSUBS 0.247431f
C9845 XM2/a_100_n155406# VSUBS 0.576721f
C9846 XM2/a_n158_n155406# VSUBS 0.576721f
C9847 XM2/a_n100_n155503# VSUBS 0.247431f
C9848 XM2/a_100_n152770# VSUBS 0.576721f
C9849 XM2/a_n158_n152770# VSUBS 0.576721f
C9850 XM2/a_n100_n152867# VSUBS 0.247431f
C9851 XM2/a_100_n150134# VSUBS 0.576721f
C9852 XM2/a_n158_n150134# VSUBS 0.576721f
C9853 XM2/a_n100_n150231# VSUBS 0.247431f
C9854 XM2/a_100_n147498# VSUBS 0.576721f
C9855 XM2/a_n158_n147498# VSUBS 0.576721f
C9856 XM2/a_n100_n147595# VSUBS 0.247431f
C9857 XM2/a_100_n144862# VSUBS 0.576721f
C9858 XM2/a_n158_n144862# VSUBS 0.576721f
C9859 XM2/a_n100_n144959# VSUBS 0.247431f
C9860 XM2/a_100_n142226# VSUBS 0.576721f
C9861 XM2/a_n158_n142226# VSUBS 0.576721f
C9862 XM2/a_n100_n142323# VSUBS 0.247431f
C9863 XM2/a_100_n139590# VSUBS 0.576721f
C9864 XM2/a_n158_n139590# VSUBS 0.576721f
C9865 XM2/a_n100_n139687# VSUBS 0.247431f
C9866 XM2/a_100_n136954# VSUBS 0.576721f
C9867 XM2/a_n158_n136954# VSUBS 0.576721f
C9868 XM2/a_n100_n137051# VSUBS 0.247431f
C9869 XM2/a_100_n134318# VSUBS 0.576721f
C9870 XM2/a_n158_n134318# VSUBS 0.576721f
C9871 XM2/a_n100_n134415# VSUBS 0.247431f
C9872 XM2/a_100_n131682# VSUBS 0.576721f
C9873 XM2/a_n158_n131682# VSUBS 0.576721f
C9874 XM2/a_n100_n131779# VSUBS 0.247431f
C9875 XM2/a_100_n129046# VSUBS 0.576721f
C9876 XM2/a_n158_n129046# VSUBS 0.576721f
C9877 XM2/a_n100_n129143# VSUBS 0.247431f
C9878 XM2/a_100_n126410# VSUBS 0.576721f
C9879 XM2/a_n158_n126410# VSUBS 0.576721f
C9880 XM2/a_n100_n126507# VSUBS 0.247431f
C9881 XM2/a_100_n123774# VSUBS 0.576721f
C9882 XM2/a_n158_n123774# VSUBS 0.576721f
C9883 XM2/a_n100_n123871# VSUBS 0.247431f
C9884 XM2/a_100_n121138# VSUBS 0.576721f
C9885 XM2/a_n158_n121138# VSUBS 0.576721f
C9886 XM2/a_n100_n121235# VSUBS 0.247431f
C9887 XM2/a_100_n118502# VSUBS 0.576721f
C9888 XM2/a_n158_n118502# VSUBS 0.576721f
C9889 XM2/a_n100_n118599# VSUBS 0.247431f
C9890 XM2/a_100_n115866# VSUBS 0.576721f
C9891 XM2/a_n158_n115866# VSUBS 0.576721f
C9892 XM2/a_n100_n115963# VSUBS 0.247431f
C9893 XM2/a_100_n113230# VSUBS 0.576721f
C9894 XM2/a_n158_n113230# VSUBS 0.576721f
C9895 XM2/a_n100_n113327# VSUBS 0.247431f
C9896 XM2/a_100_n110594# VSUBS 0.576721f
C9897 XM2/a_n158_n110594# VSUBS 0.576721f
C9898 XM2/a_n100_n110691# VSUBS 0.247431f
C9899 XM2/a_100_n107958# VSUBS 0.576721f
C9900 XM2/a_n158_n107958# VSUBS 0.576721f
C9901 XM2/a_n100_n108055# VSUBS 0.247431f
C9902 XM2/a_100_n105322# VSUBS 0.576721f
C9903 XM2/a_n158_n105322# VSUBS 0.576721f
C9904 XM2/a_n100_n105419# VSUBS 0.247431f
C9905 XM2/a_100_n102686# VSUBS 0.576721f
C9906 XM2/a_n158_n102686# VSUBS 0.576721f
C9907 XM2/a_n100_n102783# VSUBS 0.247431f
C9908 XM2/a_100_n100050# VSUBS 0.576721f
C9909 XM2/a_n158_n100050# VSUBS 0.576721f
C9910 XM2/a_n100_n100147# VSUBS 0.247431f
C9911 XM2/a_100_n97414# VSUBS 0.576721f
C9912 XM2/a_n158_n97414# VSUBS 0.576721f
C9913 XM2/a_n100_n97511# VSUBS 0.247431f
C9914 XM2/a_100_n94778# VSUBS 0.576721f
C9915 XM2/a_n158_n94778# VSUBS 0.576721f
C9916 XM2/a_n100_n94875# VSUBS 0.247431f
C9917 XM2/a_100_n92142# VSUBS 0.576721f
C9918 XM2/a_n158_n92142# VSUBS 0.576721f
C9919 XM2/a_n100_n92239# VSUBS 0.247431f
C9920 XM2/a_100_n89506# VSUBS 0.576721f
C9921 XM2/a_n158_n89506# VSUBS 0.576721f
C9922 XM2/a_n100_n89603# VSUBS 0.247431f
C9923 XM2/a_100_n86870# VSUBS 0.576721f
C9924 XM2/a_n158_n86870# VSUBS 0.576721f
C9925 XM2/a_n100_n86967# VSUBS 0.247431f
C9926 XM2/a_100_n84234# VSUBS 0.576721f
C9927 XM2/a_n158_n84234# VSUBS 0.576721f
C9928 XM2/a_n100_n84331# VSUBS 0.247431f
C9929 XM2/a_100_n81598# VSUBS 0.576721f
C9930 XM2/a_n158_n81598# VSUBS 0.576721f
C9931 XM2/a_n100_n81695# VSUBS 0.247431f
C9932 XM2/a_100_n78962# VSUBS 0.576721f
C9933 XM2/a_n158_n78962# VSUBS 0.576721f
C9934 XM2/a_n100_n79059# VSUBS 0.247431f
C9935 XM2/a_100_n76326# VSUBS 0.576721f
C9936 XM2/a_n158_n76326# VSUBS 0.576721f
C9937 XM2/a_n100_n76423# VSUBS 0.247431f
C9938 XM2/a_100_n73690# VSUBS 0.576721f
C9939 XM2/a_n158_n73690# VSUBS 0.576721f
C9940 XM2/a_n100_n73787# VSUBS 0.247431f
C9941 XM2/a_100_n71054# VSUBS 0.576721f
C9942 XM2/a_n158_n71054# VSUBS 0.576721f
C9943 XM2/a_n100_n71151# VSUBS 0.247431f
C9944 XM2/a_100_n68418# VSUBS 0.576721f
C9945 XM2/a_n158_n68418# VSUBS 0.576721f
C9946 XM2/a_n100_n68515# VSUBS 0.247431f
C9947 XM2/a_100_n65782# VSUBS 0.576721f
C9948 XM2/a_n158_n65782# VSUBS 0.576721f
C9949 XM2/a_n100_n65879# VSUBS 0.247431f
C9950 XM2/a_100_n63146# VSUBS 0.576721f
C9951 XM2/a_n158_n63146# VSUBS 0.576721f
C9952 XM2/a_n100_n63243# VSUBS 0.247431f
C9953 XM2/a_100_n60510# VSUBS 0.576721f
C9954 XM2/a_n158_n60510# VSUBS 0.576721f
C9955 XM2/a_n100_n60607# VSUBS 0.247431f
C9956 XM2/a_100_n57874# VSUBS 0.576721f
C9957 XM2/a_n158_n57874# VSUBS 0.576721f
C9958 XM2/a_n100_n57971# VSUBS 0.247431f
C9959 XM2/a_100_n55238# VSUBS 0.576721f
C9960 XM2/a_n158_n55238# VSUBS 0.576721f
C9961 XM2/a_n100_n55335# VSUBS 0.247431f
C9962 XM2/a_100_n52602# VSUBS 0.576721f
C9963 XM2/a_n158_n52602# VSUBS 0.576721f
C9964 XM2/a_n100_n52699# VSUBS 0.247431f
C9965 XM2/a_100_n49966# VSUBS 0.576721f
C9966 XM2/a_n158_n49966# VSUBS 0.576721f
C9967 XM2/a_n100_n50063# VSUBS 0.247431f
C9968 XM2/a_100_n47330# VSUBS 0.576721f
C9969 XM2/a_n158_n47330# VSUBS 0.576721f
C9970 XM2/a_n100_n47427# VSUBS 0.247431f
C9971 XM2/a_100_n44694# VSUBS 0.576721f
C9972 XM2/a_n158_n44694# VSUBS 0.576721f
C9973 XM2/a_n100_n44791# VSUBS 0.247431f
C9974 XM2/a_100_n42058# VSUBS 0.576721f
C9975 XM2/a_n158_n42058# VSUBS 0.576721f
C9976 XM2/a_n100_n42155# VSUBS 0.247431f
C9977 XM2/a_100_n39422# VSUBS 0.576721f
C9978 XM2/a_n158_n39422# VSUBS 0.576721f
C9979 XM2/a_n100_n39519# VSUBS 0.247431f
C9980 XM2/a_100_n36786# VSUBS 0.576721f
C9981 XM2/a_n158_n36786# VSUBS 0.576721f
C9982 XM2/a_n100_n36883# VSUBS 0.247431f
C9983 XM2/a_100_n34150# VSUBS 0.576721f
C9984 XM2/a_n158_n34150# VSUBS 0.576721f
C9985 XM2/a_n100_n34247# VSUBS 0.247431f
C9986 XM2/a_100_n31514# VSUBS 0.576721f
C9987 XM2/a_n158_n31514# VSUBS 0.576721f
C9988 XM2/a_n100_n31611# VSUBS 0.247431f
C9989 XM2/a_100_n28878# VSUBS 0.576721f
C9990 XM2/a_n158_n28878# VSUBS 0.576721f
C9991 XM2/a_n100_n28975# VSUBS 0.247431f
C9992 XM2/a_100_n26242# VSUBS 0.576721f
C9993 XM2/a_n158_n26242# VSUBS 0.576721f
C9994 XM2/a_n100_n26339# VSUBS 0.247431f
C9995 XM2/a_100_n23606# VSUBS 0.576721f
C9996 XM2/a_n158_n23606# VSUBS 0.576721f
C9997 XM2/a_n100_n23703# VSUBS 0.247431f
C9998 XM2/a_100_n20970# VSUBS 0.576721f
C9999 XM2/a_n158_n20970# VSUBS 0.576721f
C10000 XM2/a_n100_n21067# VSUBS 0.247431f
C10001 XM2/a_100_n18334# VSUBS 0.576721f
C10002 XM2/a_n158_n18334# VSUBS 0.576721f
C10003 XM2/a_n100_n18431# VSUBS 0.247431f
C10004 XM2/a_100_n15698# VSUBS 0.576721f
C10005 XM2/a_n158_n15698# VSUBS 0.576721f
C10006 XM2/a_n100_n15795# VSUBS 0.247431f
C10007 XM2/a_100_n13062# VSUBS 0.576721f
C10008 XM2/a_n158_n13062# VSUBS 0.576721f
C10009 XM2/a_n100_n13159# VSUBS 0.247431f
C10010 XM2/a_100_n10426# VSUBS 0.576721f
C10011 XM2/a_n158_n10426# VSUBS 0.576721f
C10012 XM2/a_n100_n10523# VSUBS 0.247431f
C10013 XM2/a_100_n7790# VSUBS 0.576721f
C10014 XM2/a_n158_n7790# VSUBS 0.576721f
C10015 XM2/a_n100_n7887# VSUBS 0.247431f
C10016 XM2/a_100_n5154# VSUBS 0.576721f
C10017 XM2/a_n158_n5154# VSUBS 0.576721f
C10018 XM2/a_n100_n5251# VSUBS 0.247431f
C10019 XM2/a_100_n2518# VSUBS 0.576721f
C10020 XM2/a_n158_n2518# VSUBS 0.576721f
C10021 XM2/a_n100_n2615# VSUBS 0.247431f
C10022 XM2/a_100_118# VSUBS 0.576721f
C10023 XM2/a_n158_118# VSUBS 0.576721f
C10024 XM2/a_n100_21# VSUBS 0.247431f
C10025 XM2/a_100_2754# VSUBS 0.576721f
C10026 XM2/a_n158_2754# VSUBS 0.576721f
C10027 XM2/a_n100_2657# VSUBS 0.247431f
C10028 XM2/a_100_5390# VSUBS 0.576721f
C10029 XM2/a_n158_5390# VSUBS 0.576721f
C10030 XM2/a_n100_5293# VSUBS 0.247431f
C10031 XM2/a_100_8026# VSUBS 0.576721f
C10032 XM2/a_n158_8026# VSUBS 0.576721f
C10033 XM2/a_n100_7929# VSUBS 0.247431f
C10034 XM2/a_100_10662# VSUBS 0.576721f
C10035 XM2/a_n158_10662# VSUBS 0.576721f
C10036 XM2/a_n100_10565# VSUBS 0.247431f
C10037 XM2/a_100_13298# VSUBS 0.576721f
C10038 XM2/a_n158_13298# VSUBS 0.576721f
C10039 XM2/a_n100_13201# VSUBS 0.247431f
C10040 XM2/a_100_15934# VSUBS 0.576721f
C10041 XM2/a_n158_15934# VSUBS 0.576721f
C10042 XM2/a_n100_15837# VSUBS 0.247431f
C10043 XM2/a_100_18570# VSUBS 0.576721f
C10044 XM2/a_n158_18570# VSUBS 0.576721f
C10045 XM2/a_n100_18473# VSUBS 0.247431f
C10046 XM2/a_100_21206# VSUBS 0.576721f
C10047 XM2/a_n158_21206# VSUBS 0.576721f
C10048 XM2/a_n100_21109# VSUBS 0.247431f
C10049 XM2/a_100_23842# VSUBS 0.576721f
C10050 XM2/a_n158_23842# VSUBS 0.576721f
C10051 XM2/a_n100_23745# VSUBS 0.247431f
C10052 XM2/a_100_26478# VSUBS 0.576721f
C10053 XM2/a_n158_26478# VSUBS 0.576721f
C10054 XM2/a_n100_26381# VSUBS 0.247431f
C10055 XM2/a_100_29114# VSUBS 0.576721f
C10056 XM2/a_n158_29114# VSUBS 0.576721f
C10057 XM2/a_n100_29017# VSUBS 0.247431f
C10058 XM2/a_100_31750# VSUBS 0.576721f $ **FLOATING
C10059 XM2/a_n158_31750# VSUBS 0.576721f $ **FLOATING
C10060 XM2/a_n100_31653# VSUBS 0.247431f $ **FLOATING
C10061 XM2/a_100_34386# VSUBS 0.576721f $ **FLOATING
C10062 XM2/a_n158_34386# VSUBS 0.576721f $ **FLOATING
C10063 XM2/a_n100_34289# VSUBS 0.247431f $ **FLOATING
C10064 XM2/a_100_37022# VSUBS 0.576721f $ **FLOATING
C10065 XM2/a_n158_37022# VSUBS 0.576721f $ **FLOATING
C10066 XM2/a_n100_36925# VSUBS 0.247431f $ **FLOATING
C10067 XM2/a_100_39658# VSUBS 0.576721f $ **FLOATING
C10068 XM2/a_n158_39658# VSUBS 0.576721f $ **FLOATING
C10069 XM2/a_n100_39561# VSUBS 0.247431f $ **FLOATING
C10070 XM2/a_100_42294# VSUBS 0.576721f $ **FLOATING
C10071 XM2/a_n158_42294# VSUBS 0.576721f $ **FLOATING
C10072 XM2/a_n100_42197# VSUBS 0.247431f $ **FLOATING
C10073 XM2/a_100_44930# VSUBS 0.576721f $ **FLOATING
C10074 XM2/a_n158_44930# VSUBS 0.576721f $ **FLOATING
C10075 XM2/a_n100_44833# VSUBS 0.247431f $ **FLOATING
C10076 XM2/a_100_47566# VSUBS 0.576721f $ **FLOATING
C10077 XM2/a_n158_47566# VSUBS 0.576721f $ **FLOATING
C10078 XM2/a_n100_47469# VSUBS 0.247431f $ **FLOATING
C10079 XM2/a_100_50202# VSUBS 0.576721f $ **FLOATING
C10080 XM2/a_n158_50202# VSUBS 0.576721f $ **FLOATING
C10081 XM2/a_n100_50105# VSUBS 0.247431f $ **FLOATING
C10082 XM2/a_100_52838# VSUBS 0.576721f $ **FLOATING
C10083 XM2/a_n158_52838# VSUBS 0.576721f $ **FLOATING
C10084 XM2/a_n100_52741# VSUBS 0.247431f $ **FLOATING
C10085 XM2/a_100_55474# VSUBS 0.576721f $ **FLOATING
C10086 XM2/a_n158_55474# VSUBS 0.576721f $ **FLOATING
C10087 XM2/a_n100_55377# VSUBS 0.247431f $ **FLOATING
C10088 XM2/a_100_58110# VSUBS 0.576721f $ **FLOATING
C10089 XM2/a_n158_58110# VSUBS 0.576721f $ **FLOATING
C10090 XM2/a_n100_58013# VSUBS 0.247431f $ **FLOATING
C10091 XM2/a_100_60746# VSUBS 0.576721f $ **FLOATING
C10092 XM2/a_n158_60746# VSUBS 0.576721f $ **FLOATING
C10093 XM2/a_n100_60649# VSUBS 0.247431f $ **FLOATING
C10094 XM2/a_100_63382# VSUBS 0.576721f $ **FLOATING
C10095 XM2/a_n158_63382# VSUBS 0.576721f $ **FLOATING
C10096 XM2/a_n100_63285# VSUBS 0.247431f $ **FLOATING
C10097 XM2/a_100_66018# VSUBS 0.576721f $ **FLOATING
C10098 XM2/a_n158_66018# VSUBS 0.576721f $ **FLOATING
C10099 XM2/a_n100_65921# VSUBS 0.247431f $ **FLOATING
C10100 XM2/a_100_68654# VSUBS 0.576721f $ **FLOATING
C10101 XM2/a_n158_68654# VSUBS 0.576721f $ **FLOATING
C10102 XM2/a_n100_68557# VSUBS 0.247431f $ **FLOATING
C10103 XM2/a_100_71290# VSUBS 0.576721f $ **FLOATING
C10104 XM2/a_n158_71290# VSUBS 0.576721f $ **FLOATING
C10105 XM2/a_n100_71193# VSUBS 0.247431f $ **FLOATING
C10106 XM2/a_100_73926# VSUBS 0.576721f $ **FLOATING
C10107 XM2/a_n158_73926# VSUBS 0.576721f $ **FLOATING
C10108 XM2/a_n100_73829# VSUBS 0.247431f $ **FLOATING
C10109 XM2/a_100_76562# VSUBS 0.576721f $ **FLOATING
C10110 XM2/a_n158_76562# VSUBS 0.576721f $ **FLOATING
C10111 XM2/a_n100_76465# VSUBS 0.247431f $ **FLOATING
C10112 XM2/a_100_79198# VSUBS 0.576721f $ **FLOATING
C10113 XM2/a_n158_79198# VSUBS 0.576721f $ **FLOATING
C10114 XM2/a_n100_79101# VSUBS 0.247431f $ **FLOATING
C10115 XM2/a_100_81834# VSUBS 0.576721f $ **FLOATING
C10116 XM2/a_n158_81834# VSUBS 0.576721f $ **FLOATING
C10117 XM2/a_n100_81737# VSUBS 0.247431f $ **FLOATING
C10118 XM2/a_100_84470# VSUBS 0.576721f $ **FLOATING
C10119 XM2/a_n158_84470# VSUBS 0.576721f $ **FLOATING
C10120 XM2/a_n100_84373# VSUBS 0.247431f $ **FLOATING
C10121 XM2/a_100_87106# VSUBS 0.576721f $ **FLOATING
C10122 XM2/a_n158_87106# VSUBS 0.576721f $ **FLOATING
C10123 XM2/a_n100_87009# VSUBS 0.247431f $ **FLOATING
C10124 XM2/a_100_89742# VSUBS 0.576721f $ **FLOATING
C10125 XM2/a_n158_89742# VSUBS 0.576721f $ **FLOATING
C10126 XM2/a_n100_89645# VSUBS 0.247431f $ **FLOATING
C10127 XM2/a_100_92378# VSUBS 0.576721f $ **FLOATING
C10128 XM2/a_n158_92378# VSUBS 0.576721f $ **FLOATING
C10129 XM2/a_n100_92281# VSUBS 0.247431f $ **FLOATING
C10130 XM2/a_100_95014# VSUBS 0.576721f $ **FLOATING
C10131 XM2/a_n158_95014# VSUBS 0.576721f $ **FLOATING
C10132 XM2/a_n100_94917# VSUBS 0.247431f $ **FLOATING
C10133 XM2/a_100_97650# VSUBS 0.576721f $ **FLOATING
C10134 XM2/a_n158_97650# VSUBS 0.576721f $ **FLOATING
C10135 XM2/a_n100_97553# VSUBS 0.247431f $ **FLOATING
C10136 XM2/a_100_100286# VSUBS 0.576721f $ **FLOATING
C10137 XM2/a_n158_100286# VSUBS 0.576721f $ **FLOATING
C10138 XM2/a_n100_100189# VSUBS 0.247431f $ **FLOATING
C10139 XM2/a_100_102922# VSUBS 0.576721f $ **FLOATING
C10140 XM2/a_n158_102922# VSUBS 0.576721f $ **FLOATING
C10141 XM2/a_n100_102825# VSUBS 0.247431f $ **FLOATING
C10142 XM2/a_100_105558# VSUBS 0.576721f $ **FLOATING
C10143 XM2/a_n158_105558# VSUBS 0.576721f $ **FLOATING
C10144 XM2/a_n100_105461# VSUBS 0.247431f $ **FLOATING
C10145 XM2/a_100_108194# VSUBS 0.576721f $ **FLOATING
C10146 XM2/a_n158_108194# VSUBS 0.576721f $ **FLOATING
C10147 XM2/a_n100_108097# VSUBS 0.247431f $ **FLOATING
C10148 XM2/a_100_110830# VSUBS 0.576721f $ **FLOATING
C10149 XM2/a_n158_110830# VSUBS 0.576721f $ **FLOATING
C10150 XM2/a_n100_110733# VSUBS 0.247431f $ **FLOATING
C10151 XM2/a_100_113466# VSUBS 0.576721f $ **FLOATING
C10152 XM2/a_n158_113466# VSUBS 0.576721f $ **FLOATING
C10153 XM2/a_n100_113369# VSUBS 0.247431f $ **FLOATING
C10154 XM2/a_100_116102# VSUBS 0.576721f $ **FLOATING
C10155 XM2/a_n158_116102# VSUBS 0.576721f $ **FLOATING
C10156 XM2/a_n100_116005# VSUBS 0.247431f $ **FLOATING
C10157 XM2/a_100_118738# VSUBS 0.576721f $ **FLOATING
C10158 XM2/a_n158_118738# VSUBS 0.576721f $ **FLOATING
C10159 XM2/a_n100_118641# VSUBS 0.247431f $ **FLOATING
C10160 XM2/a_100_121374# VSUBS 0.576721f $ **FLOATING
C10161 XM2/a_n158_121374# VSUBS 0.576721f $ **FLOATING
C10162 XM2/a_n100_121277# VSUBS 0.247431f $ **FLOATING
C10163 XM2/a_100_124010# VSUBS 0.576721f $ **FLOATING
C10164 XM2/a_n158_124010# VSUBS 0.576721f $ **FLOATING
C10165 XM2/a_n100_123913# VSUBS 0.247431f $ **FLOATING
C10166 XM2/a_100_126646# VSUBS 0.576721f $ **FLOATING
C10167 XM2/a_n158_126646# VSUBS 0.576721f $ **FLOATING
C10168 XM2/a_n100_126549# VSUBS 0.247431f $ **FLOATING
C10169 XM2/a_100_129282# VSUBS 0.576721f $ **FLOATING
C10170 XM2/a_n158_129282# VSUBS 0.576721f $ **FLOATING
C10171 XM2/a_n100_129185# VSUBS 0.247431f $ **FLOATING
C10172 XM2/a_100_131918# VSUBS 0.576721f $ **FLOATING
C10173 XM2/a_n158_131918# VSUBS 0.576721f $ **FLOATING
C10174 XM2/a_n100_131821# VSUBS 0.247431f $ **FLOATING
C10175 XM2/a_100_134554# VSUBS 0.576721f $ **FLOATING
C10176 XM2/a_n158_134554# VSUBS 0.576721f $ **FLOATING
C10177 XM2/a_n100_134457# VSUBS 0.247431f $ **FLOATING
C10178 XM2/a_100_137190# VSUBS 0.576721f $ **FLOATING
C10179 XM2/a_n158_137190# VSUBS 0.576721f $ **FLOATING
C10180 XM2/a_n100_137093# VSUBS 0.247431f $ **FLOATING
C10181 XM2/a_100_139826# VSUBS 0.576721f $ **FLOATING
C10182 XM2/a_n158_139826# VSUBS 0.576721f $ **FLOATING
C10183 XM2/a_n100_139729# VSUBS 0.247431f $ **FLOATING
C10184 XM2/a_100_142462# VSUBS 0.576721f $ **FLOATING
C10185 XM2/a_n158_142462# VSUBS 0.576721f $ **FLOATING
C10186 XM2/a_n100_142365# VSUBS 0.247431f $ **FLOATING
C10187 XM2/a_100_145098# VSUBS 0.576721f $ **FLOATING
C10188 XM2/a_n158_145098# VSUBS 0.576721f $ **FLOATING
C10189 XM2/a_n100_145001# VSUBS 0.247431f $ **FLOATING
C10190 XM2/a_100_147734# VSUBS 0.576721f $ **FLOATING
C10191 XM2/a_n158_147734# VSUBS 0.576721f $ **FLOATING
C10192 XM2/a_n100_147637# VSUBS 0.247431f $ **FLOATING
C10193 XM2/a_100_150370# VSUBS 0.576721f $ **FLOATING
C10194 XM2/a_n158_150370# VSUBS 0.576721f $ **FLOATING
C10195 XM2/a_n100_150273# VSUBS 0.247431f $ **FLOATING
C10196 XM2/a_100_153006# VSUBS 0.576721f $ **FLOATING
C10197 XM2/a_n158_153006# VSUBS 0.576721f $ **FLOATING
C10198 XM2/a_n100_152909# VSUBS 0.247431f $ **FLOATING
C10199 XM2/a_100_155642# VSUBS 0.576721f $ **FLOATING
C10200 XM2/a_n158_155642# VSUBS 0.576721f $ **FLOATING
C10201 XM2/a_n100_155545# VSUBS 0.247431f $ **FLOATING
C10202 XM2/a_100_158278# VSUBS 0.576721f $ **FLOATING
C10203 XM2/a_n158_158278# VSUBS 0.576721f $ **FLOATING
C10204 XM2/a_n100_158181# VSUBS 0.247431f $ **FLOATING
C10205 XM2/a_100_160914# VSUBS 0.576721f $ **FLOATING
C10206 XM2/a_n158_160914# VSUBS 0.576721f $ **FLOATING
C10207 XM2/a_n100_160817# VSUBS 0.247431f $ **FLOATING
C10208 XM2/a_100_163550# VSUBS 0.576721f $ **FLOATING
C10209 XM2/a_n158_163550# VSUBS 0.576721f $ **FLOATING
C10210 XM2/a_n100_163453# VSUBS 0.247431f $ **FLOATING
C10211 XM2/a_100_166186# VSUBS 0.576721f $ **FLOATING
C10212 XM2/a_n158_166186# VSUBS 0.576721f $ **FLOATING
C10213 XM2/a_n100_166089# VSUBS 0.247431f $ **FLOATING
C10214 XM2/a_100_168822# VSUBS 0.576721f $ **FLOATING
C10215 XM2/a_n158_168822# VSUBS 0.576721f $ **FLOATING
C10216 XM2/a_n100_168725# VSUBS 0.247431f $ **FLOATING
C10217 XM2/a_100_171458# VSUBS 0.576721f $ **FLOATING
C10218 XM2/a_n158_171458# VSUBS 0.576721f $ **FLOATING
C10219 XM2/a_n100_171361# VSUBS 0.247431f $ **FLOATING
C10220 XM2/a_100_174094# VSUBS 0.576721f $ **FLOATING
C10221 XM2/a_n158_174094# VSUBS 0.576721f $ **FLOATING
C10222 XM2/a_n100_173997# VSUBS 0.247431f $ **FLOATING
C10223 XM2/a_100_176730# VSUBS 0.576721f $ **FLOATING
C10224 XM2/a_n158_176730# VSUBS 0.576721f $ **FLOATING
C10225 XM2/a_n100_176633# VSUBS 0.247431f $ **FLOATING
C10226 XM2/a_100_179366# VSUBS 0.576721f $ **FLOATING
C10227 XM2/a_n158_179366# VSUBS 0.576721f $ **FLOATING
C10228 XM2/a_n100_179269# VSUBS 0.247431f $ **FLOATING
C10229 XM2/a_100_182002# VSUBS 0.576721f $ **FLOATING
C10230 XM2/a_n158_182002# VSUBS 0.576721f $ **FLOATING
C10231 XM2/a_n100_181905# VSUBS 0.247431f $ **FLOATING
C10232 XM2/a_100_184638# VSUBS 0.576721f $ **FLOATING
C10233 XM2/a_n158_184638# VSUBS 0.576721f $ **FLOATING
C10234 XM2/a_n100_184541# VSUBS 0.247431f $ **FLOATING
C10235 XM2/a_100_187274# VSUBS 0.576721f $ **FLOATING
C10236 XM2/a_n158_187274# VSUBS 0.576721f $ **FLOATING
C10237 XM2/a_n100_187177# VSUBS 0.247431f $ **FLOATING
C10238 XM2/a_100_189910# VSUBS 0.576721f $ **FLOATING
C10239 XM2/a_n158_189910# VSUBS 0.576721f $ **FLOATING
C10240 XM2/a_n100_189813# VSUBS 0.247431f $ **FLOATING
C10241 XM2/a_100_192546# VSUBS 0.576721f $ **FLOATING
C10242 XM2/a_n158_192546# VSUBS 0.576721f $ **FLOATING
C10243 XM2/a_n100_192449# VSUBS 0.247431f $ **FLOATING
C10244 XM2/a_100_195182# VSUBS 0.576721f $ **FLOATING
C10245 XM2/a_n158_195182# VSUBS 0.576721f $ **FLOATING
C10246 XM2/a_n100_195085# VSUBS 0.247431f $ **FLOATING
C10247 XM2/a_100_197818# VSUBS 0.576721f $ **FLOATING
C10248 XM2/a_n158_197818# VSUBS 0.576721f $ **FLOATING
C10249 XM2/a_n100_197721# VSUBS 0.247431f $ **FLOATING
C10250 XM2/a_100_200454# VSUBS 0.576721f $ **FLOATING
C10251 XM2/a_n158_200454# VSUBS 0.576721f $ **FLOATING
C10252 XM2/a_n100_200357# VSUBS 0.247431f $ **FLOATING
C10253 XM2/a_100_203090# VSUBS 0.576721f $ **FLOATING
C10254 XM2/a_n158_203090# VSUBS 0.576721f $ **FLOATING
C10255 XM2/a_n100_202993# VSUBS 0.247431f $ **FLOATING
C10256 XM2/a_100_205726# VSUBS 0.576721f $ **FLOATING
C10257 XM2/a_n158_205726# VSUBS 0.576721f $ **FLOATING
C10258 XM2/a_n100_205629# VSUBS 0.247431f $ **FLOATING
C10259 XM2/a_100_208362# VSUBS 0.576721f $ **FLOATING
C10260 XM2/a_n158_208362# VSUBS 0.576721f $ **FLOATING
C10261 XM2/a_n100_208265# VSUBS 0.247431f $ **FLOATING
C10262 XM2/a_100_210998# VSUBS 0.576721f $ **FLOATING
C10263 XM2/a_n158_210998# VSUBS 0.576721f $ **FLOATING
C10264 XM2/a_n100_210901# VSUBS 0.247431f $ **FLOATING
C10265 XM2/a_100_213634# VSUBS 0.576721f $ **FLOATING
C10266 XM2/a_n158_213634# VSUBS 0.576721f $ **FLOATING
C10267 XM2/a_n100_213537# VSUBS 0.247431f $ **FLOATING
C10268 XM2/a_100_216270# VSUBS 0.576721f $ **FLOATING
C10269 XM2/a_n158_216270# VSUBS 0.576721f $ **FLOATING
C10270 XM2/a_n100_216173# VSUBS 0.247431f $ **FLOATING
C10271 XM2/a_100_218906# VSUBS 0.576721f $ **FLOATING
C10272 XM2/a_n158_218906# VSUBS 0.576721f $ **FLOATING
C10273 XM2/a_n100_218809# VSUBS 0.247431f $ **FLOATING
C10274 XM2/a_100_221542# VSUBS 0.576721f $ **FLOATING
C10275 XM2/a_n158_221542# VSUBS 0.576721f $ **FLOATING
C10276 XM2/a_n100_221445# VSUBS 0.247431f $ **FLOATING
C10277 XM2/a_100_224178# VSUBS 0.576721f $ **FLOATING
C10278 XM2/a_n158_224178# VSUBS 0.576721f $ **FLOATING
C10279 XM2/a_n100_224081# VSUBS 0.247431f $ **FLOATING
C10280 XM2/a_100_226814# VSUBS 0.576721f $ **FLOATING
C10281 XM2/a_n158_226814# VSUBS 0.576721f $ **FLOATING
C10282 XM2/a_n100_226717# VSUBS 0.247431f $ **FLOATING
C10283 XM2/a_100_229450# VSUBS 0.576721f $ **FLOATING
C10284 XM2/a_n158_229450# VSUBS 0.576721f $ **FLOATING
C10285 XM2/a_n100_229353# VSUBS 0.247431f $ **FLOATING
C10286 XM2/a_100_232086# VSUBS 0.576721f $ **FLOATING
C10287 XM2/a_n158_232086# VSUBS 0.576721f $ **FLOATING
C10288 XM2/a_n100_231989# VSUBS 0.247431f $ **FLOATING
C10289 XM2/a_100_234722# VSUBS 0.576721f $ **FLOATING
C10290 XM2/a_n158_234722# VSUBS 0.576721f $ **FLOATING
C10291 XM2/a_n100_234625# VSUBS 0.247431f $ **FLOATING
C10292 XM2/a_100_237358# VSUBS 0.576721f $ **FLOATING
C10293 XM2/a_n158_237358# VSUBS 0.576721f $ **FLOATING
C10294 XM2/a_n100_237261# VSUBS 0.247431f $ **FLOATING
C10295 XM2/a_100_239994# VSUBS 0.576721f $ **FLOATING
C10296 XM2/a_n158_239994# VSUBS 0.576721f $ **FLOATING
C10297 XM2/a_n100_239897# VSUBS 0.247431f $ **FLOATING
C10298 XM2/a_100_242630# VSUBS 0.576721f $ **FLOATING
C10299 XM2/a_n158_242630# VSUBS 0.576721f $ **FLOATING
C10300 XM2/a_n100_242533# VSUBS 0.247431f $ **FLOATING
C10301 XM2/a_100_245266# VSUBS 0.576721f $ **FLOATING
C10302 XM2/a_n158_245266# VSUBS 0.576721f $ **FLOATING
C10303 XM2/a_n100_245169# VSUBS 0.247431f $ **FLOATING
C10304 XM2/a_100_247902# VSUBS 0.576721f $ **FLOATING
C10305 XM2/a_n158_247902# VSUBS 0.576721f $ **FLOATING
C10306 XM2/a_n100_247805# VSUBS 0.247431f $ **FLOATING
C10307 XM2/a_100_250538# VSUBS 0.576721f $ **FLOATING
C10308 XM2/a_n158_250538# VSUBS 0.576721f $ **FLOATING
C10309 XM2/a_n100_250441# VSUBS 0.247431f $ **FLOATING
C10310 XM2/a_100_253174# VSUBS 0.576721f $ **FLOATING
C10311 XM2/a_n158_253174# VSUBS 0.576721f $ **FLOATING
C10312 XM2/a_n100_253077# VSUBS 0.247431f $ **FLOATING
C10313 XM2/a_100_255810# VSUBS 0.576721f $ **FLOATING
C10314 XM2/a_n158_255810# VSUBS 0.576721f $ **FLOATING
C10315 XM2/a_n100_255713# VSUBS 0.247431f $ **FLOATING
C10316 XM2/a_100_258446# VSUBS 0.576721f $ **FLOATING
C10317 XM2/a_n158_258446# VSUBS 0.576721f $ **FLOATING
C10318 XM2/a_n100_258349# VSUBS 0.247431f $ **FLOATING
C10319 XM2/a_100_261082# VSUBS 0.576721f $ **FLOATING
C10320 XM2/a_n158_261082# VSUBS 0.576721f $ **FLOATING
C10321 XM2/a_n100_260985# VSUBS 0.247431f $ **FLOATING
C10322 XM2/a_100_263718# VSUBS 0.576721f $ **FLOATING
C10323 XM2/a_n158_263718# VSUBS 0.576721f $ **FLOATING
C10324 XM2/a_n100_263621# VSUBS 0.247431f $ **FLOATING
C10325 XM2/a_100_266354# VSUBS 0.576721f $ **FLOATING
C10326 XM2/a_n158_266354# VSUBS 0.576721f $ **FLOATING
C10327 XM2/a_n100_266257# VSUBS 0.247431f $ **FLOATING
C10328 XM2/a_100_268990# VSUBS 0.576721f $ **FLOATING
C10329 XM2/a_n158_268990# VSUBS 0.576721f $ **FLOATING
C10330 XM2/a_n100_268893# VSUBS 0.247431f $ **FLOATING
C10331 XM2/a_100_271626# VSUBS 0.576721f $ **FLOATING
C10332 XM2/a_n158_271626# VSUBS 0.576721f $ **FLOATING
C10333 XM2/a_n100_271529# VSUBS 0.247431f $ **FLOATING
C10334 XM2/a_100_274262# VSUBS 0.576721f $ **FLOATING
C10335 XM2/a_n158_274262# VSUBS 0.576721f $ **FLOATING
C10336 XM2/a_n100_274165# VSUBS 0.247431f $ **FLOATING
C10337 XM2/a_100_276898# VSUBS 0.576721f $ **FLOATING
C10338 XM2/a_n158_276898# VSUBS 0.576721f $ **FLOATING
C10339 XM2/a_n100_276801# VSUBS 0.247431f $ **FLOATING
C10340 XM2/a_100_279534# VSUBS 0.576721f $ **FLOATING
C10341 XM2/a_n158_279534# VSUBS 0.576721f $ **FLOATING
C10342 XM2/a_n100_279437# VSUBS 0.247431f $ **FLOATING
C10343 XM2/a_100_282170# VSUBS 0.576721f $ **FLOATING
C10344 XM2/a_n158_282170# VSUBS 0.576721f $ **FLOATING
C10345 XM2/a_n100_282073# VSUBS 0.247431f $ **FLOATING
C10346 XM2/a_100_284806# VSUBS 0.576721f $ **FLOATING
C10347 XM2/a_n158_284806# VSUBS 0.576721f $ **FLOATING
C10348 XM2/a_n100_284709# VSUBS 0.247431f $ **FLOATING
C10349 XM2/a_100_287442# VSUBS 0.576721f $ **FLOATING
C10350 XM2/a_n158_287442# VSUBS 0.576721f $ **FLOATING
C10351 XM2/a_n100_287345# VSUBS 0.247431f $ **FLOATING
C10352 XM2/a_100_290078# VSUBS 0.576721f $ **FLOATING
C10353 XM2/a_n158_290078# VSUBS 0.576721f $ **FLOATING
C10354 XM2/a_n100_289981# VSUBS 0.247431f $ **FLOATING
C10355 XM2/a_100_292714# VSUBS 0.576721f $ **FLOATING
C10356 XM2/a_n158_292714# VSUBS 0.576721f $ **FLOATING
C10357 XM2/a_n100_292617# VSUBS 0.247431f $ **FLOATING
C10358 XM2/a_100_295350# VSUBS 0.576721f $ **FLOATING
C10359 XM2/a_n158_295350# VSUBS 0.576721f $ **FLOATING
C10360 XM2/a_n100_295253# VSUBS 0.247431f $ **FLOATING
C10361 XM2/a_100_297986# VSUBS 0.576721f $ **FLOATING
C10362 XM2/a_n158_297986# VSUBS 0.576721f $ **FLOATING
C10363 XM2/a_n100_297889# VSUBS 0.247431f $ **FLOATING
C10364 XM2/a_100_300622# VSUBS 0.576721f $ **FLOATING
C10365 XM2/a_n158_300622# VSUBS 0.576721f $ **FLOATING
C10366 XM2/a_n100_300525# VSUBS 0.247431f $ **FLOATING
C10367 XM2/a_100_303258# VSUBS 0.576721f $ **FLOATING
C10368 XM2/a_n158_303258# VSUBS 0.576721f $ **FLOATING
C10369 XM2/a_n100_303161# VSUBS 0.247431f $ **FLOATING
C10370 XM2/a_100_305894# VSUBS 0.576721f $ **FLOATING
C10371 XM2/a_n158_305894# VSUBS 0.576721f $ **FLOATING
C10372 XM2/a_n100_305797# VSUBS 0.247431f $ **FLOATING
C10373 XM2/a_100_308530# VSUBS 0.576721f $ **FLOATING
C10374 XM2/a_n158_308530# VSUBS 0.576721f $ **FLOATING
C10375 XM2/a_n100_308433# VSUBS 0.247431f $ **FLOATING
C10376 XM2/a_100_311166# VSUBS 0.576721f $ **FLOATING
C10377 XM2/a_n158_311166# VSUBS 0.576721f $ **FLOATING
C10378 XM2/a_n100_311069# VSUBS 0.247431f $ **FLOATING
C10379 XM2/a_100_313802# VSUBS 0.576721f $ **FLOATING
C10380 XM2/a_n158_313802# VSUBS 0.576721f $ **FLOATING
C10381 XM2/a_n100_313705# VSUBS 0.247431f $ **FLOATING
C10382 XM2/a_100_316438# VSUBS 0.576721f $ **FLOATING
C10383 XM2/a_n158_316438# VSUBS 0.576721f $ **FLOATING
C10384 XM2/a_n100_316341# VSUBS 0.247431f $ **FLOATING
C10385 XM2/a_100_319074# VSUBS 0.576721f $ **FLOATING
C10386 XM2/a_n158_319074# VSUBS 0.576721f $ **FLOATING
C10387 XM2/a_n100_318977# VSUBS 0.247431f $ **FLOATING
C10388 XM2/a_100_321710# VSUBS 0.576721f $ **FLOATING
C10389 XM2/a_n158_321710# VSUBS 0.576721f $ **FLOATING
C10390 XM2/a_n100_321613# VSUBS 0.247431f $ **FLOATING
C10391 XM2/a_100_324346# VSUBS 0.576721f $ **FLOATING
C10392 XM2/a_n158_324346# VSUBS 0.576721f $ **FLOATING
C10393 XM2/a_n100_324249# VSUBS 0.247431f $ **FLOATING
C10394 XM2/a_100_326982# VSUBS 0.576721f $ **FLOATING
C10395 XM2/a_n158_326982# VSUBS 0.576721f $ **FLOATING
C10396 XM2/a_n100_326885# VSUBS 0.247431f $ **FLOATING
C10397 XM2/a_100_329618# VSUBS 0.576721f $ **FLOATING
C10398 XM2/a_n158_329618# VSUBS 0.576721f $ **FLOATING
C10399 XM2/a_n100_329521# VSUBS 0.247431f $ **FLOATING
C10400 XM2/a_100_332254# VSUBS 0.576721f $ **FLOATING
C10401 XM2/a_n158_332254# VSUBS 0.576721f $ **FLOATING
C10402 XM2/a_n100_332157# VSUBS 0.247431f $ **FLOATING
C10403 XM2/a_100_334890# VSUBS 0.58217f $ **FLOATING
C10404 XM2/a_n158_334890# VSUBS 0.58217f $ **FLOATING
C10405 XM2/a_n100_334793# VSUBS 0.291162f $ **FLOATING
C10406 XM4/w_n358_n132787# VSUBS 4.196118p
C10407 XM1/a_100_n183690# VSUBS 0.292592f
C10408 XM1/a_n158_n183690# VSUBS 0.292592f
C10409 XM1/a_n100_n183787# VSUBS 0.265338f
C10410 XM1/a_100_n182254# VSUBS 0.287142f
C10411 XM1/a_n158_n182254# VSUBS 0.287142f
C10412 XM1/a_n100_n182351# VSUBS 0.221608f
C10413 XM1/a_100_n180818# VSUBS 0.287142f
C10414 XM1/a_n158_n180818# VSUBS 0.287142f
C10415 XM1/a_n100_n180915# VSUBS 0.221608f
C10416 XM1/a_100_n179382# VSUBS 0.287142f
C10417 XM1/a_n158_n179382# VSUBS 0.287142f
C10418 XM1/a_n100_n179479# VSUBS 0.221608f
C10419 XM1/a_100_n177946# VSUBS 0.287142f
C10420 XM1/a_n158_n177946# VSUBS 0.287142f
C10421 XM1/a_n100_n178043# VSUBS 0.221608f
C10422 XM1/a_100_n176510# VSUBS 0.287142f
C10423 XM1/a_n158_n176510# VSUBS 0.287142f
C10424 XM1/a_n100_n176607# VSUBS 0.221608f
C10425 XM1/a_100_n175074# VSUBS 0.287142f
C10426 XM1/a_n158_n175074# VSUBS 0.287142f
C10427 XM1/a_n100_n175171# VSUBS 0.221608f
C10428 XM1/a_100_n173638# VSUBS 0.287142f
C10429 XM1/a_n158_n173638# VSUBS 0.287142f
C10430 XM1/a_n100_n173735# VSUBS 0.221608f
C10431 XM1/a_100_n172202# VSUBS 0.287142f
C10432 XM1/a_n158_n172202# VSUBS 0.287142f
C10433 XM1/a_n100_n172299# VSUBS 0.221608f
C10434 XM1/a_100_n170766# VSUBS 0.287142f
C10435 XM1/a_n158_n170766# VSUBS 0.287142f
C10436 XM1/a_n100_n170863# VSUBS 0.221608f
C10437 XM1/a_100_n169330# VSUBS 0.287142f
C10438 XM1/a_n158_n169330# VSUBS 0.287142f
C10439 XM1/a_n100_n169427# VSUBS 0.221608f
C10440 XM1/a_100_n167894# VSUBS 0.287142f
C10441 XM1/a_n158_n167894# VSUBS 0.287142f
C10442 XM1/a_n100_n167991# VSUBS 0.221608f
C10443 XM1/a_100_n166458# VSUBS 0.287142f
C10444 XM1/a_n158_n166458# VSUBS 0.287142f
C10445 XM1/a_n100_n166555# VSUBS 0.221608f
C10446 XM1/a_100_n165022# VSUBS 0.287142f
C10447 XM1/a_n158_n165022# VSUBS 0.287142f
C10448 XM1/a_n100_n165119# VSUBS 0.221608f
C10449 XM1/a_100_n163586# VSUBS 0.287142f
C10450 XM1/a_n158_n163586# VSUBS 0.287142f
C10451 XM1/a_n100_n163683# VSUBS 0.221608f
C10452 XM1/a_100_n162150# VSUBS 0.287142f
C10453 XM1/a_n158_n162150# VSUBS 0.287142f
C10454 XM1/a_n100_n162247# VSUBS 0.221608f
C10455 XM1/a_100_n160714# VSUBS 0.287142f
C10456 XM1/a_n158_n160714# VSUBS 0.287142f
C10457 XM1/a_n100_n160811# VSUBS 0.221608f
C10458 XM1/a_100_n159278# VSUBS 0.287142f
C10459 XM1/a_n158_n159278# VSUBS 0.287142f
C10460 XM1/a_n100_n159375# VSUBS 0.221608f
C10461 XM1/a_100_n157842# VSUBS 0.287142f
C10462 XM1/a_n158_n157842# VSUBS 0.287142f
C10463 XM1/a_n100_n157939# VSUBS 0.221608f
C10464 XM1/a_100_n156406# VSUBS 0.287142f
C10465 XM1/a_n158_n156406# VSUBS 0.287142f
C10466 XM1/a_n100_n156503# VSUBS 0.221608f
C10467 XM1/a_100_n154970# VSUBS 0.287142f
C10468 XM1/a_n158_n154970# VSUBS 0.287142f
C10469 XM1/a_n100_n155067# VSUBS 0.221608f
C10470 XM1/a_100_n153534# VSUBS 0.287142f
C10471 XM1/a_n158_n153534# VSUBS 0.287142f
C10472 XM1/a_n100_n153631# VSUBS 0.221608f
C10473 XM1/a_100_n152098# VSUBS 0.287142f
C10474 XM1/a_n158_n152098# VSUBS 0.287142f
C10475 XM1/a_n100_n152195# VSUBS 0.221608f
C10476 XM1/a_100_n150662# VSUBS 0.287142f
C10477 XM1/a_n158_n150662# VSUBS 0.287142f
C10478 XM1/a_n100_n150759# VSUBS 0.221608f
C10479 XM1/a_100_n149226# VSUBS 0.287142f
C10480 XM1/a_n158_n149226# VSUBS 0.287142f
C10481 XM1/a_n100_n149323# VSUBS 0.221608f
C10482 XM1/a_100_n147790# VSUBS 0.287142f
C10483 XM1/a_n158_n147790# VSUBS 0.287142f
C10484 XM1/a_n100_n147887# VSUBS 0.221608f
C10485 XM1/a_100_n146354# VSUBS 0.287142f
C10486 XM1/a_n158_n146354# VSUBS 0.287142f
C10487 XM1/a_n100_n146451# VSUBS 0.221608f
C10488 XM1/a_100_n144918# VSUBS 0.287142f
C10489 XM1/a_n158_n144918# VSUBS 0.287142f
C10490 XM1/a_n100_n145015# VSUBS 0.221608f
C10491 XM1/a_100_n143482# VSUBS 0.287142f
C10492 XM1/a_n158_n143482# VSUBS 0.287142f
C10493 XM1/a_n100_n143579# VSUBS 0.221608f
C10494 XM1/a_100_n142046# VSUBS 0.287142f
C10495 XM1/a_n158_n142046# VSUBS 0.287142f
C10496 XM1/a_n100_n142143# VSUBS 0.221608f
C10497 XM1/a_100_n140610# VSUBS 0.287142f
C10498 XM1/a_n158_n140610# VSUBS 0.287142f
C10499 XM1/a_n100_n140707# VSUBS 0.221608f
C10500 XM1/a_100_n139174# VSUBS 0.287142f
C10501 XM1/a_n158_n139174# VSUBS 0.287142f
C10502 XM1/a_n100_n139271# VSUBS 0.221608f
C10503 XM1/a_100_n137738# VSUBS 0.287142f
C10504 XM1/a_n158_n137738# VSUBS 0.287142f
C10505 XM1/a_n100_n137835# VSUBS 0.221608f
C10506 XM1/a_100_n136302# VSUBS 0.287142f
C10507 XM1/a_n158_n136302# VSUBS 0.287142f
C10508 XM1/a_n100_n136399# VSUBS 0.221608f
C10509 XM1/a_100_n134866# VSUBS 0.287142f
C10510 XM1/a_n158_n134866# VSUBS 0.287142f
C10511 XM1/a_n100_n134963# VSUBS 0.221608f
C10512 XM1/a_100_n133430# VSUBS 0.287142f
C10513 XM1/a_n158_n133430# VSUBS 0.287142f
C10514 XM1/a_n100_n133527# VSUBS 0.221608f
C10515 XM1/a_100_n131994# VSUBS 0.287142f
C10516 XM1/a_n158_n131994# VSUBS 0.287142f
C10517 XM1/a_n100_n132091# VSUBS 0.221608f
C10518 XM1/a_100_n130558# VSUBS 0.287142f
C10519 XM1/a_n158_n130558# VSUBS 0.287142f
C10520 XM1/a_n100_n130655# VSUBS 0.221608f
C10521 XM1/a_100_n129122# VSUBS 0.287142f
C10522 XM1/a_n158_n129122# VSUBS 0.287142f
C10523 XM1/a_n100_n129219# VSUBS 0.221608f
C10524 XM1/a_100_n127686# VSUBS 0.287142f
C10525 XM1/a_n158_n127686# VSUBS 0.287142f
C10526 XM1/a_n100_n127783# VSUBS 0.221608f
C10527 XM1/a_100_n126250# VSUBS 0.287142f
C10528 XM1/a_n158_n126250# VSUBS 0.287142f
C10529 XM1/a_n100_n126347# VSUBS 0.221608f
C10530 XM1/a_100_n124814# VSUBS 0.287142f
C10531 XM1/a_n158_n124814# VSUBS 0.287142f
C10532 XM1/a_n100_n124911# VSUBS 0.221608f
C10533 XM1/a_100_n123378# VSUBS 0.287142f
C10534 XM1/a_n158_n123378# VSUBS 0.287142f
C10535 XM1/a_n100_n123475# VSUBS 0.221608f
C10536 XM1/a_100_n121942# VSUBS 0.287142f
C10537 XM1/a_n158_n121942# VSUBS 0.287142f
C10538 XM1/a_n100_n122039# VSUBS 0.221608f
C10539 XM1/a_100_n120506# VSUBS 0.287142f
C10540 XM1/a_n158_n120506# VSUBS 0.287142f
C10541 XM1/a_n100_n120603# VSUBS 0.221608f
C10542 XM1/a_100_n119070# VSUBS 0.287142f
C10543 XM1/a_n158_n119070# VSUBS 0.287142f
C10544 XM1/a_n100_n119167# VSUBS 0.221608f
C10545 XM1/a_100_n117634# VSUBS 0.287142f
C10546 XM1/a_n158_n117634# VSUBS 0.287142f
C10547 XM1/a_n100_n117731# VSUBS 0.221608f
C10548 XM1/a_100_n116198# VSUBS 0.287142f
C10549 XM1/a_n158_n116198# VSUBS 0.287142f
C10550 XM1/a_n100_n116295# VSUBS 0.221608f
C10551 XM1/a_100_n114762# VSUBS 0.287142f
C10552 XM1/a_n158_n114762# VSUBS 0.287142f
C10553 XM1/a_n100_n114859# VSUBS 0.221608f
C10554 XM1/a_100_n113326# VSUBS 0.287142f
C10555 XM1/a_n158_n113326# VSUBS 0.287142f
C10556 XM1/a_n100_n113423# VSUBS 0.221608f
C10557 XM1/a_100_n111890# VSUBS 0.287142f
C10558 XM1/a_n158_n111890# VSUBS 0.287142f
C10559 XM1/a_n100_n111987# VSUBS 0.221608f
C10560 XM1/a_100_n110454# VSUBS 0.287142f
C10561 XM1/a_n158_n110454# VSUBS 0.287142f
C10562 XM1/a_n100_n110551# VSUBS 0.221608f
C10563 XM1/a_100_n109018# VSUBS 0.287142f
C10564 XM1/a_n158_n109018# VSUBS 0.287142f
C10565 XM1/a_n100_n109115# VSUBS 0.221608f
C10566 XM1/a_100_n107582# VSUBS 0.287142f
C10567 XM1/a_n158_n107582# VSUBS 0.287142f
C10568 XM1/a_n100_n107679# VSUBS 0.221608f
C10569 XM1/a_100_n106146# VSUBS 0.287142f
C10570 XM1/a_n158_n106146# VSUBS 0.287142f
C10571 XM1/a_n100_n106243# VSUBS 0.221608f
C10572 XM1/a_100_n104710# VSUBS 0.287142f
C10573 XM1/a_n158_n104710# VSUBS 0.287142f
C10574 XM1/a_n100_n104807# VSUBS 0.221608f
C10575 XM1/a_100_n103274# VSUBS 0.287142f
C10576 XM1/a_n158_n103274# VSUBS 0.287142f
C10577 XM1/a_n100_n103371# VSUBS 0.221608f
C10578 XM1/a_100_n101838# VSUBS 0.287142f
C10579 XM1/a_n158_n101838# VSUBS 0.287142f
C10580 XM1/a_n100_n101935# VSUBS 0.221608f
C10581 XM1/a_100_n100402# VSUBS 0.287142f
C10582 XM1/a_n158_n100402# VSUBS 0.287142f
C10583 XM1/a_n100_n100499# VSUBS 0.221608f
C10584 XM1/a_100_n98966# VSUBS 0.287142f
C10585 XM1/a_n158_n98966# VSUBS 0.287142f
C10586 XM1/a_n100_n99063# VSUBS 0.221608f
C10587 XM1/a_100_n97530# VSUBS 0.287142f
C10588 XM1/a_n158_n97530# VSUBS 0.287142f
C10589 XM1/a_n100_n97627# VSUBS 0.221608f
C10590 XM1/a_100_n96094# VSUBS 0.287142f
C10591 XM1/a_n158_n96094# VSUBS 0.287142f
C10592 XM1/a_n100_n96191# VSUBS 0.221608f
C10593 XM1/a_100_n94658# VSUBS 0.287142f
C10594 XM1/a_n158_n94658# VSUBS 0.287142f
C10595 XM1/a_n100_n94755# VSUBS 0.221608f
C10596 XM1/a_100_n93222# VSUBS 0.287142f
C10597 XM1/a_n158_n93222# VSUBS 0.287142f
C10598 XM1/a_n100_n93319# VSUBS 0.221608f
C10599 XM1/a_100_n91786# VSUBS 0.287142f
C10600 XM1/a_n158_n91786# VSUBS 0.287142f
C10601 XM1/a_n100_n91883# VSUBS 0.221608f
C10602 XM1/a_100_n90350# VSUBS 0.287142f
C10603 XM1/a_n158_n90350# VSUBS 0.287142f
C10604 XM1/a_n100_n90447# VSUBS 0.221608f
C10605 XM1/a_100_n88914# VSUBS 0.287142f
C10606 XM1/a_n158_n88914# VSUBS 0.287142f
C10607 XM1/a_n100_n89011# VSUBS 0.221608f
C10608 XM1/a_100_n87478# VSUBS 0.287142f
C10609 XM1/a_n158_n87478# VSUBS 0.287142f
C10610 XM1/a_n100_n87575# VSUBS 0.221608f
C10611 XM1/a_100_n86042# VSUBS 0.287142f
C10612 XM1/a_n158_n86042# VSUBS 0.287142f
C10613 XM1/a_n100_n86139# VSUBS 0.221608f
C10614 XM1/a_100_n84606# VSUBS 0.287142f
C10615 XM1/a_n158_n84606# VSUBS 0.287142f
C10616 XM1/a_n100_n84703# VSUBS 0.221608f
C10617 XM1/a_100_n83170# VSUBS 0.287142f
C10618 XM1/a_n158_n83170# VSUBS 0.287142f
C10619 XM1/a_n100_n83267# VSUBS 0.221608f
C10620 XM1/a_100_n81734# VSUBS 0.287142f
C10621 XM1/a_n158_n81734# VSUBS 0.287142f
C10622 XM1/a_n100_n81831# VSUBS 0.221608f
C10623 XM1/a_100_n80298# VSUBS 0.287142f
C10624 XM1/a_n158_n80298# VSUBS 0.287142f
C10625 XM1/a_n100_n80395# VSUBS 0.221608f
C10626 XM1/a_100_n78862# VSUBS 0.287142f
C10627 XM1/a_n158_n78862# VSUBS 0.287142f
C10628 XM1/a_n100_n78959# VSUBS 0.221608f
C10629 XM1/a_100_n77426# VSUBS 0.287142f
C10630 XM1/a_n158_n77426# VSUBS 0.287142f
C10631 XM1/a_n100_n77523# VSUBS 0.221608f
C10632 XM1/a_100_n75990# VSUBS 0.287142f
C10633 XM1/a_n158_n75990# VSUBS 0.287142f
C10634 XM1/a_n100_n76087# VSUBS 0.221608f
C10635 XM1/a_100_n74554# VSUBS 0.287142f
C10636 XM1/a_n158_n74554# VSUBS 0.287142f
C10637 XM1/a_n100_n74651# VSUBS 0.221608f
C10638 XM1/a_100_n73118# VSUBS 0.287142f
C10639 XM1/a_n158_n73118# VSUBS 0.287142f
C10640 XM1/a_n100_n73215# VSUBS 0.221608f
C10641 XM1/a_100_n71682# VSUBS 0.287142f
C10642 XM1/a_n158_n71682# VSUBS 0.287142f
C10643 XM1/a_n100_n71779# VSUBS 0.221608f
C10644 XM1/a_100_n70246# VSUBS 0.287142f
C10645 XM1/a_n158_n70246# VSUBS 0.287142f
C10646 XM1/a_n100_n70343# VSUBS 0.221608f
C10647 XM1/a_100_n68810# VSUBS 0.287142f
C10648 XM1/a_n158_n68810# VSUBS 0.287142f
C10649 XM1/a_n100_n68907# VSUBS 0.221608f
C10650 XM1/a_100_n67374# VSUBS 0.287142f
C10651 XM1/a_n158_n67374# VSUBS 0.287142f
C10652 XM1/a_n100_n67471# VSUBS 0.221608f
C10653 XM1/a_100_n65938# VSUBS 0.287142f
C10654 XM1/a_n158_n65938# VSUBS 0.287142f
C10655 XM1/a_n100_n66035# VSUBS 0.221608f
C10656 XM1/a_100_n64502# VSUBS 0.287142f
C10657 XM1/a_n158_n64502# VSUBS 0.287142f
C10658 XM1/a_n100_n64599# VSUBS 0.221608f
C10659 XM1/a_100_n63066# VSUBS 0.287142f
C10660 XM1/a_n158_n63066# VSUBS 0.287142f
C10661 XM1/a_n100_n63163# VSUBS 0.221608f
C10662 XM1/a_100_n61630# VSUBS 0.287142f
C10663 XM1/a_n158_n61630# VSUBS 0.287142f
C10664 XM1/a_n100_n61727# VSUBS 0.221608f
C10665 XM1/a_100_n60194# VSUBS 0.287142f
C10666 XM1/a_n158_n60194# VSUBS 0.287142f
C10667 XM1/a_n100_n60291# VSUBS 0.221608f
C10668 XM1/a_100_n58758# VSUBS 0.287142f
C10669 XM1/a_n158_n58758# VSUBS 0.287142f
C10670 XM1/a_n100_n58855# VSUBS 0.221608f
C10671 XM1/a_100_n57322# VSUBS 0.287142f
C10672 XM1/a_n158_n57322# VSUBS 0.287142f
C10673 XM1/a_n100_n57419# VSUBS 0.221608f
C10674 XM1/a_100_n55886# VSUBS 0.287142f
C10675 XM1/a_n158_n55886# VSUBS 0.287142f
C10676 XM1/a_n100_n55983# VSUBS 0.221608f
C10677 XM1/a_100_n54450# VSUBS 0.287142f
C10678 XM1/a_n158_n54450# VSUBS 0.287142f
C10679 XM1/a_n100_n54547# VSUBS 0.221608f
C10680 XM1/a_100_n53014# VSUBS 0.287142f
C10681 XM1/a_n158_n53014# VSUBS 0.287142f
C10682 XM1/a_n100_n53111# VSUBS 0.221608f
C10683 XM1/a_100_n51578# VSUBS 0.287142f
C10684 XM1/a_n158_n51578# VSUBS 0.287142f
C10685 XM1/a_n100_n51675# VSUBS 0.221608f
C10686 XM1/a_100_n50142# VSUBS 0.287142f
C10687 XM1/a_n158_n50142# VSUBS 0.287142f
C10688 XM1/a_n100_n50239# VSUBS 0.221608f
C10689 XM1/a_100_n48706# VSUBS 0.287142f
C10690 XM1/a_n158_n48706# VSUBS 0.287142f
C10691 XM1/a_n100_n48803# VSUBS 0.221608f
C10692 XM1/a_100_n47270# VSUBS 0.287142f
C10693 XM1/a_n158_n47270# VSUBS 0.287142f
C10694 XM1/a_n100_n47367# VSUBS 0.221608f
C10695 XM1/a_100_n45834# VSUBS 0.287142f
C10696 XM1/a_n158_n45834# VSUBS 0.287142f
C10697 XM1/a_n100_n45931# VSUBS 0.221608f
C10698 XM1/a_100_n44398# VSUBS 0.287142f
C10699 XM1/a_n158_n44398# VSUBS 0.287142f
C10700 XM1/a_n100_n44495# VSUBS 0.221608f
C10701 XM1/a_100_n42962# VSUBS 0.287142f
C10702 XM1/a_n158_n42962# VSUBS 0.287142f
C10703 XM1/a_n100_n43059# VSUBS 0.221608f
C10704 XM1/a_100_n41526# VSUBS 0.287142f
C10705 XM1/a_n158_n41526# VSUBS 0.287142f
C10706 XM1/a_n100_n41623# VSUBS 0.221608f
C10707 XM1/a_100_n40090# VSUBS 0.287142f
C10708 XM1/a_n158_n40090# VSUBS 0.287142f
C10709 XM1/a_n100_n40187# VSUBS 0.221608f
C10710 XM1/a_100_n38654# VSUBS 0.287142f
C10711 XM1/a_n158_n38654# VSUBS 0.287142f
C10712 XM1/a_n100_n38751# VSUBS 0.221608f
C10713 XM1/a_100_n37218# VSUBS 0.287142f
C10714 XM1/a_n158_n37218# VSUBS 0.287142f
C10715 XM1/a_n100_n37315# VSUBS 0.221608f
C10716 XM1/a_100_n35782# VSUBS 0.287142f
C10717 XM1/a_n158_n35782# VSUBS 0.287142f
C10718 XM1/a_n100_n35879# VSUBS 0.221608f
C10719 XM1/a_100_n34346# VSUBS 0.287142f
C10720 XM1/a_n158_n34346# VSUBS 0.287142f
C10721 XM1/a_n100_n34443# VSUBS 0.221608f
C10722 XM1/a_100_n32910# VSUBS 0.287142f
C10723 XM1/a_n158_n32910# VSUBS 0.287142f
C10724 XM1/a_n100_n33007# VSUBS 0.221608f
C10725 XM1/a_100_n31474# VSUBS 0.287142f
C10726 XM1/a_n158_n31474# VSUBS 0.287142f
C10727 XM1/a_n100_n31571# VSUBS 0.221608f
C10728 XM1/a_100_n30038# VSUBS 0.287142f
C10729 XM1/a_n158_n30038# VSUBS 0.287142f
C10730 XM1/a_n100_n30135# VSUBS 0.221608f
C10731 XM1/a_100_n28602# VSUBS 0.287142f
C10732 XM1/a_n158_n28602# VSUBS 0.287142f
C10733 XM1/a_n100_n28699# VSUBS 0.221608f
C10734 XM1/a_100_n27166# VSUBS 0.287142f
C10735 XM1/a_n158_n27166# VSUBS 0.287142f
C10736 XM1/a_n100_n27263# VSUBS 0.221608f
C10737 XM1/a_100_n25730# VSUBS 0.287142f
C10738 XM1/a_n158_n25730# VSUBS 0.287142f
C10739 XM1/a_n100_n25827# VSUBS 0.221608f
C10740 XM1/a_100_n24294# VSUBS 0.287142f
C10741 XM1/a_n158_n24294# VSUBS 0.287142f
C10742 XM1/a_n100_n24391# VSUBS 0.221608f
C10743 XM1/a_100_n22858# VSUBS 0.287142f
C10744 XM1/a_n158_n22858# VSUBS 0.287142f
C10745 XM1/a_n100_n22955# VSUBS 0.221608f
C10746 XM1/a_100_n21422# VSUBS 0.287142f
C10747 XM1/a_n158_n21422# VSUBS 0.287142f
C10748 XM1/a_n100_n21519# VSUBS 0.221608f
C10749 XM1/a_100_n19986# VSUBS 0.287142f
C10750 XM1/a_n158_n19986# VSUBS 0.287142f
C10751 XM1/a_n100_n20083# VSUBS 0.221608f
C10752 XM1/a_100_n18550# VSUBS 0.287142f
C10753 XM1/a_n158_n18550# VSUBS 0.287142f
C10754 XM1/a_n100_n18647# VSUBS 0.221608f
C10755 XM1/a_100_n17114# VSUBS 0.287142f
C10756 XM1/a_n158_n17114# VSUBS 0.287142f
C10757 XM1/a_n100_n17211# VSUBS 0.221608f
C10758 XM1/a_100_n15678# VSUBS 0.287142f
C10759 XM1/a_n158_n15678# VSUBS 0.287142f
C10760 XM1/a_n100_n15775# VSUBS 0.221608f
C10761 XM1/a_100_n14242# VSUBS 0.287142f
C10762 XM1/a_n158_n14242# VSUBS 0.287142f
C10763 XM1/a_n100_n14339# VSUBS 0.221608f
C10764 XM1/a_100_n12806# VSUBS 0.287142f
C10765 XM1/a_n158_n12806# VSUBS 0.287142f
C10766 XM1/a_n100_n12903# VSUBS 0.221608f
C10767 XM1/a_100_n11370# VSUBS 0.287142f
C10768 XM1/a_n158_n11370# VSUBS 0.287142f
C10769 XM1/a_n100_n11467# VSUBS 0.221608f
C10770 XM1/a_100_n9934# VSUBS 0.287142f
C10771 XM1/a_n158_n9934# VSUBS 0.287142f
C10772 XM1/a_n100_n10031# VSUBS 0.221608f
C10773 XM1/a_100_n8498# VSUBS 0.287142f
C10774 XM1/a_n158_n8498# VSUBS 0.287142f
C10775 XM1/a_n100_n8595# VSUBS 0.221608f
C10776 XM1/a_100_n7062# VSUBS 0.287142f
C10777 XM1/a_n158_n7062# VSUBS 0.287142f
C10778 XM1/a_n100_n7159# VSUBS 0.221608f
C10779 XM1/a_100_n5626# VSUBS 0.287142f
C10780 XM1/a_n158_n5626# VSUBS 0.287142f
C10781 XM1/a_n100_n5723# VSUBS 0.221608f
C10782 XM1/a_100_n4190# VSUBS 0.287142f
C10783 XM1/a_n158_n4190# VSUBS 0.287142f
C10784 XM1/a_n100_n4287# VSUBS 0.221608f
C10785 XM1/a_100_n2754# VSUBS 0.287142f
C10786 XM1/a_n158_n2754# VSUBS 0.287142f
C10787 XM1/a_n100_n2851# VSUBS 0.221608f
C10788 XM1/a_100_n1318# VSUBS 0.287142f
C10789 XM1/a_n158_n1318# VSUBS 0.287142f
C10790 XM1/a_n100_n1415# VSUBS 0.221608f
C10791 XM1/a_100_118# VSUBS 0.287142f
C10792 XM1/a_n158_118# VSUBS 0.287142f
C10793 XM1/a_n100_21# VSUBS 0.221608f
C10794 XM1/a_100_1554# VSUBS 0.287142f
C10795 XM1/a_n158_1554# VSUBS 0.287142f
C10796 XM1/a_n100_1457# VSUBS 0.221608f
C10797 XM1/a_100_2990# VSUBS 0.287142f
C10798 XM1/a_n158_2990# VSUBS 0.287142f
C10799 XM1/a_n100_2893# VSUBS 0.221608f
C10800 XM1/a_100_4426# VSUBS 0.287142f
C10801 XM1/a_n158_4426# VSUBS 0.287142f
C10802 XM1/a_n100_4329# VSUBS 0.221608f
C10803 XM1/a_100_5862# VSUBS 0.287142f
C10804 XM1/a_n158_5862# VSUBS 0.287142f
C10805 XM1/a_n100_5765# VSUBS 0.221608f
C10806 XM1/a_100_7298# VSUBS 0.287142f
C10807 XM1/a_n158_7298# VSUBS 0.287142f
C10808 XM1/a_n100_7201# VSUBS 0.221608f
C10809 XM1/a_100_8734# VSUBS 0.287142f
C10810 XM1/a_n158_8734# VSUBS 0.287142f
C10811 XM1/a_n100_8637# VSUBS 0.221608f
C10812 XM1/a_100_10170# VSUBS 0.287142f
C10813 XM1/a_n158_10170# VSUBS 0.287142f
C10814 XM1/a_n100_10073# VSUBS 0.221608f
C10815 XM1/a_100_11606# VSUBS 0.287142f
C10816 XM1/a_n158_11606# VSUBS 0.287142f
C10817 XM1/a_n100_11509# VSUBS 0.221608f
C10818 XM1/a_100_13042# VSUBS 0.287142f
C10819 XM1/a_n158_13042# VSUBS 0.287142f
C10820 XM1/a_n100_12945# VSUBS 0.221608f
C10821 XM1/a_100_14478# VSUBS 0.287142f
C10822 XM1/a_n158_14478# VSUBS 0.287142f
C10823 XM1/a_n100_14381# VSUBS 0.221608f
C10824 XM1/a_100_15914# VSUBS 0.287142f
C10825 XM1/a_n158_15914# VSUBS 0.287142f
C10826 XM1/a_n100_15817# VSUBS 0.221608f
C10827 XM1/a_100_17350# VSUBS 0.287142f
C10828 XM1/a_n158_17350# VSUBS 0.287142f
C10829 XM1/a_n100_17253# VSUBS 0.221608f
C10830 XM1/a_100_18786# VSUBS 0.287142f
C10831 XM1/a_n158_18786# VSUBS 0.287142f
C10832 XM1/a_n100_18689# VSUBS 0.221608f
C10833 XM1/a_100_20222# VSUBS 0.287142f
C10834 XM1/a_n158_20222# VSUBS 0.287142f
C10835 XM1/a_n100_20125# VSUBS 0.221608f
C10836 XM1/a_100_21658# VSUBS 0.287142f
C10837 XM1/a_n158_21658# VSUBS 0.287142f
C10838 XM1/a_n100_21561# VSUBS 0.221608f
C10839 XM1/a_100_23094# VSUBS 0.287142f
C10840 XM1/a_n158_23094# VSUBS 0.287142f
C10841 XM1/a_n100_22997# VSUBS 0.221608f
C10842 XM1/a_100_24530# VSUBS 0.287142f
C10843 XM1/a_n158_24530# VSUBS 0.287142f
C10844 XM1/a_n100_24433# VSUBS 0.221608f
C10845 XM1/a_100_25966# VSUBS 0.287142f
C10846 XM1/a_n158_25966# VSUBS 0.287142f
C10847 XM1/a_n100_25869# VSUBS 0.221608f
C10848 XM1/a_100_27402# VSUBS 0.287142f
C10849 XM1/a_n158_27402# VSUBS 0.287142f
C10850 XM1/a_n100_27305# VSUBS 0.221608f
C10851 XM1/a_100_28838# VSUBS 0.287142f
C10852 XM1/a_n158_28838# VSUBS 0.287142f
C10853 XM1/a_n100_28741# VSUBS 0.221608f
C10854 XM1/a_100_30274# VSUBS 0.287142f
C10855 XM1/a_n158_30274# VSUBS 0.287142f
C10856 XM1/a_n100_30177# VSUBS 0.221608f
C10857 XM1/a_100_31710# VSUBS 0.287142f
C10858 XM1/a_n158_31710# VSUBS 0.287142f
C10859 XM1/a_n100_31613# VSUBS 0.221608f
C10860 XM1/a_100_33146# VSUBS 0.287142f
C10861 XM1/a_n158_33146# VSUBS 0.287142f
C10862 XM1/a_n100_33049# VSUBS 0.221608f
C10863 XM1/a_100_34582# VSUBS 0.287142f
C10864 XM1/a_n158_34582# VSUBS 0.287142f
C10865 XM1/a_n100_34485# VSUBS 0.221608f
C10866 XM1/a_100_36018# VSUBS 0.287142f
C10867 XM1/a_n158_36018# VSUBS 0.287142f
C10868 XM1/a_n100_35921# VSUBS 0.221608f
C10869 XM1/a_100_37454# VSUBS 0.287142f
C10870 XM1/a_n158_37454# VSUBS 0.287142f
C10871 XM1/a_n100_37357# VSUBS 0.221608f
C10872 XM1/a_100_38890# VSUBS 0.287142f
C10873 XM1/a_n158_38890# VSUBS 0.287142f
C10874 XM1/a_n100_38793# VSUBS 0.221608f
C10875 XM1/a_100_40326# VSUBS 0.287142f
C10876 XM1/a_n158_40326# VSUBS 0.287142f
C10877 XM1/a_n100_40229# VSUBS 0.221608f
C10878 XM1/a_100_41762# VSUBS 0.287142f
C10879 XM1/a_n158_41762# VSUBS 0.287142f
C10880 XM1/a_n100_41665# VSUBS 0.221608f
C10881 XM1/a_100_43198# VSUBS 0.287142f
C10882 XM1/a_n158_43198# VSUBS 0.287142f
C10883 XM1/a_n100_43101# VSUBS 0.221608f
C10884 XM1/a_100_44634# VSUBS 0.287142f
C10885 XM1/a_n158_44634# VSUBS 0.287142f
C10886 XM1/a_n100_44537# VSUBS 0.221608f
C10887 XM1/a_100_46070# VSUBS 0.287142f
C10888 XM1/a_n158_46070# VSUBS 0.287142f
C10889 XM1/a_n100_45973# VSUBS 0.221608f
C10890 XM1/a_100_47506# VSUBS 0.287142f
C10891 XM1/a_n158_47506# VSUBS 0.287142f
C10892 XM1/a_n100_47409# VSUBS 0.221608f
C10893 XM1/a_100_48942# VSUBS 0.287142f
C10894 XM1/a_n158_48942# VSUBS 0.287142f
C10895 XM1/a_n100_48845# VSUBS 0.221608f
C10896 XM1/a_100_50378# VSUBS 0.287142f
C10897 XM1/a_n158_50378# VSUBS 0.287142f
C10898 XM1/a_n100_50281# VSUBS 0.221608f
C10899 XM1/a_100_51814# VSUBS 0.287142f
C10900 XM1/a_n158_51814# VSUBS 0.287142f
C10901 XM1/a_n100_51717# VSUBS 0.221608f
C10902 XM1/a_100_53250# VSUBS 0.287142f
C10903 XM1/a_n158_53250# VSUBS 0.287142f
C10904 XM1/a_n100_53153# VSUBS 0.221608f
C10905 XM1/a_100_54686# VSUBS 0.287142f
C10906 XM1/a_n158_54686# VSUBS 0.287142f
C10907 XM1/a_n100_54589# VSUBS 0.221608f
C10908 XM1/a_100_56122# VSUBS 0.287142f
C10909 XM1/a_n158_56122# VSUBS 0.287142f
C10910 XM1/a_n100_56025# VSUBS 0.221608f
C10911 XM1/a_100_57558# VSUBS 0.287142f
C10912 XM1/a_n158_57558# VSUBS 0.287142f
C10913 XM1/a_n100_57461# VSUBS 0.221608f
C10914 XM1/a_100_58994# VSUBS 0.287142f
C10915 XM1/a_n158_58994# VSUBS 0.287142f
C10916 XM1/a_n100_58897# VSUBS 0.221608f
C10917 XM1/a_100_60430# VSUBS 0.287142f
C10918 XM1/a_n158_60430# VSUBS 0.287142f
C10919 XM1/a_n100_60333# VSUBS 0.221608f
C10920 XM1/a_100_61866# VSUBS 0.287142f
C10921 XM1/a_n158_61866# VSUBS 0.287142f
C10922 XM1/a_n100_61769# VSUBS 0.221608f
C10923 XM1/a_100_63302# VSUBS 0.287142f
C10924 XM1/a_n158_63302# VSUBS 0.287142f
C10925 XM1/a_n100_63205# VSUBS 0.221608f
C10926 XM1/a_100_64738# VSUBS 0.287142f
C10927 XM1/a_n158_64738# VSUBS 0.287142f
C10928 XM1/a_n100_64641# VSUBS 0.221608f
C10929 XM1/a_100_66174# VSUBS 0.287142f
C10930 XM1/a_n158_66174# VSUBS 0.287142f
C10931 XM1/a_n100_66077# VSUBS 0.221608f
C10932 XM1/a_100_67610# VSUBS 0.287142f
C10933 XM1/a_n158_67610# VSUBS 0.287142f
C10934 XM1/a_n100_67513# VSUBS 0.221608f
C10935 XM1/a_100_69046# VSUBS 0.287142f
C10936 XM1/a_n158_69046# VSUBS 0.287142f
C10937 XM1/a_n100_68949# VSUBS 0.221608f
C10938 XM1/a_100_70482# VSUBS 0.287142f
C10939 XM1/a_n158_70482# VSUBS 0.287142f
C10940 XM1/a_n100_70385# VSUBS 0.221608f
C10941 XM1/a_100_71918# VSUBS 0.287142f
C10942 XM1/a_n158_71918# VSUBS 0.287142f
C10943 XM1/a_n100_71821# VSUBS 0.221608f
C10944 XM1/a_100_73354# VSUBS 0.287142f
C10945 XM1/a_n158_73354# VSUBS 0.287142f
C10946 XM1/a_n100_73257# VSUBS 0.221608f
C10947 XM1/a_100_74790# VSUBS 0.287142f
C10948 XM1/a_n158_74790# VSUBS 0.287142f
C10949 XM1/a_n100_74693# VSUBS 0.221608f
C10950 XM1/a_100_76226# VSUBS 0.287142f
C10951 XM1/a_n158_76226# VSUBS 0.287142f
C10952 XM1/a_n100_76129# VSUBS 0.221608f
C10953 XM1/a_100_77662# VSUBS 0.287142f
C10954 XM1/a_n158_77662# VSUBS 0.287142f
C10955 XM1/a_n100_77565# VSUBS 0.221608f
C10956 XM1/a_100_79098# VSUBS 0.287142f
C10957 XM1/a_n158_79098# VSUBS 0.287142f
C10958 XM1/a_n100_79001# VSUBS 0.221608f
C10959 XM1/a_100_80534# VSUBS 0.287142f
C10960 XM1/a_n158_80534# VSUBS 0.287142f
C10961 XM1/a_n100_80437# VSUBS 0.221608f
C10962 XM1/a_100_81970# VSUBS 0.287142f
C10963 XM1/a_n158_81970# VSUBS 0.287142f
C10964 XM1/a_n100_81873# VSUBS 0.221608f
C10965 XM1/a_100_83406# VSUBS 0.287142f
C10966 XM1/a_n158_83406# VSUBS 0.287142f
C10967 XM1/a_n100_83309# VSUBS 0.221608f
C10968 XM1/a_100_84842# VSUBS 0.287142f
C10969 XM1/a_n158_84842# VSUBS 0.287142f
C10970 XM1/a_n100_84745# VSUBS 0.221608f
C10971 XM1/a_100_86278# VSUBS 0.287142f
C10972 XM1/a_n158_86278# VSUBS 0.287142f
C10973 XM1/a_n100_86181# VSUBS 0.221608f
C10974 XM1/a_100_87714# VSUBS 0.287142f
C10975 XM1/a_n158_87714# VSUBS 0.287142f
C10976 XM1/a_n100_87617# VSUBS 0.221608f
C10977 XM1/a_100_89150# VSUBS 0.287142f
C10978 XM1/a_n158_89150# VSUBS 0.287142f
C10979 XM1/a_n100_89053# VSUBS 0.221608f
C10980 XM1/a_100_90586# VSUBS 0.287142f
C10981 XM1/a_n158_90586# VSUBS 0.287142f
C10982 XM1/a_n100_90489# VSUBS 0.221608f
C10983 XM1/a_100_92022# VSUBS 0.287142f
C10984 XM1/a_n158_92022# VSUBS 0.287142f
C10985 XM1/a_n100_91925# VSUBS 0.221608f
C10986 XM1/a_100_93458# VSUBS 0.287142f
C10987 XM1/a_n158_93458# VSUBS 0.287142f
C10988 XM1/a_n100_93361# VSUBS 0.221608f
C10989 XM1/a_100_94894# VSUBS 0.287142f
C10990 XM1/a_n158_94894# VSUBS 0.287142f
C10991 XM1/a_n100_94797# VSUBS 0.221608f
C10992 XM1/a_100_96330# VSUBS 0.287142f
C10993 XM1/a_n158_96330# VSUBS 0.287142f
C10994 XM1/a_n100_96233# VSUBS 0.221608f
C10995 XM1/a_100_97766# VSUBS 0.287142f
C10996 XM1/a_n158_97766# VSUBS 0.287142f
C10997 XM1/a_n100_97669# VSUBS 0.221608f
C10998 XM1/a_100_99202# VSUBS 0.287142f
C10999 XM1/a_n158_99202# VSUBS 0.287142f
C11000 XM1/a_n100_99105# VSUBS 0.221608f
C11001 XM1/a_100_100638# VSUBS 0.287142f
C11002 XM1/a_n158_100638# VSUBS 0.287142f
C11003 XM1/a_n100_100541# VSUBS 0.221608f
C11004 XM1/a_100_102074# VSUBS 0.287142f
C11005 XM1/a_n158_102074# VSUBS 0.287142f
C11006 XM1/a_n100_101977# VSUBS 0.221608f
C11007 XM1/a_100_103510# VSUBS 0.287142f
C11008 XM1/a_n158_103510# VSUBS 0.287142f
C11009 XM1/a_n100_103413# VSUBS 0.221608f
C11010 XM1/a_100_104946# VSUBS 0.287142f
C11011 XM1/a_n158_104946# VSUBS 0.287142f
C11012 XM1/a_n100_104849# VSUBS 0.221608f
C11013 XM1/a_100_106382# VSUBS 0.287142f
C11014 XM1/a_n158_106382# VSUBS 0.287142f
C11015 XM1/a_n100_106285# VSUBS 0.221608f
C11016 XM1/a_100_107818# VSUBS 0.287142f
C11017 XM1/a_n158_107818# VSUBS 0.287142f
C11018 XM1/a_n100_107721# VSUBS 0.221608f
C11019 XM1/a_100_109254# VSUBS 0.287142f
C11020 XM1/a_n158_109254# VSUBS 0.287142f
C11021 XM1/a_n100_109157# VSUBS 0.221608f
C11022 XM1/a_100_110690# VSUBS 0.287142f
C11023 XM1/a_n158_110690# VSUBS 0.287142f
C11024 XM1/a_n100_110593# VSUBS 0.221608f
C11025 XM1/a_100_112126# VSUBS 0.287142f
C11026 XM1/a_n158_112126# VSUBS 0.287142f
C11027 XM1/a_n100_112029# VSUBS 0.221608f
C11028 XM1/a_100_113562# VSUBS 0.287142f
C11029 XM1/a_n158_113562# VSUBS 0.287142f
C11030 XM1/a_n100_113465# VSUBS 0.221608f
C11031 XM1/a_100_114998# VSUBS 0.287142f
C11032 XM1/a_n158_114998# VSUBS 0.287142f
C11033 XM1/a_n100_114901# VSUBS 0.221608f
C11034 XM1/a_100_116434# VSUBS 0.287142f
C11035 XM1/a_n158_116434# VSUBS 0.287142f
C11036 XM1/a_n100_116337# VSUBS 0.221608f
C11037 XM1/a_100_117870# VSUBS 0.287142f
C11038 XM1/a_n158_117870# VSUBS 0.287142f
C11039 XM1/a_n100_117773# VSUBS 0.221608f
C11040 XM1/a_100_119306# VSUBS 0.287142f
C11041 XM1/a_n158_119306# VSUBS 0.287142f
C11042 XM1/a_n100_119209# VSUBS 0.221608f
C11043 XM1/a_100_120742# VSUBS 0.287142f
C11044 XM1/a_n158_120742# VSUBS 0.287142f
C11045 XM1/a_n100_120645# VSUBS 0.221608f
C11046 XM1/a_100_122178# VSUBS 0.287142f
C11047 XM1/a_n158_122178# VSUBS 0.287142f
C11048 XM1/a_n100_122081# VSUBS 0.221608f
C11049 XM1/a_100_123614# VSUBS 0.287142f
C11050 XM1/a_n158_123614# VSUBS 0.287142f
C11051 XM1/a_n100_123517# VSUBS 0.221608f
C11052 XM1/a_100_125050# VSUBS 0.287142f
C11053 XM1/a_n158_125050# VSUBS 0.287142f
C11054 XM1/a_n100_124953# VSUBS 0.221608f
C11055 XM1/a_100_126486# VSUBS 0.287142f
C11056 XM1/a_n158_126486# VSUBS 0.287142f
C11057 XM1/a_n100_126389# VSUBS 0.221608f
C11058 XM1/a_100_127922# VSUBS 0.287142f
C11059 XM1/a_n158_127922# VSUBS 0.287142f
C11060 XM1/a_n100_127825# VSUBS 0.221608f
C11061 XM1/a_100_129358# VSUBS 0.287142f
C11062 XM1/a_n158_129358# VSUBS 0.287142f
C11063 XM1/a_n100_129261# VSUBS 0.221608f
C11064 XM1/a_100_130794# VSUBS 0.287142f
C11065 XM1/a_n158_130794# VSUBS 0.287142f
C11066 XM1/a_n100_130697# VSUBS 0.221608f
C11067 XM1/a_100_132230# VSUBS 0.287142f
C11068 XM1/a_n158_132230# VSUBS 0.287142f
C11069 XM1/a_n100_132133# VSUBS 0.221608f
C11070 XM1/a_100_133666# VSUBS 0.287142f
C11071 XM1/a_n158_133666# VSUBS 0.287142f
C11072 XM1/a_n100_133569# VSUBS 0.221608f
C11073 XM1/a_100_135102# VSUBS 0.287142f
C11074 XM1/a_n158_135102# VSUBS 0.287142f
C11075 XM1/a_n100_135005# VSUBS 0.221608f
C11076 XM1/a_100_136538# VSUBS 0.287142f
C11077 XM1/a_n158_136538# VSUBS 0.287142f
C11078 XM1/a_n100_136441# VSUBS 0.221608f
C11079 XM1/a_100_137974# VSUBS 0.287142f
C11080 XM1/a_n158_137974# VSUBS 0.287142f
C11081 XM1/a_n100_137877# VSUBS 0.221608f
C11082 XM1/a_100_139410# VSUBS 0.287142f
C11083 XM1/a_n158_139410# VSUBS 0.287142f
C11084 XM1/a_n100_139313# VSUBS 0.221608f
C11085 XM1/a_100_140846# VSUBS 0.287142f
C11086 XM1/a_n158_140846# VSUBS 0.287142f
C11087 XM1/a_n100_140749# VSUBS 0.221608f
C11088 XM1/a_100_142282# VSUBS 0.287142f
C11089 XM1/a_n158_142282# VSUBS 0.287142f
C11090 XM1/a_n100_142185# VSUBS 0.221608f
C11091 XM1/a_100_143718# VSUBS 0.287142f
C11092 XM1/a_n158_143718# VSUBS 0.287142f
C11093 XM1/a_n100_143621# VSUBS 0.221608f
C11094 XM1/a_100_145154# VSUBS 0.287142f
C11095 XM1/a_n158_145154# VSUBS 0.287142f
C11096 XM1/a_n100_145057# VSUBS 0.221608f
C11097 XM1/a_100_146590# VSUBS 0.287142f
C11098 XM1/a_n158_146590# VSUBS 0.287142f
C11099 XM1/a_n100_146493# VSUBS 0.221608f
C11100 XM1/a_100_148026# VSUBS 0.287142f
C11101 XM1/a_n158_148026# VSUBS 0.287142f
C11102 XM1/a_n100_147929# VSUBS 0.221608f
C11103 XM1/a_100_149462# VSUBS 0.287142f
C11104 XM1/a_n158_149462# VSUBS 0.287142f
C11105 XM1/a_n100_149365# VSUBS 0.221608f
C11106 XM1/a_100_150898# VSUBS 0.287142f
C11107 XM1/a_n158_150898# VSUBS 0.287142f
C11108 XM1/a_n100_150801# VSUBS 0.221608f
C11109 XM1/a_100_152334# VSUBS 0.287142f
C11110 XM1/a_n158_152334# VSUBS 0.287142f
C11111 XM1/a_n100_152237# VSUBS 0.221608f
C11112 XM1/a_100_153770# VSUBS 0.287142f
C11113 XM1/a_n158_153770# VSUBS 0.287142f
C11114 XM1/a_n100_153673# VSUBS 0.221608f
C11115 XM1/a_100_155206# VSUBS 0.287142f
C11116 XM1/a_n158_155206# VSUBS 0.287142f
C11117 XM1/a_n100_155109# VSUBS 0.221608f
C11118 XM1/a_100_156642# VSUBS 0.287142f
C11119 XM1/a_n158_156642# VSUBS 0.287142f
C11120 XM1/a_n100_156545# VSUBS 0.221608f
C11121 XM1/a_100_158078# VSUBS 0.287142f
C11122 XM1/a_n158_158078# VSUBS 0.287142f
C11123 XM1/a_n100_157981# VSUBS 0.221608f
C11124 XM1/a_100_159514# VSUBS 0.287142f
C11125 XM1/a_n158_159514# VSUBS 0.287142f
C11126 XM1/a_n100_159417# VSUBS 0.221608f
C11127 XM1/a_100_160950# VSUBS 0.287142f
C11128 XM1/a_n158_160950# VSUBS 0.287142f
C11129 XM1/a_n100_160853# VSUBS 0.221608f
C11130 XM1/a_100_162386# VSUBS 0.287142f
C11131 XM1/a_n158_162386# VSUBS 0.287142f
C11132 XM1/a_n100_162289# VSUBS 0.221608f
C11133 XM1/a_100_163822# VSUBS 0.287142f
C11134 XM1/a_n158_163822# VSUBS 0.287142f
C11135 XM1/a_n100_163725# VSUBS 0.221608f
C11136 XM1/a_100_165258# VSUBS 0.287142f
C11137 XM1/a_n158_165258# VSUBS 0.287142f
C11138 XM1/a_n100_165161# VSUBS 0.221608f
C11139 XM1/a_100_166694# VSUBS 0.287142f
C11140 XM1/a_n158_166694# VSUBS 0.287142f
C11141 XM1/a_n100_166597# VSUBS 0.221608f
C11142 XM1/a_100_168130# VSUBS 0.287142f
C11143 XM1/a_n158_168130# VSUBS 0.287142f
C11144 XM1/a_n100_168033# VSUBS 0.221608f
C11145 XM1/a_100_169566# VSUBS 0.287142f
C11146 XM1/a_n158_169566# VSUBS 0.287142f
C11147 XM1/a_n100_169469# VSUBS 0.221608f
C11148 XM1/a_100_171002# VSUBS 0.287142f
C11149 XM1/a_n158_171002# VSUBS 0.287142f
C11150 XM1/a_n100_170905# VSUBS 0.221608f
C11151 XM1/a_100_172438# VSUBS 0.287142f
C11152 XM1/a_n158_172438# VSUBS 0.287142f
C11153 XM1/a_n100_172341# VSUBS 0.221608f
C11154 XM1/a_100_173874# VSUBS 0.287142f
C11155 XM1/a_n158_173874# VSUBS 0.287142f
C11156 XM1/a_n100_173777# VSUBS 0.221608f
C11157 XM1/a_100_175310# VSUBS 0.287142f
C11158 XM1/a_n158_175310# VSUBS 0.287142f
C11159 XM1/a_n100_175213# VSUBS 0.221608f
C11160 XM1/a_100_176746# VSUBS 0.287142f
C11161 XM1/a_n158_176746# VSUBS 0.287142f
C11162 XM1/a_n100_176649# VSUBS 0.221608f
C11163 XM1/a_100_178182# VSUBS 0.287142f
C11164 XM1/a_n158_178182# VSUBS 0.287142f
C11165 XM1/a_n100_178085# VSUBS 0.221608f
C11166 XM1/a_100_179618# VSUBS 0.287142f
C11167 XM1/a_n158_179618# VSUBS 0.287142f
C11168 XM1/a_n100_179521# VSUBS 0.221608f
C11169 XM1/a_100_181054# VSUBS 0.287142f
C11170 XM1/a_n158_181054# VSUBS 0.287142f
C11171 XM1/a_n100_180957# VSUBS 0.221608f
C11172 XM1/a_100_182490# VSUBS 0.292592f
C11173 XM1/a_n158_182490# VSUBS 0.292592f
C11174 XM1/a_n100_182393# VSUBS 0.265338f
.ends

