magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 16720 -2965 16836 -2899
rect 20064 -2965 20180 -2899
rect 23408 -2965 23524 -2899
rect 16572 -3232 16582 -3219
rect 16506 -3274 16582 -3232
rect 16634 -3274 16836 -3219
rect 16650 -3277 16836 -3274
rect 20180 -3219 20566 -3153
rect 23524 -3219 23910 -3153
rect 19916 -3232 19926 -3219
rect 19850 -3274 19926 -3232
rect 19978 -3274 20566 -3219
rect 23260 -3232 23270 -3219
rect 19850 -3277 20566 -3274
rect 16764 -3393 16964 -3385
rect 16780 -3397 16948 -3393
rect 16706 -3574 16806 -3450
rect 19850 -3514 19994 -3277
rect 20180 -3299 20566 -3277
rect 20104 -3385 20566 -3299
rect 23194 -3274 23270 -3232
rect 23322 -3274 23910 -3219
rect 26604 -3232 26614 -3219
rect 23194 -3277 23910 -3274
rect 20108 -3393 20308 -3385
rect 20124 -3397 20292 -3393
rect 16706 -3628 16708 -3574
rect 19850 -3600 20024 -3514
rect 20050 -3574 20150 -3450
rect 23194 -3514 23338 -3277
rect 23524 -3299 23910 -3277
rect 23448 -3385 23910 -3299
rect 26538 -3274 26614 -3232
rect 23452 -3393 23652 -3385
rect 23468 -3397 23636 -3393
rect 20050 -3628 20052 -3574
rect 23194 -3600 23368 -3514
rect 23394 -3574 23494 -3450
rect 26538 -3514 26682 -3274
rect 23394 -3628 23396 -3574
rect 26538 -3600 26712 -3514
rect 26738 -3574 26838 -3450
rect 26738 -3628 26740 -3574
rect 16391 -4371 16535 -4324
rect 16572 -4371 16589 -4270
rect 19735 -4371 19879 -4324
rect 19916 -4371 19933 -4270
rect 23079 -4371 23223 -4324
rect 23260 -4371 23277 -4270
rect 26423 -4371 26567 -4324
rect 26604 -4371 26621 -4270
rect 16391 -4382 16507 -4371
rect 16477 -4407 16507 -4382
rect 16489 -4906 16507 -4407
rect 19735 -4382 20507 -4371
rect 23079 -4382 23851 -4371
rect 26423 -4382 27195 -4371
rect 19821 -4407 20507 -4382
rect 23165 -4407 23851 -4382
rect 26509 -4407 27195 -4382
rect 19833 -4436 20507 -4407
rect 23177 -4436 23851 -4407
rect 26521 -4436 27195 -4407
rect 17671 -4848 17718 -4483
rect 17725 -4848 17772 -4537
rect 19833 -4848 20566 -4436
rect 21015 -4848 21062 -4483
rect 21069 -4848 21116 -4537
rect 23177 -4848 23910 -4436
rect 24359 -4848 24406 -4483
rect 24413 -4848 24460 -4537
rect 26521 -4848 27254 -4436
rect 27703 -4848 27750 -4483
rect 27757 -4848 27804 -4537
rect 17640 -4943 17843 -4848
rect 19833 -4906 21187 -4848
rect 23177 -4906 24531 -4848
rect 26521 -4906 27875 -4848
rect 19260 -4943 21187 -4906
rect 22604 -4943 24531 -4906
rect 25948 -4943 27875 -4906
rect 17640 -5067 18345 -4943
rect 19260 -5067 21689 -4943
rect 22604 -5067 25033 -4943
rect 25948 -5067 28377 -4943
rect 17640 -6152 18398 -5067
rect 19260 -6022 21742 -5067
rect 22604 -6022 25086 -5067
rect 25948 -6022 28430 -5067
rect 19851 -6087 21742 -6022
rect 23195 -6087 25086 -6022
rect 26539 -6087 28430 -6022
rect 20442 -6147 21742 -6087
rect 23786 -6147 25086 -6087
rect 27130 -6147 28430 -6087
rect 20471 -6152 21742 -6147
rect 23815 -6152 25086 -6147
rect 27159 -6152 28430 -6147
rect 17251 -6170 18398 -6152
rect 20595 -6170 21742 -6152
rect 23939 -6170 25086 -6152
rect 27283 -6170 28430 -6152
rect 17689 -6181 18398 -6170
rect 21033 -6181 21742 -6170
rect 24377 -6181 25086 -6170
rect 27721 -6181 28430 -6170
rect 17689 -6217 18363 -6181
rect 21033 -6217 21707 -6181
rect 24377 -6217 25051 -6181
rect 27721 -6217 28395 -6181
rect 17872 -6235 18363 -6217
rect 21216 -6235 21707 -6217
rect 24560 -6235 25051 -6217
rect 27904 -6235 28395 -6217
<< error_s >>
rect 3344 -2965 3460 -2899
rect 6688 -2965 6804 -2899
rect 10032 -2965 10148 -2899
rect 13376 -2965 13492 -2899
rect 3460 -3219 3846 -3153
rect 6804 -3219 7190 -3153
rect 10148 -3219 10534 -3153
rect 13492 -3219 13878 -3153
rect 3196 -3232 3206 -3219
rect 3130 -3274 3206 -3232
rect 3258 -3274 3846 -3219
rect 6540 -3232 6550 -3219
rect 3130 -3277 3846 -3274
rect 3130 -3514 3274 -3277
rect 3460 -3299 3846 -3277
rect 3384 -3385 3846 -3299
rect 6474 -3274 6550 -3232
rect 6602 -3274 7190 -3219
rect 9884 -3232 9894 -3219
rect 6474 -3277 7190 -3274
rect 3388 -3393 3588 -3385
rect 3404 -3397 3572 -3393
rect 3130 -3600 3304 -3514
rect 3330 -3574 3430 -3450
rect 6474 -3514 6618 -3277
rect 6804 -3299 7190 -3277
rect 6728 -3385 7190 -3299
rect 9818 -3274 9894 -3232
rect 9946 -3274 10534 -3219
rect 13228 -3232 13238 -3219
rect 9818 -3277 10534 -3274
rect 6732 -3393 6932 -3385
rect 6748 -3397 6916 -3393
rect 3330 -3628 3332 -3574
rect 6474 -3600 6648 -3514
rect 6674 -3574 6774 -3450
rect 9818 -3514 9962 -3277
rect 10148 -3299 10534 -3277
rect 10072 -3385 10534 -3299
rect 13162 -3274 13238 -3232
rect 13290 -3274 13878 -3219
rect 13162 -3277 13878 -3274
rect 10076 -3393 10276 -3385
rect 10092 -3397 10260 -3393
rect 6674 -3628 6676 -3574
rect 9818 -3600 9992 -3514
rect 10018 -3574 10118 -3450
rect 13162 -3514 13306 -3277
rect 13492 -3299 13878 -3277
rect 13416 -3385 13878 -3299
rect 13420 -3393 13620 -3385
rect 13436 -3397 13604 -3393
rect 10018 -3628 10020 -3574
rect 13162 -3600 13336 -3514
rect 13362 -3574 13462 -3450
rect 13362 -3628 13364 -3574
rect 3015 -4371 3159 -4324
rect 3196 -4371 3213 -4270
rect 6359 -4371 6503 -4324
rect 6540 -4371 6557 -4270
rect 9703 -4371 9847 -4324
rect 9884 -4371 9901 -4270
rect 13047 -4371 13191 -4324
rect 13228 -4371 13245 -4270
rect 3015 -4382 3787 -4371
rect 6359 -4382 7131 -4371
rect 9703 -4382 10475 -4371
rect 13047 -4382 13819 -4371
rect 3101 -4407 3787 -4382
rect 6445 -4407 7131 -4382
rect 9789 -4407 10475 -4382
rect 13133 -4407 13819 -4382
rect 3113 -4436 3787 -4407
rect 6457 -4436 7131 -4407
rect 9801 -4436 10475 -4407
rect 13145 -4436 13819 -4407
rect 3113 -4848 3846 -4436
rect 4295 -4848 4342 -4483
rect 4349 -4848 4396 -4537
rect 6457 -4848 7190 -4436
rect 7639 -4848 7686 -4483
rect 7693 -4848 7740 -4537
rect 9801 -4848 10534 -4436
rect 10983 -4848 11030 -4483
rect 11037 -4848 11084 -4537
rect 13145 -4848 13878 -4436
rect 14327 -4848 14374 -4483
rect 14381 -4848 14428 -4537
rect 3113 -4906 4467 -4848
rect 6457 -4906 7811 -4848
rect 9801 -4906 11155 -4848
rect 13145 -4906 14499 -4848
rect 2540 -4943 4467 -4906
rect 5884 -4943 7811 -4906
rect 9228 -4943 11155 -4906
rect 12572 -4943 14499 -4906
rect 2540 -5067 4969 -4943
rect 5884 -5067 8313 -4943
rect 9228 -5067 11657 -4943
rect 12572 -5067 15001 -4943
rect 2540 -6022 5022 -5067
rect 5884 -6022 8366 -5067
rect 9228 -6022 11710 -5067
rect 12572 -6022 15054 -5067
rect 15916 -6022 16380 -4906
rect 3131 -6087 5022 -6022
rect 6475 -6087 8366 -6022
rect 9819 -6087 11710 -6022
rect 13163 -6087 15054 -6022
rect 3722 -6147 5022 -6087
rect 7066 -6147 8366 -6087
rect 10410 -6147 11710 -6087
rect 13754 -6147 15054 -6087
rect 3751 -6152 5022 -6147
rect 7095 -6152 8366 -6147
rect 10439 -6152 11710 -6147
rect 13783 -6152 15054 -6147
rect 3875 -6170 5022 -6152
rect 7219 -6170 8366 -6152
rect 10563 -6170 11710 -6152
rect 13907 -6170 15054 -6152
rect 4313 -6181 5022 -6170
rect 7657 -6181 8366 -6170
rect 11001 -6181 11710 -6170
rect 14345 -6181 15054 -6170
rect 4313 -6217 4987 -6181
rect 7657 -6217 8331 -6181
rect 11001 -6217 11675 -6181
rect 14345 -6217 15019 -6181
rect 4496 -6235 4987 -6217
rect 7840 -6235 8331 -6217
rect 11184 -6235 11675 -6217
rect 14528 -6235 15019 -6217
<< error_ps >>
rect 16506 -3514 16650 -3274
rect 16836 -3299 17222 -3153
rect 16760 -3385 17222 -3299
rect 16506 -3600 16680 -3514
rect 16507 -4436 17163 -4371
rect 16507 -4848 17222 -4436
rect 16507 -4906 17640 -4848
rect 16380 -6022 17640 -4906
rect 16507 -6087 17640 -6022
rect 17098 -6147 17640 -6087
rect 17127 -6152 17640 -6147
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use icell4scs  x1
timestamp 1717439242
transform 1 0 0 0 1 0
box 0 -6337 15120 458
use icell4scs  x2
timestamp 1717439242
transform 1 0 13376 0 1 0
box 0 -6337 15120 458
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
