magic
tech sky130A
magscale 1 2
timestamp 1717414943
<< pwell >>
rect 149 -2436 805 -1930
rect 1239 -2272 1811 -2088
rect 149 -2472 806 -2436
rect 149 -2530 805 -2472
<< viali >>
rect 949 -2483 1317 -2448
<< metal1 >>
rect 149 -428 2514 -422
rect 149 -481 1599 -428
rect 1719 -481 2514 -428
rect 149 -622 2514 -481
rect 149 -656 2514 -650
rect 149 -709 2124 -656
rect 2244 -709 2514 -656
rect 149 -850 2514 -709
rect 1563 -987 1755 -980
rect 1563 -1040 1599 -987
rect 1719 -1040 1755 -987
rect 2089 -987 2281 -980
rect 2089 -1040 2124 -987
rect 2244 -1040 2281 -987
rect 307 -1500 371 -1488
rect 307 -1660 313 -1500
rect 365 -1660 371 -1500
rect 307 -1672 371 -1660
rect 583 -1672 1027 -1072
rect 382 -1710 573 -1704
rect 382 -1763 416 -1710
rect 536 -1763 573 -1710
rect 382 -1769 573 -1763
rect 1765 -2088 2079 -1072
rect 1239 -2100 1297 -2088
rect 1239 -2260 1245 -2100
rect 1239 -2272 1297 -2260
rect 1747 -2100 2079 -2088
rect 1747 -2260 1753 -2100
rect 1805 -2260 2079 -2100
rect 1747 -2271 2079 -2260
rect 1765 -2272 2079 -2271
rect 1036 -2357 1073 -2304
rect 1193 -2357 1229 -2304
rect 1036 -2363 1229 -2357
rect 1563 -2357 1599 -2304
rect 1719 -2357 1755 -2304
rect 1563 -2363 1755 -2357
rect 2089 -2357 2124 -2304
rect 2244 -2357 2281 -2304
rect 2089 -2363 2281 -2357
rect 149 -2448 2514 -2436
rect 149 -2470 949 -2448
rect 149 -2630 314 -2470
rect 366 -2483 949 -2470
rect 1317 -2483 2514 -2448
rect 366 -2630 2514 -2483
rect 149 -2636 2514 -2630
rect 149 -2805 2514 -2664
rect 149 -2858 1600 -2805
rect 1720 -2858 2514 -2805
rect 149 -2864 2514 -2858
rect 149 -3033 2514 -2892
rect 149 -3086 2125 -3033
rect 2245 -3086 2514 -3033
rect 149 -3092 2514 -3086
rect 149 -3261 2514 -3120
rect 149 -3314 417 -3261
rect 537 -3314 2514 -3261
rect 149 -3320 2514 -3314
rect 149 -3489 2514 -3348
rect 149 -3542 1074 -3489
rect 1194 -3542 2514 -3489
rect 149 -3548 2514 -3542
<< via1 >>
rect 1599 -481 1719 -428
rect 2124 -709 2244 -656
rect 1599 -1040 1719 -987
rect 2124 -1040 2244 -987
rect 313 -1660 365 -1500
rect 416 -1763 536 -1710
rect 1245 -2260 1297 -2100
rect 1753 -2260 1805 -2100
rect 1073 -2357 1193 -2304
rect 1599 -2357 1719 -2304
rect 2124 -2357 2244 -2304
rect 314 -2630 366 -2470
rect 1600 -2858 1720 -2805
rect 2125 -3086 2245 -3033
rect 417 -3314 537 -3261
rect 1074 -3542 1194 -3489
<< metal2 >>
rect 1593 -428 1725 -422
rect 1593 -481 1599 -428
rect 1719 -481 1725 -428
rect 1593 -987 1725 -481
rect 1593 -1040 1599 -987
rect 1719 -1040 1725 -987
rect 1593 -1046 1725 -1040
rect 2118 -656 2250 -650
rect 2118 -709 2124 -656
rect 2244 -709 2250 -656
rect 2118 -987 2250 -709
rect 2118 -1040 2124 -987
rect 2244 -1040 2250 -987
rect 2118 -1046 2250 -1040
rect 307 -1500 371 -1488
rect 307 -1660 313 -1500
rect 365 -1660 371 -1500
rect 307 -2470 371 -1660
rect 307 -2630 314 -2470
rect 366 -2630 371 -2470
rect 410 -1710 542 -1703
rect 410 -1763 416 -1710
rect 536 -1763 542 -1710
rect 410 -2436 542 -1763
rect 1239 -2100 1811 -2088
rect 1239 -2260 1245 -2100
rect 1297 -2260 1753 -2100
rect 1805 -2260 1811 -2100
rect 1239 -2270 1811 -2260
rect 1067 -2304 1199 -2298
rect 1067 -2357 1073 -2304
rect 1193 -2357 1199 -2304
rect 410 -2494 543 -2436
rect 307 -2636 371 -2630
rect 411 -3261 543 -2494
rect 411 -3314 417 -3261
rect 537 -3314 543 -3261
rect 411 -3320 543 -3314
rect 1067 -3489 1199 -2357
rect 1593 -2304 1725 -2298
rect 1593 -2357 1599 -2304
rect 1719 -2357 1725 -2304
rect 1593 -2805 1725 -2357
rect 1593 -2858 1600 -2805
rect 1720 -2858 1725 -2805
rect 1593 -2864 1725 -2858
rect 2118 -2304 2250 -2298
rect 2118 -2357 2124 -2304
rect 2244 -2357 2250 -2304
rect 2118 -3033 2250 -2357
rect 2118 -3086 2125 -3033
rect 2245 -3086 2250 -3033
rect 2118 -3092 2250 -3086
rect 1067 -3542 1074 -3489
rect 1194 -3542 1199 -3489
rect 1067 -3548 1199 -3542
use sky130_fd_pr__nfet_g5v0d10v5_BHMQGH  sky130_fd_pr__nfet_g5v0d10v5_BHMQGH_0
timestamp 1717401419
transform 1 0 1133 0 1 -1672
box -328 -858 328 858
use sky130_fd_pr__nfet_g5v0d10v5_D8TNYB  sky130_fd_pr__nfet_g5v0d10v5_D8TNYB_0
timestamp 1717401419
transform 1 0 477 0 1 -1372
box -328 -558 328 558
use sky130_fd_pr__nfet_g5v0d10v5_BHMQGH  XM1
timestamp 1717401419
transform 1 0 1659 0 1 -1672
box -328 -858 328 858
use sky130_fd_pr__nfet_g5v0d10v5_BHMQGH  XM2
timestamp 1717401419
transform 1 0 2185 0 1 -1672
box -328 -858 328 858
<< labels >>
flabel metal1 149 -2636 349 -2436 0 FreeSans 128 0 0 0 avss
port 6 nsew
flabel metal1 149 -2864 349 -2664 0 FreeSans 128 0 0 0 sw
port 3 nsew
flabel metal1 149 -3548 349 -3348 0 FreeSans 128 0 0 0 ncbias
port 4 nsew
flabel metal1 149 -3320 349 -3120 0 FreeSans 128 0 0 0 nbias
port 5 nsew
flabel metal1 149 -3092 349 -2892 0 FreeSans 128 0 0 0 swn
port 2 nsew
flabel metal1 149 -622 349 -422 0 FreeSans 128 0 0 0 iout
port 0 nsew
flabel metal1 149 -850 349 -650 0 FreeSans 128 0 0 0 ioutn
port 1 nsew
<< end >>
