magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< pwell >>
rect -328 -104853 328 104853
<< mvnmos >>
rect -100 103995 100 104595
rect -100 103177 100 103777
rect -100 102359 100 102959
rect -100 101541 100 102141
rect -100 100723 100 101323
rect -100 99905 100 100505
rect -100 99087 100 99687
rect -100 98269 100 98869
rect -100 97451 100 98051
rect -100 96633 100 97233
rect -100 95815 100 96415
rect -100 94997 100 95597
rect -100 94179 100 94779
rect -100 93361 100 93961
rect -100 92543 100 93143
rect -100 91725 100 92325
rect -100 90907 100 91507
rect -100 90089 100 90689
rect -100 89271 100 89871
rect -100 88453 100 89053
rect -100 87635 100 88235
rect -100 86817 100 87417
rect -100 85999 100 86599
rect -100 85181 100 85781
rect -100 84363 100 84963
rect -100 83545 100 84145
rect -100 82727 100 83327
rect -100 81909 100 82509
rect -100 81091 100 81691
rect -100 80273 100 80873
rect -100 79455 100 80055
rect -100 78637 100 79237
rect -100 77819 100 78419
rect -100 77001 100 77601
rect -100 76183 100 76783
rect -100 75365 100 75965
rect -100 74547 100 75147
rect -100 73729 100 74329
rect -100 72911 100 73511
rect -100 72093 100 72693
rect -100 71275 100 71875
rect -100 70457 100 71057
rect -100 69639 100 70239
rect -100 68821 100 69421
rect -100 68003 100 68603
rect -100 67185 100 67785
rect -100 66367 100 66967
rect -100 65549 100 66149
rect -100 64731 100 65331
rect -100 63913 100 64513
rect -100 63095 100 63695
rect -100 62277 100 62877
rect -100 61459 100 62059
rect -100 60641 100 61241
rect -100 59823 100 60423
rect -100 59005 100 59605
rect -100 58187 100 58787
rect -100 57369 100 57969
rect -100 56551 100 57151
rect -100 55733 100 56333
rect -100 54915 100 55515
rect -100 54097 100 54697
rect -100 53279 100 53879
rect -100 52461 100 53061
rect -100 51643 100 52243
rect -100 50825 100 51425
rect -100 50007 100 50607
rect -100 49189 100 49789
rect -100 48371 100 48971
rect -100 47553 100 48153
rect -100 46735 100 47335
rect -100 45917 100 46517
rect -100 45099 100 45699
rect -100 44281 100 44881
rect -100 43463 100 44063
rect -100 42645 100 43245
rect -100 41827 100 42427
rect -100 41009 100 41609
rect -100 40191 100 40791
rect -100 39373 100 39973
rect -100 38555 100 39155
rect -100 37737 100 38337
rect -100 36919 100 37519
rect -100 36101 100 36701
rect -100 35283 100 35883
rect -100 34465 100 35065
rect -100 33647 100 34247
rect -100 32829 100 33429
rect -100 32011 100 32611
rect -100 31193 100 31793
rect -100 30375 100 30975
rect -100 29557 100 30157
rect -100 28739 100 29339
rect -100 27921 100 28521
rect -100 27103 100 27703
rect -100 26285 100 26885
rect -100 25467 100 26067
rect -100 24649 100 25249
rect -100 23831 100 24431
rect -100 23013 100 23613
rect -100 22195 100 22795
rect -100 21377 100 21977
rect -100 20559 100 21159
rect -100 19741 100 20341
rect -100 18923 100 19523
rect -100 18105 100 18705
rect -100 17287 100 17887
rect -100 16469 100 17069
rect -100 15651 100 16251
rect -100 14833 100 15433
rect -100 14015 100 14615
rect -100 13197 100 13797
rect -100 12379 100 12979
rect -100 11561 100 12161
rect -100 10743 100 11343
rect -100 9925 100 10525
rect -100 9107 100 9707
rect -100 8289 100 8889
rect -100 7471 100 8071
rect -100 6653 100 7253
rect -100 5835 100 6435
rect -100 5017 100 5617
rect -100 4199 100 4799
rect -100 3381 100 3981
rect -100 2563 100 3163
rect -100 1745 100 2345
rect -100 927 100 1527
rect -100 109 100 709
rect -100 -709 100 -109
rect -100 -1527 100 -927
rect -100 -2345 100 -1745
rect -100 -3163 100 -2563
rect -100 -3981 100 -3381
rect -100 -4799 100 -4199
rect -100 -5617 100 -5017
rect -100 -6435 100 -5835
rect -100 -7253 100 -6653
rect -100 -8071 100 -7471
rect -100 -8889 100 -8289
rect -100 -9707 100 -9107
rect -100 -10525 100 -9925
rect -100 -11343 100 -10743
rect -100 -12161 100 -11561
rect -100 -12979 100 -12379
rect -100 -13797 100 -13197
rect -100 -14615 100 -14015
rect -100 -15433 100 -14833
rect -100 -16251 100 -15651
rect -100 -17069 100 -16469
rect -100 -17887 100 -17287
rect -100 -18705 100 -18105
rect -100 -19523 100 -18923
rect -100 -20341 100 -19741
rect -100 -21159 100 -20559
rect -100 -21977 100 -21377
rect -100 -22795 100 -22195
rect -100 -23613 100 -23013
rect -100 -24431 100 -23831
rect -100 -25249 100 -24649
rect -100 -26067 100 -25467
rect -100 -26885 100 -26285
rect -100 -27703 100 -27103
rect -100 -28521 100 -27921
rect -100 -29339 100 -28739
rect -100 -30157 100 -29557
rect -100 -30975 100 -30375
rect -100 -31793 100 -31193
rect -100 -32611 100 -32011
rect -100 -33429 100 -32829
rect -100 -34247 100 -33647
rect -100 -35065 100 -34465
rect -100 -35883 100 -35283
rect -100 -36701 100 -36101
rect -100 -37519 100 -36919
rect -100 -38337 100 -37737
rect -100 -39155 100 -38555
rect -100 -39973 100 -39373
rect -100 -40791 100 -40191
rect -100 -41609 100 -41009
rect -100 -42427 100 -41827
rect -100 -43245 100 -42645
rect -100 -44063 100 -43463
rect -100 -44881 100 -44281
rect -100 -45699 100 -45099
rect -100 -46517 100 -45917
rect -100 -47335 100 -46735
rect -100 -48153 100 -47553
rect -100 -48971 100 -48371
rect -100 -49789 100 -49189
rect -100 -50607 100 -50007
rect -100 -51425 100 -50825
rect -100 -52243 100 -51643
rect -100 -53061 100 -52461
rect -100 -53879 100 -53279
rect -100 -54697 100 -54097
rect -100 -55515 100 -54915
rect -100 -56333 100 -55733
rect -100 -57151 100 -56551
rect -100 -57969 100 -57369
rect -100 -58787 100 -58187
rect -100 -59605 100 -59005
rect -100 -60423 100 -59823
rect -100 -61241 100 -60641
rect -100 -62059 100 -61459
rect -100 -62877 100 -62277
rect -100 -63695 100 -63095
rect -100 -64513 100 -63913
rect -100 -65331 100 -64731
rect -100 -66149 100 -65549
rect -100 -66967 100 -66367
rect -100 -67785 100 -67185
rect -100 -68603 100 -68003
rect -100 -69421 100 -68821
rect -100 -70239 100 -69639
rect -100 -71057 100 -70457
rect -100 -71875 100 -71275
rect -100 -72693 100 -72093
rect -100 -73511 100 -72911
rect -100 -74329 100 -73729
rect -100 -75147 100 -74547
rect -100 -75965 100 -75365
rect -100 -76783 100 -76183
rect -100 -77601 100 -77001
rect -100 -78419 100 -77819
rect -100 -79237 100 -78637
rect -100 -80055 100 -79455
rect -100 -80873 100 -80273
rect -100 -81691 100 -81091
rect -100 -82509 100 -81909
rect -100 -83327 100 -82727
rect -100 -84145 100 -83545
rect -100 -84963 100 -84363
rect -100 -85781 100 -85181
rect -100 -86599 100 -85999
rect -100 -87417 100 -86817
rect -100 -88235 100 -87635
rect -100 -89053 100 -88453
rect -100 -89871 100 -89271
rect -100 -90689 100 -90089
rect -100 -91507 100 -90907
rect -100 -92325 100 -91725
rect -100 -93143 100 -92543
rect -100 -93961 100 -93361
rect -100 -94779 100 -94179
rect -100 -95597 100 -94997
rect -100 -96415 100 -95815
rect -100 -97233 100 -96633
rect -100 -98051 100 -97451
rect -100 -98869 100 -98269
rect -100 -99687 100 -99087
rect -100 -100505 100 -99905
rect -100 -101323 100 -100723
rect -100 -102141 100 -101541
rect -100 -102959 100 -102359
rect -100 -103777 100 -103177
rect -100 -104595 100 -103995
<< mvndiff >>
rect -158 104583 -100 104595
rect -158 104007 -146 104583
rect -112 104007 -100 104583
rect -158 103995 -100 104007
rect 100 104583 158 104595
rect 100 104007 112 104583
rect 146 104007 158 104583
rect 100 103995 158 104007
rect -158 103765 -100 103777
rect -158 103189 -146 103765
rect -112 103189 -100 103765
rect -158 103177 -100 103189
rect 100 103765 158 103777
rect 100 103189 112 103765
rect 146 103189 158 103765
rect 100 103177 158 103189
rect -158 102947 -100 102959
rect -158 102371 -146 102947
rect -112 102371 -100 102947
rect -158 102359 -100 102371
rect 100 102947 158 102959
rect 100 102371 112 102947
rect 146 102371 158 102947
rect 100 102359 158 102371
rect -158 102129 -100 102141
rect -158 101553 -146 102129
rect -112 101553 -100 102129
rect -158 101541 -100 101553
rect 100 102129 158 102141
rect 100 101553 112 102129
rect 146 101553 158 102129
rect 100 101541 158 101553
rect -158 101311 -100 101323
rect -158 100735 -146 101311
rect -112 100735 -100 101311
rect -158 100723 -100 100735
rect 100 101311 158 101323
rect 100 100735 112 101311
rect 146 100735 158 101311
rect 100 100723 158 100735
rect -158 100493 -100 100505
rect -158 99917 -146 100493
rect -112 99917 -100 100493
rect -158 99905 -100 99917
rect 100 100493 158 100505
rect 100 99917 112 100493
rect 146 99917 158 100493
rect 100 99905 158 99917
rect -158 99675 -100 99687
rect -158 99099 -146 99675
rect -112 99099 -100 99675
rect -158 99087 -100 99099
rect 100 99675 158 99687
rect 100 99099 112 99675
rect 146 99099 158 99675
rect 100 99087 158 99099
rect -158 98857 -100 98869
rect -158 98281 -146 98857
rect -112 98281 -100 98857
rect -158 98269 -100 98281
rect 100 98857 158 98869
rect 100 98281 112 98857
rect 146 98281 158 98857
rect 100 98269 158 98281
rect -158 98039 -100 98051
rect -158 97463 -146 98039
rect -112 97463 -100 98039
rect -158 97451 -100 97463
rect 100 98039 158 98051
rect 100 97463 112 98039
rect 146 97463 158 98039
rect 100 97451 158 97463
rect -158 97221 -100 97233
rect -158 96645 -146 97221
rect -112 96645 -100 97221
rect -158 96633 -100 96645
rect 100 97221 158 97233
rect 100 96645 112 97221
rect 146 96645 158 97221
rect 100 96633 158 96645
rect -158 96403 -100 96415
rect -158 95827 -146 96403
rect -112 95827 -100 96403
rect -158 95815 -100 95827
rect 100 96403 158 96415
rect 100 95827 112 96403
rect 146 95827 158 96403
rect 100 95815 158 95827
rect -158 95585 -100 95597
rect -158 95009 -146 95585
rect -112 95009 -100 95585
rect -158 94997 -100 95009
rect 100 95585 158 95597
rect 100 95009 112 95585
rect 146 95009 158 95585
rect 100 94997 158 95009
rect -158 94767 -100 94779
rect -158 94191 -146 94767
rect -112 94191 -100 94767
rect -158 94179 -100 94191
rect 100 94767 158 94779
rect 100 94191 112 94767
rect 146 94191 158 94767
rect 100 94179 158 94191
rect -158 93949 -100 93961
rect -158 93373 -146 93949
rect -112 93373 -100 93949
rect -158 93361 -100 93373
rect 100 93949 158 93961
rect 100 93373 112 93949
rect 146 93373 158 93949
rect 100 93361 158 93373
rect -158 93131 -100 93143
rect -158 92555 -146 93131
rect -112 92555 -100 93131
rect -158 92543 -100 92555
rect 100 93131 158 93143
rect 100 92555 112 93131
rect 146 92555 158 93131
rect 100 92543 158 92555
rect -158 92313 -100 92325
rect -158 91737 -146 92313
rect -112 91737 -100 92313
rect -158 91725 -100 91737
rect 100 92313 158 92325
rect 100 91737 112 92313
rect 146 91737 158 92313
rect 100 91725 158 91737
rect -158 91495 -100 91507
rect -158 90919 -146 91495
rect -112 90919 -100 91495
rect -158 90907 -100 90919
rect 100 91495 158 91507
rect 100 90919 112 91495
rect 146 90919 158 91495
rect 100 90907 158 90919
rect -158 90677 -100 90689
rect -158 90101 -146 90677
rect -112 90101 -100 90677
rect -158 90089 -100 90101
rect 100 90677 158 90689
rect 100 90101 112 90677
rect 146 90101 158 90677
rect 100 90089 158 90101
rect -158 89859 -100 89871
rect -158 89283 -146 89859
rect -112 89283 -100 89859
rect -158 89271 -100 89283
rect 100 89859 158 89871
rect 100 89283 112 89859
rect 146 89283 158 89859
rect 100 89271 158 89283
rect -158 89041 -100 89053
rect -158 88465 -146 89041
rect -112 88465 -100 89041
rect -158 88453 -100 88465
rect 100 89041 158 89053
rect 100 88465 112 89041
rect 146 88465 158 89041
rect 100 88453 158 88465
rect -158 88223 -100 88235
rect -158 87647 -146 88223
rect -112 87647 -100 88223
rect -158 87635 -100 87647
rect 100 88223 158 88235
rect 100 87647 112 88223
rect 146 87647 158 88223
rect 100 87635 158 87647
rect -158 87405 -100 87417
rect -158 86829 -146 87405
rect -112 86829 -100 87405
rect -158 86817 -100 86829
rect 100 87405 158 87417
rect 100 86829 112 87405
rect 146 86829 158 87405
rect 100 86817 158 86829
rect -158 86587 -100 86599
rect -158 86011 -146 86587
rect -112 86011 -100 86587
rect -158 85999 -100 86011
rect 100 86587 158 86599
rect 100 86011 112 86587
rect 146 86011 158 86587
rect 100 85999 158 86011
rect -158 85769 -100 85781
rect -158 85193 -146 85769
rect -112 85193 -100 85769
rect -158 85181 -100 85193
rect 100 85769 158 85781
rect 100 85193 112 85769
rect 146 85193 158 85769
rect 100 85181 158 85193
rect -158 84951 -100 84963
rect -158 84375 -146 84951
rect -112 84375 -100 84951
rect -158 84363 -100 84375
rect 100 84951 158 84963
rect 100 84375 112 84951
rect 146 84375 158 84951
rect 100 84363 158 84375
rect -158 84133 -100 84145
rect -158 83557 -146 84133
rect -112 83557 -100 84133
rect -158 83545 -100 83557
rect 100 84133 158 84145
rect 100 83557 112 84133
rect 146 83557 158 84133
rect 100 83545 158 83557
rect -158 83315 -100 83327
rect -158 82739 -146 83315
rect -112 82739 -100 83315
rect -158 82727 -100 82739
rect 100 83315 158 83327
rect 100 82739 112 83315
rect 146 82739 158 83315
rect 100 82727 158 82739
rect -158 82497 -100 82509
rect -158 81921 -146 82497
rect -112 81921 -100 82497
rect -158 81909 -100 81921
rect 100 82497 158 82509
rect 100 81921 112 82497
rect 146 81921 158 82497
rect 100 81909 158 81921
rect -158 81679 -100 81691
rect -158 81103 -146 81679
rect -112 81103 -100 81679
rect -158 81091 -100 81103
rect 100 81679 158 81691
rect 100 81103 112 81679
rect 146 81103 158 81679
rect 100 81091 158 81103
rect -158 80861 -100 80873
rect -158 80285 -146 80861
rect -112 80285 -100 80861
rect -158 80273 -100 80285
rect 100 80861 158 80873
rect 100 80285 112 80861
rect 146 80285 158 80861
rect 100 80273 158 80285
rect -158 80043 -100 80055
rect -158 79467 -146 80043
rect -112 79467 -100 80043
rect -158 79455 -100 79467
rect 100 80043 158 80055
rect 100 79467 112 80043
rect 146 79467 158 80043
rect 100 79455 158 79467
rect -158 79225 -100 79237
rect -158 78649 -146 79225
rect -112 78649 -100 79225
rect -158 78637 -100 78649
rect 100 79225 158 79237
rect 100 78649 112 79225
rect 146 78649 158 79225
rect 100 78637 158 78649
rect -158 78407 -100 78419
rect -158 77831 -146 78407
rect -112 77831 -100 78407
rect -158 77819 -100 77831
rect 100 78407 158 78419
rect 100 77831 112 78407
rect 146 77831 158 78407
rect 100 77819 158 77831
rect -158 77589 -100 77601
rect -158 77013 -146 77589
rect -112 77013 -100 77589
rect -158 77001 -100 77013
rect 100 77589 158 77601
rect 100 77013 112 77589
rect 146 77013 158 77589
rect 100 77001 158 77013
rect -158 76771 -100 76783
rect -158 76195 -146 76771
rect -112 76195 -100 76771
rect -158 76183 -100 76195
rect 100 76771 158 76783
rect 100 76195 112 76771
rect 146 76195 158 76771
rect 100 76183 158 76195
rect -158 75953 -100 75965
rect -158 75377 -146 75953
rect -112 75377 -100 75953
rect -158 75365 -100 75377
rect 100 75953 158 75965
rect 100 75377 112 75953
rect 146 75377 158 75953
rect 100 75365 158 75377
rect -158 75135 -100 75147
rect -158 74559 -146 75135
rect -112 74559 -100 75135
rect -158 74547 -100 74559
rect 100 75135 158 75147
rect 100 74559 112 75135
rect 146 74559 158 75135
rect 100 74547 158 74559
rect -158 74317 -100 74329
rect -158 73741 -146 74317
rect -112 73741 -100 74317
rect -158 73729 -100 73741
rect 100 74317 158 74329
rect 100 73741 112 74317
rect 146 73741 158 74317
rect 100 73729 158 73741
rect -158 73499 -100 73511
rect -158 72923 -146 73499
rect -112 72923 -100 73499
rect -158 72911 -100 72923
rect 100 73499 158 73511
rect 100 72923 112 73499
rect 146 72923 158 73499
rect 100 72911 158 72923
rect -158 72681 -100 72693
rect -158 72105 -146 72681
rect -112 72105 -100 72681
rect -158 72093 -100 72105
rect 100 72681 158 72693
rect 100 72105 112 72681
rect 146 72105 158 72681
rect 100 72093 158 72105
rect -158 71863 -100 71875
rect -158 71287 -146 71863
rect -112 71287 -100 71863
rect -158 71275 -100 71287
rect 100 71863 158 71875
rect 100 71287 112 71863
rect 146 71287 158 71863
rect 100 71275 158 71287
rect -158 71045 -100 71057
rect -158 70469 -146 71045
rect -112 70469 -100 71045
rect -158 70457 -100 70469
rect 100 71045 158 71057
rect 100 70469 112 71045
rect 146 70469 158 71045
rect 100 70457 158 70469
rect -158 70227 -100 70239
rect -158 69651 -146 70227
rect -112 69651 -100 70227
rect -158 69639 -100 69651
rect 100 70227 158 70239
rect 100 69651 112 70227
rect 146 69651 158 70227
rect 100 69639 158 69651
rect -158 69409 -100 69421
rect -158 68833 -146 69409
rect -112 68833 -100 69409
rect -158 68821 -100 68833
rect 100 69409 158 69421
rect 100 68833 112 69409
rect 146 68833 158 69409
rect 100 68821 158 68833
rect -158 68591 -100 68603
rect -158 68015 -146 68591
rect -112 68015 -100 68591
rect -158 68003 -100 68015
rect 100 68591 158 68603
rect 100 68015 112 68591
rect 146 68015 158 68591
rect 100 68003 158 68015
rect -158 67773 -100 67785
rect -158 67197 -146 67773
rect -112 67197 -100 67773
rect -158 67185 -100 67197
rect 100 67773 158 67785
rect 100 67197 112 67773
rect 146 67197 158 67773
rect 100 67185 158 67197
rect -158 66955 -100 66967
rect -158 66379 -146 66955
rect -112 66379 -100 66955
rect -158 66367 -100 66379
rect 100 66955 158 66967
rect 100 66379 112 66955
rect 146 66379 158 66955
rect 100 66367 158 66379
rect -158 66137 -100 66149
rect -158 65561 -146 66137
rect -112 65561 -100 66137
rect -158 65549 -100 65561
rect 100 66137 158 66149
rect 100 65561 112 66137
rect 146 65561 158 66137
rect 100 65549 158 65561
rect -158 65319 -100 65331
rect -158 64743 -146 65319
rect -112 64743 -100 65319
rect -158 64731 -100 64743
rect 100 65319 158 65331
rect 100 64743 112 65319
rect 146 64743 158 65319
rect 100 64731 158 64743
rect -158 64501 -100 64513
rect -158 63925 -146 64501
rect -112 63925 -100 64501
rect -158 63913 -100 63925
rect 100 64501 158 64513
rect 100 63925 112 64501
rect 146 63925 158 64501
rect 100 63913 158 63925
rect -158 63683 -100 63695
rect -158 63107 -146 63683
rect -112 63107 -100 63683
rect -158 63095 -100 63107
rect 100 63683 158 63695
rect 100 63107 112 63683
rect 146 63107 158 63683
rect 100 63095 158 63107
rect -158 62865 -100 62877
rect -158 62289 -146 62865
rect -112 62289 -100 62865
rect -158 62277 -100 62289
rect 100 62865 158 62877
rect 100 62289 112 62865
rect 146 62289 158 62865
rect 100 62277 158 62289
rect -158 62047 -100 62059
rect -158 61471 -146 62047
rect -112 61471 -100 62047
rect -158 61459 -100 61471
rect 100 62047 158 62059
rect 100 61471 112 62047
rect 146 61471 158 62047
rect 100 61459 158 61471
rect -158 61229 -100 61241
rect -158 60653 -146 61229
rect -112 60653 -100 61229
rect -158 60641 -100 60653
rect 100 61229 158 61241
rect 100 60653 112 61229
rect 146 60653 158 61229
rect 100 60641 158 60653
rect -158 60411 -100 60423
rect -158 59835 -146 60411
rect -112 59835 -100 60411
rect -158 59823 -100 59835
rect 100 60411 158 60423
rect 100 59835 112 60411
rect 146 59835 158 60411
rect 100 59823 158 59835
rect -158 59593 -100 59605
rect -158 59017 -146 59593
rect -112 59017 -100 59593
rect -158 59005 -100 59017
rect 100 59593 158 59605
rect 100 59017 112 59593
rect 146 59017 158 59593
rect 100 59005 158 59017
rect -158 58775 -100 58787
rect -158 58199 -146 58775
rect -112 58199 -100 58775
rect -158 58187 -100 58199
rect 100 58775 158 58787
rect 100 58199 112 58775
rect 146 58199 158 58775
rect 100 58187 158 58199
rect -158 57957 -100 57969
rect -158 57381 -146 57957
rect -112 57381 -100 57957
rect -158 57369 -100 57381
rect 100 57957 158 57969
rect 100 57381 112 57957
rect 146 57381 158 57957
rect 100 57369 158 57381
rect -158 57139 -100 57151
rect -158 56563 -146 57139
rect -112 56563 -100 57139
rect -158 56551 -100 56563
rect 100 57139 158 57151
rect 100 56563 112 57139
rect 146 56563 158 57139
rect 100 56551 158 56563
rect -158 56321 -100 56333
rect -158 55745 -146 56321
rect -112 55745 -100 56321
rect -158 55733 -100 55745
rect 100 56321 158 56333
rect 100 55745 112 56321
rect 146 55745 158 56321
rect 100 55733 158 55745
rect -158 55503 -100 55515
rect -158 54927 -146 55503
rect -112 54927 -100 55503
rect -158 54915 -100 54927
rect 100 55503 158 55515
rect 100 54927 112 55503
rect 146 54927 158 55503
rect 100 54915 158 54927
rect -158 54685 -100 54697
rect -158 54109 -146 54685
rect -112 54109 -100 54685
rect -158 54097 -100 54109
rect 100 54685 158 54697
rect 100 54109 112 54685
rect 146 54109 158 54685
rect 100 54097 158 54109
rect -158 53867 -100 53879
rect -158 53291 -146 53867
rect -112 53291 -100 53867
rect -158 53279 -100 53291
rect 100 53867 158 53879
rect 100 53291 112 53867
rect 146 53291 158 53867
rect 100 53279 158 53291
rect -158 53049 -100 53061
rect -158 52473 -146 53049
rect -112 52473 -100 53049
rect -158 52461 -100 52473
rect 100 53049 158 53061
rect 100 52473 112 53049
rect 146 52473 158 53049
rect 100 52461 158 52473
rect -158 52231 -100 52243
rect -158 51655 -146 52231
rect -112 51655 -100 52231
rect -158 51643 -100 51655
rect 100 52231 158 52243
rect 100 51655 112 52231
rect 146 51655 158 52231
rect 100 51643 158 51655
rect -158 51413 -100 51425
rect -158 50837 -146 51413
rect -112 50837 -100 51413
rect -158 50825 -100 50837
rect 100 51413 158 51425
rect 100 50837 112 51413
rect 146 50837 158 51413
rect 100 50825 158 50837
rect -158 50595 -100 50607
rect -158 50019 -146 50595
rect -112 50019 -100 50595
rect -158 50007 -100 50019
rect 100 50595 158 50607
rect 100 50019 112 50595
rect 146 50019 158 50595
rect 100 50007 158 50019
rect -158 49777 -100 49789
rect -158 49201 -146 49777
rect -112 49201 -100 49777
rect -158 49189 -100 49201
rect 100 49777 158 49789
rect 100 49201 112 49777
rect 146 49201 158 49777
rect 100 49189 158 49201
rect -158 48959 -100 48971
rect -158 48383 -146 48959
rect -112 48383 -100 48959
rect -158 48371 -100 48383
rect 100 48959 158 48971
rect 100 48383 112 48959
rect 146 48383 158 48959
rect 100 48371 158 48383
rect -158 48141 -100 48153
rect -158 47565 -146 48141
rect -112 47565 -100 48141
rect -158 47553 -100 47565
rect 100 48141 158 48153
rect 100 47565 112 48141
rect 146 47565 158 48141
rect 100 47553 158 47565
rect -158 47323 -100 47335
rect -158 46747 -146 47323
rect -112 46747 -100 47323
rect -158 46735 -100 46747
rect 100 47323 158 47335
rect 100 46747 112 47323
rect 146 46747 158 47323
rect 100 46735 158 46747
rect -158 46505 -100 46517
rect -158 45929 -146 46505
rect -112 45929 -100 46505
rect -158 45917 -100 45929
rect 100 46505 158 46517
rect 100 45929 112 46505
rect 146 45929 158 46505
rect 100 45917 158 45929
rect -158 45687 -100 45699
rect -158 45111 -146 45687
rect -112 45111 -100 45687
rect -158 45099 -100 45111
rect 100 45687 158 45699
rect 100 45111 112 45687
rect 146 45111 158 45687
rect 100 45099 158 45111
rect -158 44869 -100 44881
rect -158 44293 -146 44869
rect -112 44293 -100 44869
rect -158 44281 -100 44293
rect 100 44869 158 44881
rect 100 44293 112 44869
rect 146 44293 158 44869
rect 100 44281 158 44293
rect -158 44051 -100 44063
rect -158 43475 -146 44051
rect -112 43475 -100 44051
rect -158 43463 -100 43475
rect 100 44051 158 44063
rect 100 43475 112 44051
rect 146 43475 158 44051
rect 100 43463 158 43475
rect -158 43233 -100 43245
rect -158 42657 -146 43233
rect -112 42657 -100 43233
rect -158 42645 -100 42657
rect 100 43233 158 43245
rect 100 42657 112 43233
rect 146 42657 158 43233
rect 100 42645 158 42657
rect -158 42415 -100 42427
rect -158 41839 -146 42415
rect -112 41839 -100 42415
rect -158 41827 -100 41839
rect 100 42415 158 42427
rect 100 41839 112 42415
rect 146 41839 158 42415
rect 100 41827 158 41839
rect -158 41597 -100 41609
rect -158 41021 -146 41597
rect -112 41021 -100 41597
rect -158 41009 -100 41021
rect 100 41597 158 41609
rect 100 41021 112 41597
rect 146 41021 158 41597
rect 100 41009 158 41021
rect -158 40779 -100 40791
rect -158 40203 -146 40779
rect -112 40203 -100 40779
rect -158 40191 -100 40203
rect 100 40779 158 40791
rect 100 40203 112 40779
rect 146 40203 158 40779
rect 100 40191 158 40203
rect -158 39961 -100 39973
rect -158 39385 -146 39961
rect -112 39385 -100 39961
rect -158 39373 -100 39385
rect 100 39961 158 39973
rect 100 39385 112 39961
rect 146 39385 158 39961
rect 100 39373 158 39385
rect -158 39143 -100 39155
rect -158 38567 -146 39143
rect -112 38567 -100 39143
rect -158 38555 -100 38567
rect 100 39143 158 39155
rect 100 38567 112 39143
rect 146 38567 158 39143
rect 100 38555 158 38567
rect -158 38325 -100 38337
rect -158 37749 -146 38325
rect -112 37749 -100 38325
rect -158 37737 -100 37749
rect 100 38325 158 38337
rect 100 37749 112 38325
rect 146 37749 158 38325
rect 100 37737 158 37749
rect -158 37507 -100 37519
rect -158 36931 -146 37507
rect -112 36931 -100 37507
rect -158 36919 -100 36931
rect 100 37507 158 37519
rect 100 36931 112 37507
rect 146 36931 158 37507
rect 100 36919 158 36931
rect -158 36689 -100 36701
rect -158 36113 -146 36689
rect -112 36113 -100 36689
rect -158 36101 -100 36113
rect 100 36689 158 36701
rect 100 36113 112 36689
rect 146 36113 158 36689
rect 100 36101 158 36113
rect -158 35871 -100 35883
rect -158 35295 -146 35871
rect -112 35295 -100 35871
rect -158 35283 -100 35295
rect 100 35871 158 35883
rect 100 35295 112 35871
rect 146 35295 158 35871
rect 100 35283 158 35295
rect -158 35053 -100 35065
rect -158 34477 -146 35053
rect -112 34477 -100 35053
rect -158 34465 -100 34477
rect 100 35053 158 35065
rect 100 34477 112 35053
rect 146 34477 158 35053
rect 100 34465 158 34477
rect -158 34235 -100 34247
rect -158 33659 -146 34235
rect -112 33659 -100 34235
rect -158 33647 -100 33659
rect 100 34235 158 34247
rect 100 33659 112 34235
rect 146 33659 158 34235
rect 100 33647 158 33659
rect -158 33417 -100 33429
rect -158 32841 -146 33417
rect -112 32841 -100 33417
rect -158 32829 -100 32841
rect 100 33417 158 33429
rect 100 32841 112 33417
rect 146 32841 158 33417
rect 100 32829 158 32841
rect -158 32599 -100 32611
rect -158 32023 -146 32599
rect -112 32023 -100 32599
rect -158 32011 -100 32023
rect 100 32599 158 32611
rect 100 32023 112 32599
rect 146 32023 158 32599
rect 100 32011 158 32023
rect -158 31781 -100 31793
rect -158 31205 -146 31781
rect -112 31205 -100 31781
rect -158 31193 -100 31205
rect 100 31781 158 31793
rect 100 31205 112 31781
rect 146 31205 158 31781
rect 100 31193 158 31205
rect -158 30963 -100 30975
rect -158 30387 -146 30963
rect -112 30387 -100 30963
rect -158 30375 -100 30387
rect 100 30963 158 30975
rect 100 30387 112 30963
rect 146 30387 158 30963
rect 100 30375 158 30387
rect -158 30145 -100 30157
rect -158 29569 -146 30145
rect -112 29569 -100 30145
rect -158 29557 -100 29569
rect 100 30145 158 30157
rect 100 29569 112 30145
rect 146 29569 158 30145
rect 100 29557 158 29569
rect -158 29327 -100 29339
rect -158 28751 -146 29327
rect -112 28751 -100 29327
rect -158 28739 -100 28751
rect 100 29327 158 29339
rect 100 28751 112 29327
rect 146 28751 158 29327
rect 100 28739 158 28751
rect -158 28509 -100 28521
rect -158 27933 -146 28509
rect -112 27933 -100 28509
rect -158 27921 -100 27933
rect 100 28509 158 28521
rect 100 27933 112 28509
rect 146 27933 158 28509
rect 100 27921 158 27933
rect -158 27691 -100 27703
rect -158 27115 -146 27691
rect -112 27115 -100 27691
rect -158 27103 -100 27115
rect 100 27691 158 27703
rect 100 27115 112 27691
rect 146 27115 158 27691
rect 100 27103 158 27115
rect -158 26873 -100 26885
rect -158 26297 -146 26873
rect -112 26297 -100 26873
rect -158 26285 -100 26297
rect 100 26873 158 26885
rect 100 26297 112 26873
rect 146 26297 158 26873
rect 100 26285 158 26297
rect -158 26055 -100 26067
rect -158 25479 -146 26055
rect -112 25479 -100 26055
rect -158 25467 -100 25479
rect 100 26055 158 26067
rect 100 25479 112 26055
rect 146 25479 158 26055
rect 100 25467 158 25479
rect -158 25237 -100 25249
rect -158 24661 -146 25237
rect -112 24661 -100 25237
rect -158 24649 -100 24661
rect 100 25237 158 25249
rect 100 24661 112 25237
rect 146 24661 158 25237
rect 100 24649 158 24661
rect -158 24419 -100 24431
rect -158 23843 -146 24419
rect -112 23843 -100 24419
rect -158 23831 -100 23843
rect 100 24419 158 24431
rect 100 23843 112 24419
rect 146 23843 158 24419
rect 100 23831 158 23843
rect -158 23601 -100 23613
rect -158 23025 -146 23601
rect -112 23025 -100 23601
rect -158 23013 -100 23025
rect 100 23601 158 23613
rect 100 23025 112 23601
rect 146 23025 158 23601
rect 100 23013 158 23025
rect -158 22783 -100 22795
rect -158 22207 -146 22783
rect -112 22207 -100 22783
rect -158 22195 -100 22207
rect 100 22783 158 22795
rect 100 22207 112 22783
rect 146 22207 158 22783
rect 100 22195 158 22207
rect -158 21965 -100 21977
rect -158 21389 -146 21965
rect -112 21389 -100 21965
rect -158 21377 -100 21389
rect 100 21965 158 21977
rect 100 21389 112 21965
rect 146 21389 158 21965
rect 100 21377 158 21389
rect -158 21147 -100 21159
rect -158 20571 -146 21147
rect -112 20571 -100 21147
rect -158 20559 -100 20571
rect 100 21147 158 21159
rect 100 20571 112 21147
rect 146 20571 158 21147
rect 100 20559 158 20571
rect -158 20329 -100 20341
rect -158 19753 -146 20329
rect -112 19753 -100 20329
rect -158 19741 -100 19753
rect 100 20329 158 20341
rect 100 19753 112 20329
rect 146 19753 158 20329
rect 100 19741 158 19753
rect -158 19511 -100 19523
rect -158 18935 -146 19511
rect -112 18935 -100 19511
rect -158 18923 -100 18935
rect 100 19511 158 19523
rect 100 18935 112 19511
rect 146 18935 158 19511
rect 100 18923 158 18935
rect -158 18693 -100 18705
rect -158 18117 -146 18693
rect -112 18117 -100 18693
rect -158 18105 -100 18117
rect 100 18693 158 18705
rect 100 18117 112 18693
rect 146 18117 158 18693
rect 100 18105 158 18117
rect -158 17875 -100 17887
rect -158 17299 -146 17875
rect -112 17299 -100 17875
rect -158 17287 -100 17299
rect 100 17875 158 17887
rect 100 17299 112 17875
rect 146 17299 158 17875
rect 100 17287 158 17299
rect -158 17057 -100 17069
rect -158 16481 -146 17057
rect -112 16481 -100 17057
rect -158 16469 -100 16481
rect 100 17057 158 17069
rect 100 16481 112 17057
rect 146 16481 158 17057
rect 100 16469 158 16481
rect -158 16239 -100 16251
rect -158 15663 -146 16239
rect -112 15663 -100 16239
rect -158 15651 -100 15663
rect 100 16239 158 16251
rect 100 15663 112 16239
rect 146 15663 158 16239
rect 100 15651 158 15663
rect -158 15421 -100 15433
rect -158 14845 -146 15421
rect -112 14845 -100 15421
rect -158 14833 -100 14845
rect 100 15421 158 15433
rect 100 14845 112 15421
rect 146 14845 158 15421
rect 100 14833 158 14845
rect -158 14603 -100 14615
rect -158 14027 -146 14603
rect -112 14027 -100 14603
rect -158 14015 -100 14027
rect 100 14603 158 14615
rect 100 14027 112 14603
rect 146 14027 158 14603
rect 100 14015 158 14027
rect -158 13785 -100 13797
rect -158 13209 -146 13785
rect -112 13209 -100 13785
rect -158 13197 -100 13209
rect 100 13785 158 13797
rect 100 13209 112 13785
rect 146 13209 158 13785
rect 100 13197 158 13209
rect -158 12967 -100 12979
rect -158 12391 -146 12967
rect -112 12391 -100 12967
rect -158 12379 -100 12391
rect 100 12967 158 12979
rect 100 12391 112 12967
rect 146 12391 158 12967
rect 100 12379 158 12391
rect -158 12149 -100 12161
rect -158 11573 -146 12149
rect -112 11573 -100 12149
rect -158 11561 -100 11573
rect 100 12149 158 12161
rect 100 11573 112 12149
rect 146 11573 158 12149
rect 100 11561 158 11573
rect -158 11331 -100 11343
rect -158 10755 -146 11331
rect -112 10755 -100 11331
rect -158 10743 -100 10755
rect 100 11331 158 11343
rect 100 10755 112 11331
rect 146 10755 158 11331
rect 100 10743 158 10755
rect -158 10513 -100 10525
rect -158 9937 -146 10513
rect -112 9937 -100 10513
rect -158 9925 -100 9937
rect 100 10513 158 10525
rect 100 9937 112 10513
rect 146 9937 158 10513
rect 100 9925 158 9937
rect -158 9695 -100 9707
rect -158 9119 -146 9695
rect -112 9119 -100 9695
rect -158 9107 -100 9119
rect 100 9695 158 9707
rect 100 9119 112 9695
rect 146 9119 158 9695
rect 100 9107 158 9119
rect -158 8877 -100 8889
rect -158 8301 -146 8877
rect -112 8301 -100 8877
rect -158 8289 -100 8301
rect 100 8877 158 8889
rect 100 8301 112 8877
rect 146 8301 158 8877
rect 100 8289 158 8301
rect -158 8059 -100 8071
rect -158 7483 -146 8059
rect -112 7483 -100 8059
rect -158 7471 -100 7483
rect 100 8059 158 8071
rect 100 7483 112 8059
rect 146 7483 158 8059
rect 100 7471 158 7483
rect -158 7241 -100 7253
rect -158 6665 -146 7241
rect -112 6665 -100 7241
rect -158 6653 -100 6665
rect 100 7241 158 7253
rect 100 6665 112 7241
rect 146 6665 158 7241
rect 100 6653 158 6665
rect -158 6423 -100 6435
rect -158 5847 -146 6423
rect -112 5847 -100 6423
rect -158 5835 -100 5847
rect 100 6423 158 6435
rect 100 5847 112 6423
rect 146 5847 158 6423
rect 100 5835 158 5847
rect -158 5605 -100 5617
rect -158 5029 -146 5605
rect -112 5029 -100 5605
rect -158 5017 -100 5029
rect 100 5605 158 5617
rect 100 5029 112 5605
rect 146 5029 158 5605
rect 100 5017 158 5029
rect -158 4787 -100 4799
rect -158 4211 -146 4787
rect -112 4211 -100 4787
rect -158 4199 -100 4211
rect 100 4787 158 4799
rect 100 4211 112 4787
rect 146 4211 158 4787
rect 100 4199 158 4211
rect -158 3969 -100 3981
rect -158 3393 -146 3969
rect -112 3393 -100 3969
rect -158 3381 -100 3393
rect 100 3969 158 3981
rect 100 3393 112 3969
rect 146 3393 158 3969
rect 100 3381 158 3393
rect -158 3151 -100 3163
rect -158 2575 -146 3151
rect -112 2575 -100 3151
rect -158 2563 -100 2575
rect 100 3151 158 3163
rect 100 2575 112 3151
rect 146 2575 158 3151
rect 100 2563 158 2575
rect -158 2333 -100 2345
rect -158 1757 -146 2333
rect -112 1757 -100 2333
rect -158 1745 -100 1757
rect 100 2333 158 2345
rect 100 1757 112 2333
rect 146 1757 158 2333
rect 100 1745 158 1757
rect -158 1515 -100 1527
rect -158 939 -146 1515
rect -112 939 -100 1515
rect -158 927 -100 939
rect 100 1515 158 1527
rect 100 939 112 1515
rect 146 939 158 1515
rect 100 927 158 939
rect -158 697 -100 709
rect -158 121 -146 697
rect -112 121 -100 697
rect -158 109 -100 121
rect 100 697 158 709
rect 100 121 112 697
rect 146 121 158 697
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -697 -146 -121
rect -112 -697 -100 -121
rect -158 -709 -100 -697
rect 100 -121 158 -109
rect 100 -697 112 -121
rect 146 -697 158 -121
rect 100 -709 158 -697
rect -158 -939 -100 -927
rect -158 -1515 -146 -939
rect -112 -1515 -100 -939
rect -158 -1527 -100 -1515
rect 100 -939 158 -927
rect 100 -1515 112 -939
rect 146 -1515 158 -939
rect 100 -1527 158 -1515
rect -158 -1757 -100 -1745
rect -158 -2333 -146 -1757
rect -112 -2333 -100 -1757
rect -158 -2345 -100 -2333
rect 100 -1757 158 -1745
rect 100 -2333 112 -1757
rect 146 -2333 158 -1757
rect 100 -2345 158 -2333
rect -158 -2575 -100 -2563
rect -158 -3151 -146 -2575
rect -112 -3151 -100 -2575
rect -158 -3163 -100 -3151
rect 100 -2575 158 -2563
rect 100 -3151 112 -2575
rect 146 -3151 158 -2575
rect 100 -3163 158 -3151
rect -158 -3393 -100 -3381
rect -158 -3969 -146 -3393
rect -112 -3969 -100 -3393
rect -158 -3981 -100 -3969
rect 100 -3393 158 -3381
rect 100 -3969 112 -3393
rect 146 -3969 158 -3393
rect 100 -3981 158 -3969
rect -158 -4211 -100 -4199
rect -158 -4787 -146 -4211
rect -112 -4787 -100 -4211
rect -158 -4799 -100 -4787
rect 100 -4211 158 -4199
rect 100 -4787 112 -4211
rect 146 -4787 158 -4211
rect 100 -4799 158 -4787
rect -158 -5029 -100 -5017
rect -158 -5605 -146 -5029
rect -112 -5605 -100 -5029
rect -158 -5617 -100 -5605
rect 100 -5029 158 -5017
rect 100 -5605 112 -5029
rect 146 -5605 158 -5029
rect 100 -5617 158 -5605
rect -158 -5847 -100 -5835
rect -158 -6423 -146 -5847
rect -112 -6423 -100 -5847
rect -158 -6435 -100 -6423
rect 100 -5847 158 -5835
rect 100 -6423 112 -5847
rect 146 -6423 158 -5847
rect 100 -6435 158 -6423
rect -158 -6665 -100 -6653
rect -158 -7241 -146 -6665
rect -112 -7241 -100 -6665
rect -158 -7253 -100 -7241
rect 100 -6665 158 -6653
rect 100 -7241 112 -6665
rect 146 -7241 158 -6665
rect 100 -7253 158 -7241
rect -158 -7483 -100 -7471
rect -158 -8059 -146 -7483
rect -112 -8059 -100 -7483
rect -158 -8071 -100 -8059
rect 100 -7483 158 -7471
rect 100 -8059 112 -7483
rect 146 -8059 158 -7483
rect 100 -8071 158 -8059
rect -158 -8301 -100 -8289
rect -158 -8877 -146 -8301
rect -112 -8877 -100 -8301
rect -158 -8889 -100 -8877
rect 100 -8301 158 -8289
rect 100 -8877 112 -8301
rect 146 -8877 158 -8301
rect 100 -8889 158 -8877
rect -158 -9119 -100 -9107
rect -158 -9695 -146 -9119
rect -112 -9695 -100 -9119
rect -158 -9707 -100 -9695
rect 100 -9119 158 -9107
rect 100 -9695 112 -9119
rect 146 -9695 158 -9119
rect 100 -9707 158 -9695
rect -158 -9937 -100 -9925
rect -158 -10513 -146 -9937
rect -112 -10513 -100 -9937
rect -158 -10525 -100 -10513
rect 100 -9937 158 -9925
rect 100 -10513 112 -9937
rect 146 -10513 158 -9937
rect 100 -10525 158 -10513
rect -158 -10755 -100 -10743
rect -158 -11331 -146 -10755
rect -112 -11331 -100 -10755
rect -158 -11343 -100 -11331
rect 100 -10755 158 -10743
rect 100 -11331 112 -10755
rect 146 -11331 158 -10755
rect 100 -11343 158 -11331
rect -158 -11573 -100 -11561
rect -158 -12149 -146 -11573
rect -112 -12149 -100 -11573
rect -158 -12161 -100 -12149
rect 100 -11573 158 -11561
rect 100 -12149 112 -11573
rect 146 -12149 158 -11573
rect 100 -12161 158 -12149
rect -158 -12391 -100 -12379
rect -158 -12967 -146 -12391
rect -112 -12967 -100 -12391
rect -158 -12979 -100 -12967
rect 100 -12391 158 -12379
rect 100 -12967 112 -12391
rect 146 -12967 158 -12391
rect 100 -12979 158 -12967
rect -158 -13209 -100 -13197
rect -158 -13785 -146 -13209
rect -112 -13785 -100 -13209
rect -158 -13797 -100 -13785
rect 100 -13209 158 -13197
rect 100 -13785 112 -13209
rect 146 -13785 158 -13209
rect 100 -13797 158 -13785
rect -158 -14027 -100 -14015
rect -158 -14603 -146 -14027
rect -112 -14603 -100 -14027
rect -158 -14615 -100 -14603
rect 100 -14027 158 -14015
rect 100 -14603 112 -14027
rect 146 -14603 158 -14027
rect 100 -14615 158 -14603
rect -158 -14845 -100 -14833
rect -158 -15421 -146 -14845
rect -112 -15421 -100 -14845
rect -158 -15433 -100 -15421
rect 100 -14845 158 -14833
rect 100 -15421 112 -14845
rect 146 -15421 158 -14845
rect 100 -15433 158 -15421
rect -158 -15663 -100 -15651
rect -158 -16239 -146 -15663
rect -112 -16239 -100 -15663
rect -158 -16251 -100 -16239
rect 100 -15663 158 -15651
rect 100 -16239 112 -15663
rect 146 -16239 158 -15663
rect 100 -16251 158 -16239
rect -158 -16481 -100 -16469
rect -158 -17057 -146 -16481
rect -112 -17057 -100 -16481
rect -158 -17069 -100 -17057
rect 100 -16481 158 -16469
rect 100 -17057 112 -16481
rect 146 -17057 158 -16481
rect 100 -17069 158 -17057
rect -158 -17299 -100 -17287
rect -158 -17875 -146 -17299
rect -112 -17875 -100 -17299
rect -158 -17887 -100 -17875
rect 100 -17299 158 -17287
rect 100 -17875 112 -17299
rect 146 -17875 158 -17299
rect 100 -17887 158 -17875
rect -158 -18117 -100 -18105
rect -158 -18693 -146 -18117
rect -112 -18693 -100 -18117
rect -158 -18705 -100 -18693
rect 100 -18117 158 -18105
rect 100 -18693 112 -18117
rect 146 -18693 158 -18117
rect 100 -18705 158 -18693
rect -158 -18935 -100 -18923
rect -158 -19511 -146 -18935
rect -112 -19511 -100 -18935
rect -158 -19523 -100 -19511
rect 100 -18935 158 -18923
rect 100 -19511 112 -18935
rect 146 -19511 158 -18935
rect 100 -19523 158 -19511
rect -158 -19753 -100 -19741
rect -158 -20329 -146 -19753
rect -112 -20329 -100 -19753
rect -158 -20341 -100 -20329
rect 100 -19753 158 -19741
rect 100 -20329 112 -19753
rect 146 -20329 158 -19753
rect 100 -20341 158 -20329
rect -158 -20571 -100 -20559
rect -158 -21147 -146 -20571
rect -112 -21147 -100 -20571
rect -158 -21159 -100 -21147
rect 100 -20571 158 -20559
rect 100 -21147 112 -20571
rect 146 -21147 158 -20571
rect 100 -21159 158 -21147
rect -158 -21389 -100 -21377
rect -158 -21965 -146 -21389
rect -112 -21965 -100 -21389
rect -158 -21977 -100 -21965
rect 100 -21389 158 -21377
rect 100 -21965 112 -21389
rect 146 -21965 158 -21389
rect 100 -21977 158 -21965
rect -158 -22207 -100 -22195
rect -158 -22783 -146 -22207
rect -112 -22783 -100 -22207
rect -158 -22795 -100 -22783
rect 100 -22207 158 -22195
rect 100 -22783 112 -22207
rect 146 -22783 158 -22207
rect 100 -22795 158 -22783
rect -158 -23025 -100 -23013
rect -158 -23601 -146 -23025
rect -112 -23601 -100 -23025
rect -158 -23613 -100 -23601
rect 100 -23025 158 -23013
rect 100 -23601 112 -23025
rect 146 -23601 158 -23025
rect 100 -23613 158 -23601
rect -158 -23843 -100 -23831
rect -158 -24419 -146 -23843
rect -112 -24419 -100 -23843
rect -158 -24431 -100 -24419
rect 100 -23843 158 -23831
rect 100 -24419 112 -23843
rect 146 -24419 158 -23843
rect 100 -24431 158 -24419
rect -158 -24661 -100 -24649
rect -158 -25237 -146 -24661
rect -112 -25237 -100 -24661
rect -158 -25249 -100 -25237
rect 100 -24661 158 -24649
rect 100 -25237 112 -24661
rect 146 -25237 158 -24661
rect 100 -25249 158 -25237
rect -158 -25479 -100 -25467
rect -158 -26055 -146 -25479
rect -112 -26055 -100 -25479
rect -158 -26067 -100 -26055
rect 100 -25479 158 -25467
rect 100 -26055 112 -25479
rect 146 -26055 158 -25479
rect 100 -26067 158 -26055
rect -158 -26297 -100 -26285
rect -158 -26873 -146 -26297
rect -112 -26873 -100 -26297
rect -158 -26885 -100 -26873
rect 100 -26297 158 -26285
rect 100 -26873 112 -26297
rect 146 -26873 158 -26297
rect 100 -26885 158 -26873
rect -158 -27115 -100 -27103
rect -158 -27691 -146 -27115
rect -112 -27691 -100 -27115
rect -158 -27703 -100 -27691
rect 100 -27115 158 -27103
rect 100 -27691 112 -27115
rect 146 -27691 158 -27115
rect 100 -27703 158 -27691
rect -158 -27933 -100 -27921
rect -158 -28509 -146 -27933
rect -112 -28509 -100 -27933
rect -158 -28521 -100 -28509
rect 100 -27933 158 -27921
rect 100 -28509 112 -27933
rect 146 -28509 158 -27933
rect 100 -28521 158 -28509
rect -158 -28751 -100 -28739
rect -158 -29327 -146 -28751
rect -112 -29327 -100 -28751
rect -158 -29339 -100 -29327
rect 100 -28751 158 -28739
rect 100 -29327 112 -28751
rect 146 -29327 158 -28751
rect 100 -29339 158 -29327
rect -158 -29569 -100 -29557
rect -158 -30145 -146 -29569
rect -112 -30145 -100 -29569
rect -158 -30157 -100 -30145
rect 100 -29569 158 -29557
rect 100 -30145 112 -29569
rect 146 -30145 158 -29569
rect 100 -30157 158 -30145
rect -158 -30387 -100 -30375
rect -158 -30963 -146 -30387
rect -112 -30963 -100 -30387
rect -158 -30975 -100 -30963
rect 100 -30387 158 -30375
rect 100 -30963 112 -30387
rect 146 -30963 158 -30387
rect 100 -30975 158 -30963
rect -158 -31205 -100 -31193
rect -158 -31781 -146 -31205
rect -112 -31781 -100 -31205
rect -158 -31793 -100 -31781
rect 100 -31205 158 -31193
rect 100 -31781 112 -31205
rect 146 -31781 158 -31205
rect 100 -31793 158 -31781
rect -158 -32023 -100 -32011
rect -158 -32599 -146 -32023
rect -112 -32599 -100 -32023
rect -158 -32611 -100 -32599
rect 100 -32023 158 -32011
rect 100 -32599 112 -32023
rect 146 -32599 158 -32023
rect 100 -32611 158 -32599
rect -158 -32841 -100 -32829
rect -158 -33417 -146 -32841
rect -112 -33417 -100 -32841
rect -158 -33429 -100 -33417
rect 100 -32841 158 -32829
rect 100 -33417 112 -32841
rect 146 -33417 158 -32841
rect 100 -33429 158 -33417
rect -158 -33659 -100 -33647
rect -158 -34235 -146 -33659
rect -112 -34235 -100 -33659
rect -158 -34247 -100 -34235
rect 100 -33659 158 -33647
rect 100 -34235 112 -33659
rect 146 -34235 158 -33659
rect 100 -34247 158 -34235
rect -158 -34477 -100 -34465
rect -158 -35053 -146 -34477
rect -112 -35053 -100 -34477
rect -158 -35065 -100 -35053
rect 100 -34477 158 -34465
rect 100 -35053 112 -34477
rect 146 -35053 158 -34477
rect 100 -35065 158 -35053
rect -158 -35295 -100 -35283
rect -158 -35871 -146 -35295
rect -112 -35871 -100 -35295
rect -158 -35883 -100 -35871
rect 100 -35295 158 -35283
rect 100 -35871 112 -35295
rect 146 -35871 158 -35295
rect 100 -35883 158 -35871
rect -158 -36113 -100 -36101
rect -158 -36689 -146 -36113
rect -112 -36689 -100 -36113
rect -158 -36701 -100 -36689
rect 100 -36113 158 -36101
rect 100 -36689 112 -36113
rect 146 -36689 158 -36113
rect 100 -36701 158 -36689
rect -158 -36931 -100 -36919
rect -158 -37507 -146 -36931
rect -112 -37507 -100 -36931
rect -158 -37519 -100 -37507
rect 100 -36931 158 -36919
rect 100 -37507 112 -36931
rect 146 -37507 158 -36931
rect 100 -37519 158 -37507
rect -158 -37749 -100 -37737
rect -158 -38325 -146 -37749
rect -112 -38325 -100 -37749
rect -158 -38337 -100 -38325
rect 100 -37749 158 -37737
rect 100 -38325 112 -37749
rect 146 -38325 158 -37749
rect 100 -38337 158 -38325
rect -158 -38567 -100 -38555
rect -158 -39143 -146 -38567
rect -112 -39143 -100 -38567
rect -158 -39155 -100 -39143
rect 100 -38567 158 -38555
rect 100 -39143 112 -38567
rect 146 -39143 158 -38567
rect 100 -39155 158 -39143
rect -158 -39385 -100 -39373
rect -158 -39961 -146 -39385
rect -112 -39961 -100 -39385
rect -158 -39973 -100 -39961
rect 100 -39385 158 -39373
rect 100 -39961 112 -39385
rect 146 -39961 158 -39385
rect 100 -39973 158 -39961
rect -158 -40203 -100 -40191
rect -158 -40779 -146 -40203
rect -112 -40779 -100 -40203
rect -158 -40791 -100 -40779
rect 100 -40203 158 -40191
rect 100 -40779 112 -40203
rect 146 -40779 158 -40203
rect 100 -40791 158 -40779
rect -158 -41021 -100 -41009
rect -158 -41597 -146 -41021
rect -112 -41597 -100 -41021
rect -158 -41609 -100 -41597
rect 100 -41021 158 -41009
rect 100 -41597 112 -41021
rect 146 -41597 158 -41021
rect 100 -41609 158 -41597
rect -158 -41839 -100 -41827
rect -158 -42415 -146 -41839
rect -112 -42415 -100 -41839
rect -158 -42427 -100 -42415
rect 100 -41839 158 -41827
rect 100 -42415 112 -41839
rect 146 -42415 158 -41839
rect 100 -42427 158 -42415
rect -158 -42657 -100 -42645
rect -158 -43233 -146 -42657
rect -112 -43233 -100 -42657
rect -158 -43245 -100 -43233
rect 100 -42657 158 -42645
rect 100 -43233 112 -42657
rect 146 -43233 158 -42657
rect 100 -43245 158 -43233
rect -158 -43475 -100 -43463
rect -158 -44051 -146 -43475
rect -112 -44051 -100 -43475
rect -158 -44063 -100 -44051
rect 100 -43475 158 -43463
rect 100 -44051 112 -43475
rect 146 -44051 158 -43475
rect 100 -44063 158 -44051
rect -158 -44293 -100 -44281
rect -158 -44869 -146 -44293
rect -112 -44869 -100 -44293
rect -158 -44881 -100 -44869
rect 100 -44293 158 -44281
rect 100 -44869 112 -44293
rect 146 -44869 158 -44293
rect 100 -44881 158 -44869
rect -158 -45111 -100 -45099
rect -158 -45687 -146 -45111
rect -112 -45687 -100 -45111
rect -158 -45699 -100 -45687
rect 100 -45111 158 -45099
rect 100 -45687 112 -45111
rect 146 -45687 158 -45111
rect 100 -45699 158 -45687
rect -158 -45929 -100 -45917
rect -158 -46505 -146 -45929
rect -112 -46505 -100 -45929
rect -158 -46517 -100 -46505
rect 100 -45929 158 -45917
rect 100 -46505 112 -45929
rect 146 -46505 158 -45929
rect 100 -46517 158 -46505
rect -158 -46747 -100 -46735
rect -158 -47323 -146 -46747
rect -112 -47323 -100 -46747
rect -158 -47335 -100 -47323
rect 100 -46747 158 -46735
rect 100 -47323 112 -46747
rect 146 -47323 158 -46747
rect 100 -47335 158 -47323
rect -158 -47565 -100 -47553
rect -158 -48141 -146 -47565
rect -112 -48141 -100 -47565
rect -158 -48153 -100 -48141
rect 100 -47565 158 -47553
rect 100 -48141 112 -47565
rect 146 -48141 158 -47565
rect 100 -48153 158 -48141
rect -158 -48383 -100 -48371
rect -158 -48959 -146 -48383
rect -112 -48959 -100 -48383
rect -158 -48971 -100 -48959
rect 100 -48383 158 -48371
rect 100 -48959 112 -48383
rect 146 -48959 158 -48383
rect 100 -48971 158 -48959
rect -158 -49201 -100 -49189
rect -158 -49777 -146 -49201
rect -112 -49777 -100 -49201
rect -158 -49789 -100 -49777
rect 100 -49201 158 -49189
rect 100 -49777 112 -49201
rect 146 -49777 158 -49201
rect 100 -49789 158 -49777
rect -158 -50019 -100 -50007
rect -158 -50595 -146 -50019
rect -112 -50595 -100 -50019
rect -158 -50607 -100 -50595
rect 100 -50019 158 -50007
rect 100 -50595 112 -50019
rect 146 -50595 158 -50019
rect 100 -50607 158 -50595
rect -158 -50837 -100 -50825
rect -158 -51413 -146 -50837
rect -112 -51413 -100 -50837
rect -158 -51425 -100 -51413
rect 100 -50837 158 -50825
rect 100 -51413 112 -50837
rect 146 -51413 158 -50837
rect 100 -51425 158 -51413
rect -158 -51655 -100 -51643
rect -158 -52231 -146 -51655
rect -112 -52231 -100 -51655
rect -158 -52243 -100 -52231
rect 100 -51655 158 -51643
rect 100 -52231 112 -51655
rect 146 -52231 158 -51655
rect 100 -52243 158 -52231
rect -158 -52473 -100 -52461
rect -158 -53049 -146 -52473
rect -112 -53049 -100 -52473
rect -158 -53061 -100 -53049
rect 100 -52473 158 -52461
rect 100 -53049 112 -52473
rect 146 -53049 158 -52473
rect 100 -53061 158 -53049
rect -158 -53291 -100 -53279
rect -158 -53867 -146 -53291
rect -112 -53867 -100 -53291
rect -158 -53879 -100 -53867
rect 100 -53291 158 -53279
rect 100 -53867 112 -53291
rect 146 -53867 158 -53291
rect 100 -53879 158 -53867
rect -158 -54109 -100 -54097
rect -158 -54685 -146 -54109
rect -112 -54685 -100 -54109
rect -158 -54697 -100 -54685
rect 100 -54109 158 -54097
rect 100 -54685 112 -54109
rect 146 -54685 158 -54109
rect 100 -54697 158 -54685
rect -158 -54927 -100 -54915
rect -158 -55503 -146 -54927
rect -112 -55503 -100 -54927
rect -158 -55515 -100 -55503
rect 100 -54927 158 -54915
rect 100 -55503 112 -54927
rect 146 -55503 158 -54927
rect 100 -55515 158 -55503
rect -158 -55745 -100 -55733
rect -158 -56321 -146 -55745
rect -112 -56321 -100 -55745
rect -158 -56333 -100 -56321
rect 100 -55745 158 -55733
rect 100 -56321 112 -55745
rect 146 -56321 158 -55745
rect 100 -56333 158 -56321
rect -158 -56563 -100 -56551
rect -158 -57139 -146 -56563
rect -112 -57139 -100 -56563
rect -158 -57151 -100 -57139
rect 100 -56563 158 -56551
rect 100 -57139 112 -56563
rect 146 -57139 158 -56563
rect 100 -57151 158 -57139
rect -158 -57381 -100 -57369
rect -158 -57957 -146 -57381
rect -112 -57957 -100 -57381
rect -158 -57969 -100 -57957
rect 100 -57381 158 -57369
rect 100 -57957 112 -57381
rect 146 -57957 158 -57381
rect 100 -57969 158 -57957
rect -158 -58199 -100 -58187
rect -158 -58775 -146 -58199
rect -112 -58775 -100 -58199
rect -158 -58787 -100 -58775
rect 100 -58199 158 -58187
rect 100 -58775 112 -58199
rect 146 -58775 158 -58199
rect 100 -58787 158 -58775
rect -158 -59017 -100 -59005
rect -158 -59593 -146 -59017
rect -112 -59593 -100 -59017
rect -158 -59605 -100 -59593
rect 100 -59017 158 -59005
rect 100 -59593 112 -59017
rect 146 -59593 158 -59017
rect 100 -59605 158 -59593
rect -158 -59835 -100 -59823
rect -158 -60411 -146 -59835
rect -112 -60411 -100 -59835
rect -158 -60423 -100 -60411
rect 100 -59835 158 -59823
rect 100 -60411 112 -59835
rect 146 -60411 158 -59835
rect 100 -60423 158 -60411
rect -158 -60653 -100 -60641
rect -158 -61229 -146 -60653
rect -112 -61229 -100 -60653
rect -158 -61241 -100 -61229
rect 100 -60653 158 -60641
rect 100 -61229 112 -60653
rect 146 -61229 158 -60653
rect 100 -61241 158 -61229
rect -158 -61471 -100 -61459
rect -158 -62047 -146 -61471
rect -112 -62047 -100 -61471
rect -158 -62059 -100 -62047
rect 100 -61471 158 -61459
rect 100 -62047 112 -61471
rect 146 -62047 158 -61471
rect 100 -62059 158 -62047
rect -158 -62289 -100 -62277
rect -158 -62865 -146 -62289
rect -112 -62865 -100 -62289
rect -158 -62877 -100 -62865
rect 100 -62289 158 -62277
rect 100 -62865 112 -62289
rect 146 -62865 158 -62289
rect 100 -62877 158 -62865
rect -158 -63107 -100 -63095
rect -158 -63683 -146 -63107
rect -112 -63683 -100 -63107
rect -158 -63695 -100 -63683
rect 100 -63107 158 -63095
rect 100 -63683 112 -63107
rect 146 -63683 158 -63107
rect 100 -63695 158 -63683
rect -158 -63925 -100 -63913
rect -158 -64501 -146 -63925
rect -112 -64501 -100 -63925
rect -158 -64513 -100 -64501
rect 100 -63925 158 -63913
rect 100 -64501 112 -63925
rect 146 -64501 158 -63925
rect 100 -64513 158 -64501
rect -158 -64743 -100 -64731
rect -158 -65319 -146 -64743
rect -112 -65319 -100 -64743
rect -158 -65331 -100 -65319
rect 100 -64743 158 -64731
rect 100 -65319 112 -64743
rect 146 -65319 158 -64743
rect 100 -65331 158 -65319
rect -158 -65561 -100 -65549
rect -158 -66137 -146 -65561
rect -112 -66137 -100 -65561
rect -158 -66149 -100 -66137
rect 100 -65561 158 -65549
rect 100 -66137 112 -65561
rect 146 -66137 158 -65561
rect 100 -66149 158 -66137
rect -158 -66379 -100 -66367
rect -158 -66955 -146 -66379
rect -112 -66955 -100 -66379
rect -158 -66967 -100 -66955
rect 100 -66379 158 -66367
rect 100 -66955 112 -66379
rect 146 -66955 158 -66379
rect 100 -66967 158 -66955
rect -158 -67197 -100 -67185
rect -158 -67773 -146 -67197
rect -112 -67773 -100 -67197
rect -158 -67785 -100 -67773
rect 100 -67197 158 -67185
rect 100 -67773 112 -67197
rect 146 -67773 158 -67197
rect 100 -67785 158 -67773
rect -158 -68015 -100 -68003
rect -158 -68591 -146 -68015
rect -112 -68591 -100 -68015
rect -158 -68603 -100 -68591
rect 100 -68015 158 -68003
rect 100 -68591 112 -68015
rect 146 -68591 158 -68015
rect 100 -68603 158 -68591
rect -158 -68833 -100 -68821
rect -158 -69409 -146 -68833
rect -112 -69409 -100 -68833
rect -158 -69421 -100 -69409
rect 100 -68833 158 -68821
rect 100 -69409 112 -68833
rect 146 -69409 158 -68833
rect 100 -69421 158 -69409
rect -158 -69651 -100 -69639
rect -158 -70227 -146 -69651
rect -112 -70227 -100 -69651
rect -158 -70239 -100 -70227
rect 100 -69651 158 -69639
rect 100 -70227 112 -69651
rect 146 -70227 158 -69651
rect 100 -70239 158 -70227
rect -158 -70469 -100 -70457
rect -158 -71045 -146 -70469
rect -112 -71045 -100 -70469
rect -158 -71057 -100 -71045
rect 100 -70469 158 -70457
rect 100 -71045 112 -70469
rect 146 -71045 158 -70469
rect 100 -71057 158 -71045
rect -158 -71287 -100 -71275
rect -158 -71863 -146 -71287
rect -112 -71863 -100 -71287
rect -158 -71875 -100 -71863
rect 100 -71287 158 -71275
rect 100 -71863 112 -71287
rect 146 -71863 158 -71287
rect 100 -71875 158 -71863
rect -158 -72105 -100 -72093
rect -158 -72681 -146 -72105
rect -112 -72681 -100 -72105
rect -158 -72693 -100 -72681
rect 100 -72105 158 -72093
rect 100 -72681 112 -72105
rect 146 -72681 158 -72105
rect 100 -72693 158 -72681
rect -158 -72923 -100 -72911
rect -158 -73499 -146 -72923
rect -112 -73499 -100 -72923
rect -158 -73511 -100 -73499
rect 100 -72923 158 -72911
rect 100 -73499 112 -72923
rect 146 -73499 158 -72923
rect 100 -73511 158 -73499
rect -158 -73741 -100 -73729
rect -158 -74317 -146 -73741
rect -112 -74317 -100 -73741
rect -158 -74329 -100 -74317
rect 100 -73741 158 -73729
rect 100 -74317 112 -73741
rect 146 -74317 158 -73741
rect 100 -74329 158 -74317
rect -158 -74559 -100 -74547
rect -158 -75135 -146 -74559
rect -112 -75135 -100 -74559
rect -158 -75147 -100 -75135
rect 100 -74559 158 -74547
rect 100 -75135 112 -74559
rect 146 -75135 158 -74559
rect 100 -75147 158 -75135
rect -158 -75377 -100 -75365
rect -158 -75953 -146 -75377
rect -112 -75953 -100 -75377
rect -158 -75965 -100 -75953
rect 100 -75377 158 -75365
rect 100 -75953 112 -75377
rect 146 -75953 158 -75377
rect 100 -75965 158 -75953
rect -158 -76195 -100 -76183
rect -158 -76771 -146 -76195
rect -112 -76771 -100 -76195
rect -158 -76783 -100 -76771
rect 100 -76195 158 -76183
rect 100 -76771 112 -76195
rect 146 -76771 158 -76195
rect 100 -76783 158 -76771
rect -158 -77013 -100 -77001
rect -158 -77589 -146 -77013
rect -112 -77589 -100 -77013
rect -158 -77601 -100 -77589
rect 100 -77013 158 -77001
rect 100 -77589 112 -77013
rect 146 -77589 158 -77013
rect 100 -77601 158 -77589
rect -158 -77831 -100 -77819
rect -158 -78407 -146 -77831
rect -112 -78407 -100 -77831
rect -158 -78419 -100 -78407
rect 100 -77831 158 -77819
rect 100 -78407 112 -77831
rect 146 -78407 158 -77831
rect 100 -78419 158 -78407
rect -158 -78649 -100 -78637
rect -158 -79225 -146 -78649
rect -112 -79225 -100 -78649
rect -158 -79237 -100 -79225
rect 100 -78649 158 -78637
rect 100 -79225 112 -78649
rect 146 -79225 158 -78649
rect 100 -79237 158 -79225
rect -158 -79467 -100 -79455
rect -158 -80043 -146 -79467
rect -112 -80043 -100 -79467
rect -158 -80055 -100 -80043
rect 100 -79467 158 -79455
rect 100 -80043 112 -79467
rect 146 -80043 158 -79467
rect 100 -80055 158 -80043
rect -158 -80285 -100 -80273
rect -158 -80861 -146 -80285
rect -112 -80861 -100 -80285
rect -158 -80873 -100 -80861
rect 100 -80285 158 -80273
rect 100 -80861 112 -80285
rect 146 -80861 158 -80285
rect 100 -80873 158 -80861
rect -158 -81103 -100 -81091
rect -158 -81679 -146 -81103
rect -112 -81679 -100 -81103
rect -158 -81691 -100 -81679
rect 100 -81103 158 -81091
rect 100 -81679 112 -81103
rect 146 -81679 158 -81103
rect 100 -81691 158 -81679
rect -158 -81921 -100 -81909
rect -158 -82497 -146 -81921
rect -112 -82497 -100 -81921
rect -158 -82509 -100 -82497
rect 100 -81921 158 -81909
rect 100 -82497 112 -81921
rect 146 -82497 158 -81921
rect 100 -82509 158 -82497
rect -158 -82739 -100 -82727
rect -158 -83315 -146 -82739
rect -112 -83315 -100 -82739
rect -158 -83327 -100 -83315
rect 100 -82739 158 -82727
rect 100 -83315 112 -82739
rect 146 -83315 158 -82739
rect 100 -83327 158 -83315
rect -158 -83557 -100 -83545
rect -158 -84133 -146 -83557
rect -112 -84133 -100 -83557
rect -158 -84145 -100 -84133
rect 100 -83557 158 -83545
rect 100 -84133 112 -83557
rect 146 -84133 158 -83557
rect 100 -84145 158 -84133
rect -158 -84375 -100 -84363
rect -158 -84951 -146 -84375
rect -112 -84951 -100 -84375
rect -158 -84963 -100 -84951
rect 100 -84375 158 -84363
rect 100 -84951 112 -84375
rect 146 -84951 158 -84375
rect 100 -84963 158 -84951
rect -158 -85193 -100 -85181
rect -158 -85769 -146 -85193
rect -112 -85769 -100 -85193
rect -158 -85781 -100 -85769
rect 100 -85193 158 -85181
rect 100 -85769 112 -85193
rect 146 -85769 158 -85193
rect 100 -85781 158 -85769
rect -158 -86011 -100 -85999
rect -158 -86587 -146 -86011
rect -112 -86587 -100 -86011
rect -158 -86599 -100 -86587
rect 100 -86011 158 -85999
rect 100 -86587 112 -86011
rect 146 -86587 158 -86011
rect 100 -86599 158 -86587
rect -158 -86829 -100 -86817
rect -158 -87405 -146 -86829
rect -112 -87405 -100 -86829
rect -158 -87417 -100 -87405
rect 100 -86829 158 -86817
rect 100 -87405 112 -86829
rect 146 -87405 158 -86829
rect 100 -87417 158 -87405
rect -158 -87647 -100 -87635
rect -158 -88223 -146 -87647
rect -112 -88223 -100 -87647
rect -158 -88235 -100 -88223
rect 100 -87647 158 -87635
rect 100 -88223 112 -87647
rect 146 -88223 158 -87647
rect 100 -88235 158 -88223
rect -158 -88465 -100 -88453
rect -158 -89041 -146 -88465
rect -112 -89041 -100 -88465
rect -158 -89053 -100 -89041
rect 100 -88465 158 -88453
rect 100 -89041 112 -88465
rect 146 -89041 158 -88465
rect 100 -89053 158 -89041
rect -158 -89283 -100 -89271
rect -158 -89859 -146 -89283
rect -112 -89859 -100 -89283
rect -158 -89871 -100 -89859
rect 100 -89283 158 -89271
rect 100 -89859 112 -89283
rect 146 -89859 158 -89283
rect 100 -89871 158 -89859
rect -158 -90101 -100 -90089
rect -158 -90677 -146 -90101
rect -112 -90677 -100 -90101
rect -158 -90689 -100 -90677
rect 100 -90101 158 -90089
rect 100 -90677 112 -90101
rect 146 -90677 158 -90101
rect 100 -90689 158 -90677
rect -158 -90919 -100 -90907
rect -158 -91495 -146 -90919
rect -112 -91495 -100 -90919
rect -158 -91507 -100 -91495
rect 100 -90919 158 -90907
rect 100 -91495 112 -90919
rect 146 -91495 158 -90919
rect 100 -91507 158 -91495
rect -158 -91737 -100 -91725
rect -158 -92313 -146 -91737
rect -112 -92313 -100 -91737
rect -158 -92325 -100 -92313
rect 100 -91737 158 -91725
rect 100 -92313 112 -91737
rect 146 -92313 158 -91737
rect 100 -92325 158 -92313
rect -158 -92555 -100 -92543
rect -158 -93131 -146 -92555
rect -112 -93131 -100 -92555
rect -158 -93143 -100 -93131
rect 100 -92555 158 -92543
rect 100 -93131 112 -92555
rect 146 -93131 158 -92555
rect 100 -93143 158 -93131
rect -158 -93373 -100 -93361
rect -158 -93949 -146 -93373
rect -112 -93949 -100 -93373
rect -158 -93961 -100 -93949
rect 100 -93373 158 -93361
rect 100 -93949 112 -93373
rect 146 -93949 158 -93373
rect 100 -93961 158 -93949
rect -158 -94191 -100 -94179
rect -158 -94767 -146 -94191
rect -112 -94767 -100 -94191
rect -158 -94779 -100 -94767
rect 100 -94191 158 -94179
rect 100 -94767 112 -94191
rect 146 -94767 158 -94191
rect 100 -94779 158 -94767
rect -158 -95009 -100 -94997
rect -158 -95585 -146 -95009
rect -112 -95585 -100 -95009
rect -158 -95597 -100 -95585
rect 100 -95009 158 -94997
rect 100 -95585 112 -95009
rect 146 -95585 158 -95009
rect 100 -95597 158 -95585
rect -158 -95827 -100 -95815
rect -158 -96403 -146 -95827
rect -112 -96403 -100 -95827
rect -158 -96415 -100 -96403
rect 100 -95827 158 -95815
rect 100 -96403 112 -95827
rect 146 -96403 158 -95827
rect 100 -96415 158 -96403
rect -158 -96645 -100 -96633
rect -158 -97221 -146 -96645
rect -112 -97221 -100 -96645
rect -158 -97233 -100 -97221
rect 100 -96645 158 -96633
rect 100 -97221 112 -96645
rect 146 -97221 158 -96645
rect 100 -97233 158 -97221
rect -158 -97463 -100 -97451
rect -158 -98039 -146 -97463
rect -112 -98039 -100 -97463
rect -158 -98051 -100 -98039
rect 100 -97463 158 -97451
rect 100 -98039 112 -97463
rect 146 -98039 158 -97463
rect 100 -98051 158 -98039
rect -158 -98281 -100 -98269
rect -158 -98857 -146 -98281
rect -112 -98857 -100 -98281
rect -158 -98869 -100 -98857
rect 100 -98281 158 -98269
rect 100 -98857 112 -98281
rect 146 -98857 158 -98281
rect 100 -98869 158 -98857
rect -158 -99099 -100 -99087
rect -158 -99675 -146 -99099
rect -112 -99675 -100 -99099
rect -158 -99687 -100 -99675
rect 100 -99099 158 -99087
rect 100 -99675 112 -99099
rect 146 -99675 158 -99099
rect 100 -99687 158 -99675
rect -158 -99917 -100 -99905
rect -158 -100493 -146 -99917
rect -112 -100493 -100 -99917
rect -158 -100505 -100 -100493
rect 100 -99917 158 -99905
rect 100 -100493 112 -99917
rect 146 -100493 158 -99917
rect 100 -100505 158 -100493
rect -158 -100735 -100 -100723
rect -158 -101311 -146 -100735
rect -112 -101311 -100 -100735
rect -158 -101323 -100 -101311
rect 100 -100735 158 -100723
rect 100 -101311 112 -100735
rect 146 -101311 158 -100735
rect 100 -101323 158 -101311
rect -158 -101553 -100 -101541
rect -158 -102129 -146 -101553
rect -112 -102129 -100 -101553
rect -158 -102141 -100 -102129
rect 100 -101553 158 -101541
rect 100 -102129 112 -101553
rect 146 -102129 158 -101553
rect 100 -102141 158 -102129
rect -158 -102371 -100 -102359
rect -158 -102947 -146 -102371
rect -112 -102947 -100 -102371
rect -158 -102959 -100 -102947
rect 100 -102371 158 -102359
rect 100 -102947 112 -102371
rect 146 -102947 158 -102371
rect 100 -102959 158 -102947
rect -158 -103189 -100 -103177
rect -158 -103765 -146 -103189
rect -112 -103765 -100 -103189
rect -158 -103777 -100 -103765
rect 100 -103189 158 -103177
rect 100 -103765 112 -103189
rect 146 -103765 158 -103189
rect 100 -103777 158 -103765
rect -158 -104007 -100 -103995
rect -158 -104583 -146 -104007
rect -112 -104583 -100 -104007
rect -158 -104595 -100 -104583
rect 100 -104007 158 -103995
rect 100 -104583 112 -104007
rect 146 -104583 158 -104007
rect 100 -104595 158 -104583
<< mvndiffc >>
rect -146 104007 -112 104583
rect 112 104007 146 104583
rect -146 103189 -112 103765
rect 112 103189 146 103765
rect -146 102371 -112 102947
rect 112 102371 146 102947
rect -146 101553 -112 102129
rect 112 101553 146 102129
rect -146 100735 -112 101311
rect 112 100735 146 101311
rect -146 99917 -112 100493
rect 112 99917 146 100493
rect -146 99099 -112 99675
rect 112 99099 146 99675
rect -146 98281 -112 98857
rect 112 98281 146 98857
rect -146 97463 -112 98039
rect 112 97463 146 98039
rect -146 96645 -112 97221
rect 112 96645 146 97221
rect -146 95827 -112 96403
rect 112 95827 146 96403
rect -146 95009 -112 95585
rect 112 95009 146 95585
rect -146 94191 -112 94767
rect 112 94191 146 94767
rect -146 93373 -112 93949
rect 112 93373 146 93949
rect -146 92555 -112 93131
rect 112 92555 146 93131
rect -146 91737 -112 92313
rect 112 91737 146 92313
rect -146 90919 -112 91495
rect 112 90919 146 91495
rect -146 90101 -112 90677
rect 112 90101 146 90677
rect -146 89283 -112 89859
rect 112 89283 146 89859
rect -146 88465 -112 89041
rect 112 88465 146 89041
rect -146 87647 -112 88223
rect 112 87647 146 88223
rect -146 86829 -112 87405
rect 112 86829 146 87405
rect -146 86011 -112 86587
rect 112 86011 146 86587
rect -146 85193 -112 85769
rect 112 85193 146 85769
rect -146 84375 -112 84951
rect 112 84375 146 84951
rect -146 83557 -112 84133
rect 112 83557 146 84133
rect -146 82739 -112 83315
rect 112 82739 146 83315
rect -146 81921 -112 82497
rect 112 81921 146 82497
rect -146 81103 -112 81679
rect 112 81103 146 81679
rect -146 80285 -112 80861
rect 112 80285 146 80861
rect -146 79467 -112 80043
rect 112 79467 146 80043
rect -146 78649 -112 79225
rect 112 78649 146 79225
rect -146 77831 -112 78407
rect 112 77831 146 78407
rect -146 77013 -112 77589
rect 112 77013 146 77589
rect -146 76195 -112 76771
rect 112 76195 146 76771
rect -146 75377 -112 75953
rect 112 75377 146 75953
rect -146 74559 -112 75135
rect 112 74559 146 75135
rect -146 73741 -112 74317
rect 112 73741 146 74317
rect -146 72923 -112 73499
rect 112 72923 146 73499
rect -146 72105 -112 72681
rect 112 72105 146 72681
rect -146 71287 -112 71863
rect 112 71287 146 71863
rect -146 70469 -112 71045
rect 112 70469 146 71045
rect -146 69651 -112 70227
rect 112 69651 146 70227
rect -146 68833 -112 69409
rect 112 68833 146 69409
rect -146 68015 -112 68591
rect 112 68015 146 68591
rect -146 67197 -112 67773
rect 112 67197 146 67773
rect -146 66379 -112 66955
rect 112 66379 146 66955
rect -146 65561 -112 66137
rect 112 65561 146 66137
rect -146 64743 -112 65319
rect 112 64743 146 65319
rect -146 63925 -112 64501
rect 112 63925 146 64501
rect -146 63107 -112 63683
rect 112 63107 146 63683
rect -146 62289 -112 62865
rect 112 62289 146 62865
rect -146 61471 -112 62047
rect 112 61471 146 62047
rect -146 60653 -112 61229
rect 112 60653 146 61229
rect -146 59835 -112 60411
rect 112 59835 146 60411
rect -146 59017 -112 59593
rect 112 59017 146 59593
rect -146 58199 -112 58775
rect 112 58199 146 58775
rect -146 57381 -112 57957
rect 112 57381 146 57957
rect -146 56563 -112 57139
rect 112 56563 146 57139
rect -146 55745 -112 56321
rect 112 55745 146 56321
rect -146 54927 -112 55503
rect 112 54927 146 55503
rect -146 54109 -112 54685
rect 112 54109 146 54685
rect -146 53291 -112 53867
rect 112 53291 146 53867
rect -146 52473 -112 53049
rect 112 52473 146 53049
rect -146 51655 -112 52231
rect 112 51655 146 52231
rect -146 50837 -112 51413
rect 112 50837 146 51413
rect -146 50019 -112 50595
rect 112 50019 146 50595
rect -146 49201 -112 49777
rect 112 49201 146 49777
rect -146 48383 -112 48959
rect 112 48383 146 48959
rect -146 47565 -112 48141
rect 112 47565 146 48141
rect -146 46747 -112 47323
rect 112 46747 146 47323
rect -146 45929 -112 46505
rect 112 45929 146 46505
rect -146 45111 -112 45687
rect 112 45111 146 45687
rect -146 44293 -112 44869
rect 112 44293 146 44869
rect -146 43475 -112 44051
rect 112 43475 146 44051
rect -146 42657 -112 43233
rect 112 42657 146 43233
rect -146 41839 -112 42415
rect 112 41839 146 42415
rect -146 41021 -112 41597
rect 112 41021 146 41597
rect -146 40203 -112 40779
rect 112 40203 146 40779
rect -146 39385 -112 39961
rect 112 39385 146 39961
rect -146 38567 -112 39143
rect 112 38567 146 39143
rect -146 37749 -112 38325
rect 112 37749 146 38325
rect -146 36931 -112 37507
rect 112 36931 146 37507
rect -146 36113 -112 36689
rect 112 36113 146 36689
rect -146 35295 -112 35871
rect 112 35295 146 35871
rect -146 34477 -112 35053
rect 112 34477 146 35053
rect -146 33659 -112 34235
rect 112 33659 146 34235
rect -146 32841 -112 33417
rect 112 32841 146 33417
rect -146 32023 -112 32599
rect 112 32023 146 32599
rect -146 31205 -112 31781
rect 112 31205 146 31781
rect -146 30387 -112 30963
rect 112 30387 146 30963
rect -146 29569 -112 30145
rect 112 29569 146 30145
rect -146 28751 -112 29327
rect 112 28751 146 29327
rect -146 27933 -112 28509
rect 112 27933 146 28509
rect -146 27115 -112 27691
rect 112 27115 146 27691
rect -146 26297 -112 26873
rect 112 26297 146 26873
rect -146 25479 -112 26055
rect 112 25479 146 26055
rect -146 24661 -112 25237
rect 112 24661 146 25237
rect -146 23843 -112 24419
rect 112 23843 146 24419
rect -146 23025 -112 23601
rect 112 23025 146 23601
rect -146 22207 -112 22783
rect 112 22207 146 22783
rect -146 21389 -112 21965
rect 112 21389 146 21965
rect -146 20571 -112 21147
rect 112 20571 146 21147
rect -146 19753 -112 20329
rect 112 19753 146 20329
rect -146 18935 -112 19511
rect 112 18935 146 19511
rect -146 18117 -112 18693
rect 112 18117 146 18693
rect -146 17299 -112 17875
rect 112 17299 146 17875
rect -146 16481 -112 17057
rect 112 16481 146 17057
rect -146 15663 -112 16239
rect 112 15663 146 16239
rect -146 14845 -112 15421
rect 112 14845 146 15421
rect -146 14027 -112 14603
rect 112 14027 146 14603
rect -146 13209 -112 13785
rect 112 13209 146 13785
rect -146 12391 -112 12967
rect 112 12391 146 12967
rect -146 11573 -112 12149
rect 112 11573 146 12149
rect -146 10755 -112 11331
rect 112 10755 146 11331
rect -146 9937 -112 10513
rect 112 9937 146 10513
rect -146 9119 -112 9695
rect 112 9119 146 9695
rect -146 8301 -112 8877
rect 112 8301 146 8877
rect -146 7483 -112 8059
rect 112 7483 146 8059
rect -146 6665 -112 7241
rect 112 6665 146 7241
rect -146 5847 -112 6423
rect 112 5847 146 6423
rect -146 5029 -112 5605
rect 112 5029 146 5605
rect -146 4211 -112 4787
rect 112 4211 146 4787
rect -146 3393 -112 3969
rect 112 3393 146 3969
rect -146 2575 -112 3151
rect 112 2575 146 3151
rect -146 1757 -112 2333
rect 112 1757 146 2333
rect -146 939 -112 1515
rect 112 939 146 1515
rect -146 121 -112 697
rect 112 121 146 697
rect -146 -697 -112 -121
rect 112 -697 146 -121
rect -146 -1515 -112 -939
rect 112 -1515 146 -939
rect -146 -2333 -112 -1757
rect 112 -2333 146 -1757
rect -146 -3151 -112 -2575
rect 112 -3151 146 -2575
rect -146 -3969 -112 -3393
rect 112 -3969 146 -3393
rect -146 -4787 -112 -4211
rect 112 -4787 146 -4211
rect -146 -5605 -112 -5029
rect 112 -5605 146 -5029
rect -146 -6423 -112 -5847
rect 112 -6423 146 -5847
rect -146 -7241 -112 -6665
rect 112 -7241 146 -6665
rect -146 -8059 -112 -7483
rect 112 -8059 146 -7483
rect -146 -8877 -112 -8301
rect 112 -8877 146 -8301
rect -146 -9695 -112 -9119
rect 112 -9695 146 -9119
rect -146 -10513 -112 -9937
rect 112 -10513 146 -9937
rect -146 -11331 -112 -10755
rect 112 -11331 146 -10755
rect -146 -12149 -112 -11573
rect 112 -12149 146 -11573
rect -146 -12967 -112 -12391
rect 112 -12967 146 -12391
rect -146 -13785 -112 -13209
rect 112 -13785 146 -13209
rect -146 -14603 -112 -14027
rect 112 -14603 146 -14027
rect -146 -15421 -112 -14845
rect 112 -15421 146 -14845
rect -146 -16239 -112 -15663
rect 112 -16239 146 -15663
rect -146 -17057 -112 -16481
rect 112 -17057 146 -16481
rect -146 -17875 -112 -17299
rect 112 -17875 146 -17299
rect -146 -18693 -112 -18117
rect 112 -18693 146 -18117
rect -146 -19511 -112 -18935
rect 112 -19511 146 -18935
rect -146 -20329 -112 -19753
rect 112 -20329 146 -19753
rect -146 -21147 -112 -20571
rect 112 -21147 146 -20571
rect -146 -21965 -112 -21389
rect 112 -21965 146 -21389
rect -146 -22783 -112 -22207
rect 112 -22783 146 -22207
rect -146 -23601 -112 -23025
rect 112 -23601 146 -23025
rect -146 -24419 -112 -23843
rect 112 -24419 146 -23843
rect -146 -25237 -112 -24661
rect 112 -25237 146 -24661
rect -146 -26055 -112 -25479
rect 112 -26055 146 -25479
rect -146 -26873 -112 -26297
rect 112 -26873 146 -26297
rect -146 -27691 -112 -27115
rect 112 -27691 146 -27115
rect -146 -28509 -112 -27933
rect 112 -28509 146 -27933
rect -146 -29327 -112 -28751
rect 112 -29327 146 -28751
rect -146 -30145 -112 -29569
rect 112 -30145 146 -29569
rect -146 -30963 -112 -30387
rect 112 -30963 146 -30387
rect -146 -31781 -112 -31205
rect 112 -31781 146 -31205
rect -146 -32599 -112 -32023
rect 112 -32599 146 -32023
rect -146 -33417 -112 -32841
rect 112 -33417 146 -32841
rect -146 -34235 -112 -33659
rect 112 -34235 146 -33659
rect -146 -35053 -112 -34477
rect 112 -35053 146 -34477
rect -146 -35871 -112 -35295
rect 112 -35871 146 -35295
rect -146 -36689 -112 -36113
rect 112 -36689 146 -36113
rect -146 -37507 -112 -36931
rect 112 -37507 146 -36931
rect -146 -38325 -112 -37749
rect 112 -38325 146 -37749
rect -146 -39143 -112 -38567
rect 112 -39143 146 -38567
rect -146 -39961 -112 -39385
rect 112 -39961 146 -39385
rect -146 -40779 -112 -40203
rect 112 -40779 146 -40203
rect -146 -41597 -112 -41021
rect 112 -41597 146 -41021
rect -146 -42415 -112 -41839
rect 112 -42415 146 -41839
rect -146 -43233 -112 -42657
rect 112 -43233 146 -42657
rect -146 -44051 -112 -43475
rect 112 -44051 146 -43475
rect -146 -44869 -112 -44293
rect 112 -44869 146 -44293
rect -146 -45687 -112 -45111
rect 112 -45687 146 -45111
rect -146 -46505 -112 -45929
rect 112 -46505 146 -45929
rect -146 -47323 -112 -46747
rect 112 -47323 146 -46747
rect -146 -48141 -112 -47565
rect 112 -48141 146 -47565
rect -146 -48959 -112 -48383
rect 112 -48959 146 -48383
rect -146 -49777 -112 -49201
rect 112 -49777 146 -49201
rect -146 -50595 -112 -50019
rect 112 -50595 146 -50019
rect -146 -51413 -112 -50837
rect 112 -51413 146 -50837
rect -146 -52231 -112 -51655
rect 112 -52231 146 -51655
rect -146 -53049 -112 -52473
rect 112 -53049 146 -52473
rect -146 -53867 -112 -53291
rect 112 -53867 146 -53291
rect -146 -54685 -112 -54109
rect 112 -54685 146 -54109
rect -146 -55503 -112 -54927
rect 112 -55503 146 -54927
rect -146 -56321 -112 -55745
rect 112 -56321 146 -55745
rect -146 -57139 -112 -56563
rect 112 -57139 146 -56563
rect -146 -57957 -112 -57381
rect 112 -57957 146 -57381
rect -146 -58775 -112 -58199
rect 112 -58775 146 -58199
rect -146 -59593 -112 -59017
rect 112 -59593 146 -59017
rect -146 -60411 -112 -59835
rect 112 -60411 146 -59835
rect -146 -61229 -112 -60653
rect 112 -61229 146 -60653
rect -146 -62047 -112 -61471
rect 112 -62047 146 -61471
rect -146 -62865 -112 -62289
rect 112 -62865 146 -62289
rect -146 -63683 -112 -63107
rect 112 -63683 146 -63107
rect -146 -64501 -112 -63925
rect 112 -64501 146 -63925
rect -146 -65319 -112 -64743
rect 112 -65319 146 -64743
rect -146 -66137 -112 -65561
rect 112 -66137 146 -65561
rect -146 -66955 -112 -66379
rect 112 -66955 146 -66379
rect -146 -67773 -112 -67197
rect 112 -67773 146 -67197
rect -146 -68591 -112 -68015
rect 112 -68591 146 -68015
rect -146 -69409 -112 -68833
rect 112 -69409 146 -68833
rect -146 -70227 -112 -69651
rect 112 -70227 146 -69651
rect -146 -71045 -112 -70469
rect 112 -71045 146 -70469
rect -146 -71863 -112 -71287
rect 112 -71863 146 -71287
rect -146 -72681 -112 -72105
rect 112 -72681 146 -72105
rect -146 -73499 -112 -72923
rect 112 -73499 146 -72923
rect -146 -74317 -112 -73741
rect 112 -74317 146 -73741
rect -146 -75135 -112 -74559
rect 112 -75135 146 -74559
rect -146 -75953 -112 -75377
rect 112 -75953 146 -75377
rect -146 -76771 -112 -76195
rect 112 -76771 146 -76195
rect -146 -77589 -112 -77013
rect 112 -77589 146 -77013
rect -146 -78407 -112 -77831
rect 112 -78407 146 -77831
rect -146 -79225 -112 -78649
rect 112 -79225 146 -78649
rect -146 -80043 -112 -79467
rect 112 -80043 146 -79467
rect -146 -80861 -112 -80285
rect 112 -80861 146 -80285
rect -146 -81679 -112 -81103
rect 112 -81679 146 -81103
rect -146 -82497 -112 -81921
rect 112 -82497 146 -81921
rect -146 -83315 -112 -82739
rect 112 -83315 146 -82739
rect -146 -84133 -112 -83557
rect 112 -84133 146 -83557
rect -146 -84951 -112 -84375
rect 112 -84951 146 -84375
rect -146 -85769 -112 -85193
rect 112 -85769 146 -85193
rect -146 -86587 -112 -86011
rect 112 -86587 146 -86011
rect -146 -87405 -112 -86829
rect 112 -87405 146 -86829
rect -146 -88223 -112 -87647
rect 112 -88223 146 -87647
rect -146 -89041 -112 -88465
rect 112 -89041 146 -88465
rect -146 -89859 -112 -89283
rect 112 -89859 146 -89283
rect -146 -90677 -112 -90101
rect 112 -90677 146 -90101
rect -146 -91495 -112 -90919
rect 112 -91495 146 -90919
rect -146 -92313 -112 -91737
rect 112 -92313 146 -91737
rect -146 -93131 -112 -92555
rect 112 -93131 146 -92555
rect -146 -93949 -112 -93373
rect 112 -93949 146 -93373
rect -146 -94767 -112 -94191
rect 112 -94767 146 -94191
rect -146 -95585 -112 -95009
rect 112 -95585 146 -95009
rect -146 -96403 -112 -95827
rect 112 -96403 146 -95827
rect -146 -97221 -112 -96645
rect 112 -97221 146 -96645
rect -146 -98039 -112 -97463
rect 112 -98039 146 -97463
rect -146 -98857 -112 -98281
rect 112 -98857 146 -98281
rect -146 -99675 -112 -99099
rect 112 -99675 146 -99099
rect -146 -100493 -112 -99917
rect 112 -100493 146 -99917
rect -146 -101311 -112 -100735
rect 112 -101311 146 -100735
rect -146 -102129 -112 -101553
rect 112 -102129 146 -101553
rect -146 -102947 -112 -102371
rect 112 -102947 146 -102371
rect -146 -103765 -112 -103189
rect 112 -103765 146 -103189
rect -146 -104583 -112 -104007
rect 112 -104583 146 -104007
<< mvpsubdiff >>
rect -292 104805 292 104817
rect -292 104771 -184 104805
rect 184 104771 292 104805
rect -292 104759 292 104771
rect -292 104709 -234 104759
rect -292 -104709 -280 104709
rect -246 -104709 -234 104709
rect 234 104709 292 104759
rect -292 -104759 -234 -104709
rect 234 -104709 246 104709
rect 280 -104709 292 104709
rect 234 -104759 292 -104709
rect -292 -104771 292 -104759
rect -292 -104805 -184 -104771
rect 184 -104805 292 -104771
rect -292 -104817 292 -104805
<< mvpsubdiffcont >>
rect -184 104771 184 104805
rect -280 -104709 -246 104709
rect 246 -104709 280 104709
rect -184 -104805 184 -104771
<< poly >>
rect -100 104667 100 104683
rect -100 104633 -84 104667
rect 84 104633 100 104667
rect -100 104595 100 104633
rect -100 103957 100 103995
rect -100 103923 -84 103957
rect 84 103923 100 103957
rect -100 103907 100 103923
rect -100 103849 100 103865
rect -100 103815 -84 103849
rect 84 103815 100 103849
rect -100 103777 100 103815
rect -100 103139 100 103177
rect -100 103105 -84 103139
rect 84 103105 100 103139
rect -100 103089 100 103105
rect -100 103031 100 103047
rect -100 102997 -84 103031
rect 84 102997 100 103031
rect -100 102959 100 102997
rect -100 102321 100 102359
rect -100 102287 -84 102321
rect 84 102287 100 102321
rect -100 102271 100 102287
rect -100 102213 100 102229
rect -100 102179 -84 102213
rect 84 102179 100 102213
rect -100 102141 100 102179
rect -100 101503 100 101541
rect -100 101469 -84 101503
rect 84 101469 100 101503
rect -100 101453 100 101469
rect -100 101395 100 101411
rect -100 101361 -84 101395
rect 84 101361 100 101395
rect -100 101323 100 101361
rect -100 100685 100 100723
rect -100 100651 -84 100685
rect 84 100651 100 100685
rect -100 100635 100 100651
rect -100 100577 100 100593
rect -100 100543 -84 100577
rect 84 100543 100 100577
rect -100 100505 100 100543
rect -100 99867 100 99905
rect -100 99833 -84 99867
rect 84 99833 100 99867
rect -100 99817 100 99833
rect -100 99759 100 99775
rect -100 99725 -84 99759
rect 84 99725 100 99759
rect -100 99687 100 99725
rect -100 99049 100 99087
rect -100 99015 -84 99049
rect 84 99015 100 99049
rect -100 98999 100 99015
rect -100 98941 100 98957
rect -100 98907 -84 98941
rect 84 98907 100 98941
rect -100 98869 100 98907
rect -100 98231 100 98269
rect -100 98197 -84 98231
rect 84 98197 100 98231
rect -100 98181 100 98197
rect -100 98123 100 98139
rect -100 98089 -84 98123
rect 84 98089 100 98123
rect -100 98051 100 98089
rect -100 97413 100 97451
rect -100 97379 -84 97413
rect 84 97379 100 97413
rect -100 97363 100 97379
rect -100 97305 100 97321
rect -100 97271 -84 97305
rect 84 97271 100 97305
rect -100 97233 100 97271
rect -100 96595 100 96633
rect -100 96561 -84 96595
rect 84 96561 100 96595
rect -100 96545 100 96561
rect -100 96487 100 96503
rect -100 96453 -84 96487
rect 84 96453 100 96487
rect -100 96415 100 96453
rect -100 95777 100 95815
rect -100 95743 -84 95777
rect 84 95743 100 95777
rect -100 95727 100 95743
rect -100 95669 100 95685
rect -100 95635 -84 95669
rect 84 95635 100 95669
rect -100 95597 100 95635
rect -100 94959 100 94997
rect -100 94925 -84 94959
rect 84 94925 100 94959
rect -100 94909 100 94925
rect -100 94851 100 94867
rect -100 94817 -84 94851
rect 84 94817 100 94851
rect -100 94779 100 94817
rect -100 94141 100 94179
rect -100 94107 -84 94141
rect 84 94107 100 94141
rect -100 94091 100 94107
rect -100 94033 100 94049
rect -100 93999 -84 94033
rect 84 93999 100 94033
rect -100 93961 100 93999
rect -100 93323 100 93361
rect -100 93289 -84 93323
rect 84 93289 100 93323
rect -100 93273 100 93289
rect -100 93215 100 93231
rect -100 93181 -84 93215
rect 84 93181 100 93215
rect -100 93143 100 93181
rect -100 92505 100 92543
rect -100 92471 -84 92505
rect 84 92471 100 92505
rect -100 92455 100 92471
rect -100 92397 100 92413
rect -100 92363 -84 92397
rect 84 92363 100 92397
rect -100 92325 100 92363
rect -100 91687 100 91725
rect -100 91653 -84 91687
rect 84 91653 100 91687
rect -100 91637 100 91653
rect -100 91579 100 91595
rect -100 91545 -84 91579
rect 84 91545 100 91579
rect -100 91507 100 91545
rect -100 90869 100 90907
rect -100 90835 -84 90869
rect 84 90835 100 90869
rect -100 90819 100 90835
rect -100 90761 100 90777
rect -100 90727 -84 90761
rect 84 90727 100 90761
rect -100 90689 100 90727
rect -100 90051 100 90089
rect -100 90017 -84 90051
rect 84 90017 100 90051
rect -100 90001 100 90017
rect -100 89943 100 89959
rect -100 89909 -84 89943
rect 84 89909 100 89943
rect -100 89871 100 89909
rect -100 89233 100 89271
rect -100 89199 -84 89233
rect 84 89199 100 89233
rect -100 89183 100 89199
rect -100 89125 100 89141
rect -100 89091 -84 89125
rect 84 89091 100 89125
rect -100 89053 100 89091
rect -100 88415 100 88453
rect -100 88381 -84 88415
rect 84 88381 100 88415
rect -100 88365 100 88381
rect -100 88307 100 88323
rect -100 88273 -84 88307
rect 84 88273 100 88307
rect -100 88235 100 88273
rect -100 87597 100 87635
rect -100 87563 -84 87597
rect 84 87563 100 87597
rect -100 87547 100 87563
rect -100 87489 100 87505
rect -100 87455 -84 87489
rect 84 87455 100 87489
rect -100 87417 100 87455
rect -100 86779 100 86817
rect -100 86745 -84 86779
rect 84 86745 100 86779
rect -100 86729 100 86745
rect -100 86671 100 86687
rect -100 86637 -84 86671
rect 84 86637 100 86671
rect -100 86599 100 86637
rect -100 85961 100 85999
rect -100 85927 -84 85961
rect 84 85927 100 85961
rect -100 85911 100 85927
rect -100 85853 100 85869
rect -100 85819 -84 85853
rect 84 85819 100 85853
rect -100 85781 100 85819
rect -100 85143 100 85181
rect -100 85109 -84 85143
rect 84 85109 100 85143
rect -100 85093 100 85109
rect -100 85035 100 85051
rect -100 85001 -84 85035
rect 84 85001 100 85035
rect -100 84963 100 85001
rect -100 84325 100 84363
rect -100 84291 -84 84325
rect 84 84291 100 84325
rect -100 84275 100 84291
rect -100 84217 100 84233
rect -100 84183 -84 84217
rect 84 84183 100 84217
rect -100 84145 100 84183
rect -100 83507 100 83545
rect -100 83473 -84 83507
rect 84 83473 100 83507
rect -100 83457 100 83473
rect -100 83399 100 83415
rect -100 83365 -84 83399
rect 84 83365 100 83399
rect -100 83327 100 83365
rect -100 82689 100 82727
rect -100 82655 -84 82689
rect 84 82655 100 82689
rect -100 82639 100 82655
rect -100 82581 100 82597
rect -100 82547 -84 82581
rect 84 82547 100 82581
rect -100 82509 100 82547
rect -100 81871 100 81909
rect -100 81837 -84 81871
rect 84 81837 100 81871
rect -100 81821 100 81837
rect -100 81763 100 81779
rect -100 81729 -84 81763
rect 84 81729 100 81763
rect -100 81691 100 81729
rect -100 81053 100 81091
rect -100 81019 -84 81053
rect 84 81019 100 81053
rect -100 81003 100 81019
rect -100 80945 100 80961
rect -100 80911 -84 80945
rect 84 80911 100 80945
rect -100 80873 100 80911
rect -100 80235 100 80273
rect -100 80201 -84 80235
rect 84 80201 100 80235
rect -100 80185 100 80201
rect -100 80127 100 80143
rect -100 80093 -84 80127
rect 84 80093 100 80127
rect -100 80055 100 80093
rect -100 79417 100 79455
rect -100 79383 -84 79417
rect 84 79383 100 79417
rect -100 79367 100 79383
rect -100 79309 100 79325
rect -100 79275 -84 79309
rect 84 79275 100 79309
rect -100 79237 100 79275
rect -100 78599 100 78637
rect -100 78565 -84 78599
rect 84 78565 100 78599
rect -100 78549 100 78565
rect -100 78491 100 78507
rect -100 78457 -84 78491
rect 84 78457 100 78491
rect -100 78419 100 78457
rect -100 77781 100 77819
rect -100 77747 -84 77781
rect 84 77747 100 77781
rect -100 77731 100 77747
rect -100 77673 100 77689
rect -100 77639 -84 77673
rect 84 77639 100 77673
rect -100 77601 100 77639
rect -100 76963 100 77001
rect -100 76929 -84 76963
rect 84 76929 100 76963
rect -100 76913 100 76929
rect -100 76855 100 76871
rect -100 76821 -84 76855
rect 84 76821 100 76855
rect -100 76783 100 76821
rect -100 76145 100 76183
rect -100 76111 -84 76145
rect 84 76111 100 76145
rect -100 76095 100 76111
rect -100 76037 100 76053
rect -100 76003 -84 76037
rect 84 76003 100 76037
rect -100 75965 100 76003
rect -100 75327 100 75365
rect -100 75293 -84 75327
rect 84 75293 100 75327
rect -100 75277 100 75293
rect -100 75219 100 75235
rect -100 75185 -84 75219
rect 84 75185 100 75219
rect -100 75147 100 75185
rect -100 74509 100 74547
rect -100 74475 -84 74509
rect 84 74475 100 74509
rect -100 74459 100 74475
rect -100 74401 100 74417
rect -100 74367 -84 74401
rect 84 74367 100 74401
rect -100 74329 100 74367
rect -100 73691 100 73729
rect -100 73657 -84 73691
rect 84 73657 100 73691
rect -100 73641 100 73657
rect -100 73583 100 73599
rect -100 73549 -84 73583
rect 84 73549 100 73583
rect -100 73511 100 73549
rect -100 72873 100 72911
rect -100 72839 -84 72873
rect 84 72839 100 72873
rect -100 72823 100 72839
rect -100 72765 100 72781
rect -100 72731 -84 72765
rect 84 72731 100 72765
rect -100 72693 100 72731
rect -100 72055 100 72093
rect -100 72021 -84 72055
rect 84 72021 100 72055
rect -100 72005 100 72021
rect -100 71947 100 71963
rect -100 71913 -84 71947
rect 84 71913 100 71947
rect -100 71875 100 71913
rect -100 71237 100 71275
rect -100 71203 -84 71237
rect 84 71203 100 71237
rect -100 71187 100 71203
rect -100 71129 100 71145
rect -100 71095 -84 71129
rect 84 71095 100 71129
rect -100 71057 100 71095
rect -100 70419 100 70457
rect -100 70385 -84 70419
rect 84 70385 100 70419
rect -100 70369 100 70385
rect -100 70311 100 70327
rect -100 70277 -84 70311
rect 84 70277 100 70311
rect -100 70239 100 70277
rect -100 69601 100 69639
rect -100 69567 -84 69601
rect 84 69567 100 69601
rect -100 69551 100 69567
rect -100 69493 100 69509
rect -100 69459 -84 69493
rect 84 69459 100 69493
rect -100 69421 100 69459
rect -100 68783 100 68821
rect -100 68749 -84 68783
rect 84 68749 100 68783
rect -100 68733 100 68749
rect -100 68675 100 68691
rect -100 68641 -84 68675
rect 84 68641 100 68675
rect -100 68603 100 68641
rect -100 67965 100 68003
rect -100 67931 -84 67965
rect 84 67931 100 67965
rect -100 67915 100 67931
rect -100 67857 100 67873
rect -100 67823 -84 67857
rect 84 67823 100 67857
rect -100 67785 100 67823
rect -100 67147 100 67185
rect -100 67113 -84 67147
rect 84 67113 100 67147
rect -100 67097 100 67113
rect -100 67039 100 67055
rect -100 67005 -84 67039
rect 84 67005 100 67039
rect -100 66967 100 67005
rect -100 66329 100 66367
rect -100 66295 -84 66329
rect 84 66295 100 66329
rect -100 66279 100 66295
rect -100 66221 100 66237
rect -100 66187 -84 66221
rect 84 66187 100 66221
rect -100 66149 100 66187
rect -100 65511 100 65549
rect -100 65477 -84 65511
rect 84 65477 100 65511
rect -100 65461 100 65477
rect -100 65403 100 65419
rect -100 65369 -84 65403
rect 84 65369 100 65403
rect -100 65331 100 65369
rect -100 64693 100 64731
rect -100 64659 -84 64693
rect 84 64659 100 64693
rect -100 64643 100 64659
rect -100 64585 100 64601
rect -100 64551 -84 64585
rect 84 64551 100 64585
rect -100 64513 100 64551
rect -100 63875 100 63913
rect -100 63841 -84 63875
rect 84 63841 100 63875
rect -100 63825 100 63841
rect -100 63767 100 63783
rect -100 63733 -84 63767
rect 84 63733 100 63767
rect -100 63695 100 63733
rect -100 63057 100 63095
rect -100 63023 -84 63057
rect 84 63023 100 63057
rect -100 63007 100 63023
rect -100 62949 100 62965
rect -100 62915 -84 62949
rect 84 62915 100 62949
rect -100 62877 100 62915
rect -100 62239 100 62277
rect -100 62205 -84 62239
rect 84 62205 100 62239
rect -100 62189 100 62205
rect -100 62131 100 62147
rect -100 62097 -84 62131
rect 84 62097 100 62131
rect -100 62059 100 62097
rect -100 61421 100 61459
rect -100 61387 -84 61421
rect 84 61387 100 61421
rect -100 61371 100 61387
rect -100 61313 100 61329
rect -100 61279 -84 61313
rect 84 61279 100 61313
rect -100 61241 100 61279
rect -100 60603 100 60641
rect -100 60569 -84 60603
rect 84 60569 100 60603
rect -100 60553 100 60569
rect -100 60495 100 60511
rect -100 60461 -84 60495
rect 84 60461 100 60495
rect -100 60423 100 60461
rect -100 59785 100 59823
rect -100 59751 -84 59785
rect 84 59751 100 59785
rect -100 59735 100 59751
rect -100 59677 100 59693
rect -100 59643 -84 59677
rect 84 59643 100 59677
rect -100 59605 100 59643
rect -100 58967 100 59005
rect -100 58933 -84 58967
rect 84 58933 100 58967
rect -100 58917 100 58933
rect -100 58859 100 58875
rect -100 58825 -84 58859
rect 84 58825 100 58859
rect -100 58787 100 58825
rect -100 58149 100 58187
rect -100 58115 -84 58149
rect 84 58115 100 58149
rect -100 58099 100 58115
rect -100 58041 100 58057
rect -100 58007 -84 58041
rect 84 58007 100 58041
rect -100 57969 100 58007
rect -100 57331 100 57369
rect -100 57297 -84 57331
rect 84 57297 100 57331
rect -100 57281 100 57297
rect -100 57223 100 57239
rect -100 57189 -84 57223
rect 84 57189 100 57223
rect -100 57151 100 57189
rect -100 56513 100 56551
rect -100 56479 -84 56513
rect 84 56479 100 56513
rect -100 56463 100 56479
rect -100 56405 100 56421
rect -100 56371 -84 56405
rect 84 56371 100 56405
rect -100 56333 100 56371
rect -100 55695 100 55733
rect -100 55661 -84 55695
rect 84 55661 100 55695
rect -100 55645 100 55661
rect -100 55587 100 55603
rect -100 55553 -84 55587
rect 84 55553 100 55587
rect -100 55515 100 55553
rect -100 54877 100 54915
rect -100 54843 -84 54877
rect 84 54843 100 54877
rect -100 54827 100 54843
rect -100 54769 100 54785
rect -100 54735 -84 54769
rect 84 54735 100 54769
rect -100 54697 100 54735
rect -100 54059 100 54097
rect -100 54025 -84 54059
rect 84 54025 100 54059
rect -100 54009 100 54025
rect -100 53951 100 53967
rect -100 53917 -84 53951
rect 84 53917 100 53951
rect -100 53879 100 53917
rect -100 53241 100 53279
rect -100 53207 -84 53241
rect 84 53207 100 53241
rect -100 53191 100 53207
rect -100 53133 100 53149
rect -100 53099 -84 53133
rect 84 53099 100 53133
rect -100 53061 100 53099
rect -100 52423 100 52461
rect -100 52389 -84 52423
rect 84 52389 100 52423
rect -100 52373 100 52389
rect -100 52315 100 52331
rect -100 52281 -84 52315
rect 84 52281 100 52315
rect -100 52243 100 52281
rect -100 51605 100 51643
rect -100 51571 -84 51605
rect 84 51571 100 51605
rect -100 51555 100 51571
rect -100 51497 100 51513
rect -100 51463 -84 51497
rect 84 51463 100 51497
rect -100 51425 100 51463
rect -100 50787 100 50825
rect -100 50753 -84 50787
rect 84 50753 100 50787
rect -100 50737 100 50753
rect -100 50679 100 50695
rect -100 50645 -84 50679
rect 84 50645 100 50679
rect -100 50607 100 50645
rect -100 49969 100 50007
rect -100 49935 -84 49969
rect 84 49935 100 49969
rect -100 49919 100 49935
rect -100 49861 100 49877
rect -100 49827 -84 49861
rect 84 49827 100 49861
rect -100 49789 100 49827
rect -100 49151 100 49189
rect -100 49117 -84 49151
rect 84 49117 100 49151
rect -100 49101 100 49117
rect -100 49043 100 49059
rect -100 49009 -84 49043
rect 84 49009 100 49043
rect -100 48971 100 49009
rect -100 48333 100 48371
rect -100 48299 -84 48333
rect 84 48299 100 48333
rect -100 48283 100 48299
rect -100 48225 100 48241
rect -100 48191 -84 48225
rect 84 48191 100 48225
rect -100 48153 100 48191
rect -100 47515 100 47553
rect -100 47481 -84 47515
rect 84 47481 100 47515
rect -100 47465 100 47481
rect -100 47407 100 47423
rect -100 47373 -84 47407
rect 84 47373 100 47407
rect -100 47335 100 47373
rect -100 46697 100 46735
rect -100 46663 -84 46697
rect 84 46663 100 46697
rect -100 46647 100 46663
rect -100 46589 100 46605
rect -100 46555 -84 46589
rect 84 46555 100 46589
rect -100 46517 100 46555
rect -100 45879 100 45917
rect -100 45845 -84 45879
rect 84 45845 100 45879
rect -100 45829 100 45845
rect -100 45771 100 45787
rect -100 45737 -84 45771
rect 84 45737 100 45771
rect -100 45699 100 45737
rect -100 45061 100 45099
rect -100 45027 -84 45061
rect 84 45027 100 45061
rect -100 45011 100 45027
rect -100 44953 100 44969
rect -100 44919 -84 44953
rect 84 44919 100 44953
rect -100 44881 100 44919
rect -100 44243 100 44281
rect -100 44209 -84 44243
rect 84 44209 100 44243
rect -100 44193 100 44209
rect -100 44135 100 44151
rect -100 44101 -84 44135
rect 84 44101 100 44135
rect -100 44063 100 44101
rect -100 43425 100 43463
rect -100 43391 -84 43425
rect 84 43391 100 43425
rect -100 43375 100 43391
rect -100 43317 100 43333
rect -100 43283 -84 43317
rect 84 43283 100 43317
rect -100 43245 100 43283
rect -100 42607 100 42645
rect -100 42573 -84 42607
rect 84 42573 100 42607
rect -100 42557 100 42573
rect -100 42499 100 42515
rect -100 42465 -84 42499
rect 84 42465 100 42499
rect -100 42427 100 42465
rect -100 41789 100 41827
rect -100 41755 -84 41789
rect 84 41755 100 41789
rect -100 41739 100 41755
rect -100 41681 100 41697
rect -100 41647 -84 41681
rect 84 41647 100 41681
rect -100 41609 100 41647
rect -100 40971 100 41009
rect -100 40937 -84 40971
rect 84 40937 100 40971
rect -100 40921 100 40937
rect -100 40863 100 40879
rect -100 40829 -84 40863
rect 84 40829 100 40863
rect -100 40791 100 40829
rect -100 40153 100 40191
rect -100 40119 -84 40153
rect 84 40119 100 40153
rect -100 40103 100 40119
rect -100 40045 100 40061
rect -100 40011 -84 40045
rect 84 40011 100 40045
rect -100 39973 100 40011
rect -100 39335 100 39373
rect -100 39301 -84 39335
rect 84 39301 100 39335
rect -100 39285 100 39301
rect -100 39227 100 39243
rect -100 39193 -84 39227
rect 84 39193 100 39227
rect -100 39155 100 39193
rect -100 38517 100 38555
rect -100 38483 -84 38517
rect 84 38483 100 38517
rect -100 38467 100 38483
rect -100 38409 100 38425
rect -100 38375 -84 38409
rect 84 38375 100 38409
rect -100 38337 100 38375
rect -100 37699 100 37737
rect -100 37665 -84 37699
rect 84 37665 100 37699
rect -100 37649 100 37665
rect -100 37591 100 37607
rect -100 37557 -84 37591
rect 84 37557 100 37591
rect -100 37519 100 37557
rect -100 36881 100 36919
rect -100 36847 -84 36881
rect 84 36847 100 36881
rect -100 36831 100 36847
rect -100 36773 100 36789
rect -100 36739 -84 36773
rect 84 36739 100 36773
rect -100 36701 100 36739
rect -100 36063 100 36101
rect -100 36029 -84 36063
rect 84 36029 100 36063
rect -100 36013 100 36029
rect -100 35955 100 35971
rect -100 35921 -84 35955
rect 84 35921 100 35955
rect -100 35883 100 35921
rect -100 35245 100 35283
rect -100 35211 -84 35245
rect 84 35211 100 35245
rect -100 35195 100 35211
rect -100 35137 100 35153
rect -100 35103 -84 35137
rect 84 35103 100 35137
rect -100 35065 100 35103
rect -100 34427 100 34465
rect -100 34393 -84 34427
rect 84 34393 100 34427
rect -100 34377 100 34393
rect -100 34319 100 34335
rect -100 34285 -84 34319
rect 84 34285 100 34319
rect -100 34247 100 34285
rect -100 33609 100 33647
rect -100 33575 -84 33609
rect 84 33575 100 33609
rect -100 33559 100 33575
rect -100 33501 100 33517
rect -100 33467 -84 33501
rect 84 33467 100 33501
rect -100 33429 100 33467
rect -100 32791 100 32829
rect -100 32757 -84 32791
rect 84 32757 100 32791
rect -100 32741 100 32757
rect -100 32683 100 32699
rect -100 32649 -84 32683
rect 84 32649 100 32683
rect -100 32611 100 32649
rect -100 31973 100 32011
rect -100 31939 -84 31973
rect 84 31939 100 31973
rect -100 31923 100 31939
rect -100 31865 100 31881
rect -100 31831 -84 31865
rect 84 31831 100 31865
rect -100 31793 100 31831
rect -100 31155 100 31193
rect -100 31121 -84 31155
rect 84 31121 100 31155
rect -100 31105 100 31121
rect -100 31047 100 31063
rect -100 31013 -84 31047
rect 84 31013 100 31047
rect -100 30975 100 31013
rect -100 30337 100 30375
rect -100 30303 -84 30337
rect 84 30303 100 30337
rect -100 30287 100 30303
rect -100 30229 100 30245
rect -100 30195 -84 30229
rect 84 30195 100 30229
rect -100 30157 100 30195
rect -100 29519 100 29557
rect -100 29485 -84 29519
rect 84 29485 100 29519
rect -100 29469 100 29485
rect -100 29411 100 29427
rect -100 29377 -84 29411
rect 84 29377 100 29411
rect -100 29339 100 29377
rect -100 28701 100 28739
rect -100 28667 -84 28701
rect 84 28667 100 28701
rect -100 28651 100 28667
rect -100 28593 100 28609
rect -100 28559 -84 28593
rect 84 28559 100 28593
rect -100 28521 100 28559
rect -100 27883 100 27921
rect -100 27849 -84 27883
rect 84 27849 100 27883
rect -100 27833 100 27849
rect -100 27775 100 27791
rect -100 27741 -84 27775
rect 84 27741 100 27775
rect -100 27703 100 27741
rect -100 27065 100 27103
rect -100 27031 -84 27065
rect 84 27031 100 27065
rect -100 27015 100 27031
rect -100 26957 100 26973
rect -100 26923 -84 26957
rect 84 26923 100 26957
rect -100 26885 100 26923
rect -100 26247 100 26285
rect -100 26213 -84 26247
rect 84 26213 100 26247
rect -100 26197 100 26213
rect -100 26139 100 26155
rect -100 26105 -84 26139
rect 84 26105 100 26139
rect -100 26067 100 26105
rect -100 25429 100 25467
rect -100 25395 -84 25429
rect 84 25395 100 25429
rect -100 25379 100 25395
rect -100 25321 100 25337
rect -100 25287 -84 25321
rect 84 25287 100 25321
rect -100 25249 100 25287
rect -100 24611 100 24649
rect -100 24577 -84 24611
rect 84 24577 100 24611
rect -100 24561 100 24577
rect -100 24503 100 24519
rect -100 24469 -84 24503
rect 84 24469 100 24503
rect -100 24431 100 24469
rect -100 23793 100 23831
rect -100 23759 -84 23793
rect 84 23759 100 23793
rect -100 23743 100 23759
rect -100 23685 100 23701
rect -100 23651 -84 23685
rect 84 23651 100 23685
rect -100 23613 100 23651
rect -100 22975 100 23013
rect -100 22941 -84 22975
rect 84 22941 100 22975
rect -100 22925 100 22941
rect -100 22867 100 22883
rect -100 22833 -84 22867
rect 84 22833 100 22867
rect -100 22795 100 22833
rect -100 22157 100 22195
rect -100 22123 -84 22157
rect 84 22123 100 22157
rect -100 22107 100 22123
rect -100 22049 100 22065
rect -100 22015 -84 22049
rect 84 22015 100 22049
rect -100 21977 100 22015
rect -100 21339 100 21377
rect -100 21305 -84 21339
rect 84 21305 100 21339
rect -100 21289 100 21305
rect -100 21231 100 21247
rect -100 21197 -84 21231
rect 84 21197 100 21231
rect -100 21159 100 21197
rect -100 20521 100 20559
rect -100 20487 -84 20521
rect 84 20487 100 20521
rect -100 20471 100 20487
rect -100 20413 100 20429
rect -100 20379 -84 20413
rect 84 20379 100 20413
rect -100 20341 100 20379
rect -100 19703 100 19741
rect -100 19669 -84 19703
rect 84 19669 100 19703
rect -100 19653 100 19669
rect -100 19595 100 19611
rect -100 19561 -84 19595
rect 84 19561 100 19595
rect -100 19523 100 19561
rect -100 18885 100 18923
rect -100 18851 -84 18885
rect 84 18851 100 18885
rect -100 18835 100 18851
rect -100 18777 100 18793
rect -100 18743 -84 18777
rect 84 18743 100 18777
rect -100 18705 100 18743
rect -100 18067 100 18105
rect -100 18033 -84 18067
rect 84 18033 100 18067
rect -100 18017 100 18033
rect -100 17959 100 17975
rect -100 17925 -84 17959
rect 84 17925 100 17959
rect -100 17887 100 17925
rect -100 17249 100 17287
rect -100 17215 -84 17249
rect 84 17215 100 17249
rect -100 17199 100 17215
rect -100 17141 100 17157
rect -100 17107 -84 17141
rect 84 17107 100 17141
rect -100 17069 100 17107
rect -100 16431 100 16469
rect -100 16397 -84 16431
rect 84 16397 100 16431
rect -100 16381 100 16397
rect -100 16323 100 16339
rect -100 16289 -84 16323
rect 84 16289 100 16323
rect -100 16251 100 16289
rect -100 15613 100 15651
rect -100 15579 -84 15613
rect 84 15579 100 15613
rect -100 15563 100 15579
rect -100 15505 100 15521
rect -100 15471 -84 15505
rect 84 15471 100 15505
rect -100 15433 100 15471
rect -100 14795 100 14833
rect -100 14761 -84 14795
rect 84 14761 100 14795
rect -100 14745 100 14761
rect -100 14687 100 14703
rect -100 14653 -84 14687
rect 84 14653 100 14687
rect -100 14615 100 14653
rect -100 13977 100 14015
rect -100 13943 -84 13977
rect 84 13943 100 13977
rect -100 13927 100 13943
rect -100 13869 100 13885
rect -100 13835 -84 13869
rect 84 13835 100 13869
rect -100 13797 100 13835
rect -100 13159 100 13197
rect -100 13125 -84 13159
rect 84 13125 100 13159
rect -100 13109 100 13125
rect -100 13051 100 13067
rect -100 13017 -84 13051
rect 84 13017 100 13051
rect -100 12979 100 13017
rect -100 12341 100 12379
rect -100 12307 -84 12341
rect 84 12307 100 12341
rect -100 12291 100 12307
rect -100 12233 100 12249
rect -100 12199 -84 12233
rect 84 12199 100 12233
rect -100 12161 100 12199
rect -100 11523 100 11561
rect -100 11489 -84 11523
rect 84 11489 100 11523
rect -100 11473 100 11489
rect -100 11415 100 11431
rect -100 11381 -84 11415
rect 84 11381 100 11415
rect -100 11343 100 11381
rect -100 10705 100 10743
rect -100 10671 -84 10705
rect 84 10671 100 10705
rect -100 10655 100 10671
rect -100 10597 100 10613
rect -100 10563 -84 10597
rect 84 10563 100 10597
rect -100 10525 100 10563
rect -100 9887 100 9925
rect -100 9853 -84 9887
rect 84 9853 100 9887
rect -100 9837 100 9853
rect -100 9779 100 9795
rect -100 9745 -84 9779
rect 84 9745 100 9779
rect -100 9707 100 9745
rect -100 9069 100 9107
rect -100 9035 -84 9069
rect 84 9035 100 9069
rect -100 9019 100 9035
rect -100 8961 100 8977
rect -100 8927 -84 8961
rect 84 8927 100 8961
rect -100 8889 100 8927
rect -100 8251 100 8289
rect -100 8217 -84 8251
rect 84 8217 100 8251
rect -100 8201 100 8217
rect -100 8143 100 8159
rect -100 8109 -84 8143
rect 84 8109 100 8143
rect -100 8071 100 8109
rect -100 7433 100 7471
rect -100 7399 -84 7433
rect 84 7399 100 7433
rect -100 7383 100 7399
rect -100 7325 100 7341
rect -100 7291 -84 7325
rect 84 7291 100 7325
rect -100 7253 100 7291
rect -100 6615 100 6653
rect -100 6581 -84 6615
rect 84 6581 100 6615
rect -100 6565 100 6581
rect -100 6507 100 6523
rect -100 6473 -84 6507
rect 84 6473 100 6507
rect -100 6435 100 6473
rect -100 5797 100 5835
rect -100 5763 -84 5797
rect 84 5763 100 5797
rect -100 5747 100 5763
rect -100 5689 100 5705
rect -100 5655 -84 5689
rect 84 5655 100 5689
rect -100 5617 100 5655
rect -100 4979 100 5017
rect -100 4945 -84 4979
rect 84 4945 100 4979
rect -100 4929 100 4945
rect -100 4871 100 4887
rect -100 4837 -84 4871
rect 84 4837 100 4871
rect -100 4799 100 4837
rect -100 4161 100 4199
rect -100 4127 -84 4161
rect 84 4127 100 4161
rect -100 4111 100 4127
rect -100 4053 100 4069
rect -100 4019 -84 4053
rect 84 4019 100 4053
rect -100 3981 100 4019
rect -100 3343 100 3381
rect -100 3309 -84 3343
rect 84 3309 100 3343
rect -100 3293 100 3309
rect -100 3235 100 3251
rect -100 3201 -84 3235
rect 84 3201 100 3235
rect -100 3163 100 3201
rect -100 2525 100 2563
rect -100 2491 -84 2525
rect 84 2491 100 2525
rect -100 2475 100 2491
rect -100 2417 100 2433
rect -100 2383 -84 2417
rect 84 2383 100 2417
rect -100 2345 100 2383
rect -100 1707 100 1745
rect -100 1673 -84 1707
rect 84 1673 100 1707
rect -100 1657 100 1673
rect -100 1599 100 1615
rect -100 1565 -84 1599
rect 84 1565 100 1599
rect -100 1527 100 1565
rect -100 889 100 927
rect -100 855 -84 889
rect 84 855 100 889
rect -100 839 100 855
rect -100 781 100 797
rect -100 747 -84 781
rect 84 747 100 781
rect -100 709 100 747
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -747 100 -709
rect -100 -781 -84 -747
rect 84 -781 100 -747
rect -100 -797 100 -781
rect -100 -855 100 -839
rect -100 -889 -84 -855
rect 84 -889 100 -855
rect -100 -927 100 -889
rect -100 -1565 100 -1527
rect -100 -1599 -84 -1565
rect 84 -1599 100 -1565
rect -100 -1615 100 -1599
rect -100 -1673 100 -1657
rect -100 -1707 -84 -1673
rect 84 -1707 100 -1673
rect -100 -1745 100 -1707
rect -100 -2383 100 -2345
rect -100 -2417 -84 -2383
rect 84 -2417 100 -2383
rect -100 -2433 100 -2417
rect -100 -2491 100 -2475
rect -100 -2525 -84 -2491
rect 84 -2525 100 -2491
rect -100 -2563 100 -2525
rect -100 -3201 100 -3163
rect -100 -3235 -84 -3201
rect 84 -3235 100 -3201
rect -100 -3251 100 -3235
rect -100 -3309 100 -3293
rect -100 -3343 -84 -3309
rect 84 -3343 100 -3309
rect -100 -3381 100 -3343
rect -100 -4019 100 -3981
rect -100 -4053 -84 -4019
rect 84 -4053 100 -4019
rect -100 -4069 100 -4053
rect -100 -4127 100 -4111
rect -100 -4161 -84 -4127
rect 84 -4161 100 -4127
rect -100 -4199 100 -4161
rect -100 -4837 100 -4799
rect -100 -4871 -84 -4837
rect 84 -4871 100 -4837
rect -100 -4887 100 -4871
rect -100 -4945 100 -4929
rect -100 -4979 -84 -4945
rect 84 -4979 100 -4945
rect -100 -5017 100 -4979
rect -100 -5655 100 -5617
rect -100 -5689 -84 -5655
rect 84 -5689 100 -5655
rect -100 -5705 100 -5689
rect -100 -5763 100 -5747
rect -100 -5797 -84 -5763
rect 84 -5797 100 -5763
rect -100 -5835 100 -5797
rect -100 -6473 100 -6435
rect -100 -6507 -84 -6473
rect 84 -6507 100 -6473
rect -100 -6523 100 -6507
rect -100 -6581 100 -6565
rect -100 -6615 -84 -6581
rect 84 -6615 100 -6581
rect -100 -6653 100 -6615
rect -100 -7291 100 -7253
rect -100 -7325 -84 -7291
rect 84 -7325 100 -7291
rect -100 -7341 100 -7325
rect -100 -7399 100 -7383
rect -100 -7433 -84 -7399
rect 84 -7433 100 -7399
rect -100 -7471 100 -7433
rect -100 -8109 100 -8071
rect -100 -8143 -84 -8109
rect 84 -8143 100 -8109
rect -100 -8159 100 -8143
rect -100 -8217 100 -8201
rect -100 -8251 -84 -8217
rect 84 -8251 100 -8217
rect -100 -8289 100 -8251
rect -100 -8927 100 -8889
rect -100 -8961 -84 -8927
rect 84 -8961 100 -8927
rect -100 -8977 100 -8961
rect -100 -9035 100 -9019
rect -100 -9069 -84 -9035
rect 84 -9069 100 -9035
rect -100 -9107 100 -9069
rect -100 -9745 100 -9707
rect -100 -9779 -84 -9745
rect 84 -9779 100 -9745
rect -100 -9795 100 -9779
rect -100 -9853 100 -9837
rect -100 -9887 -84 -9853
rect 84 -9887 100 -9853
rect -100 -9925 100 -9887
rect -100 -10563 100 -10525
rect -100 -10597 -84 -10563
rect 84 -10597 100 -10563
rect -100 -10613 100 -10597
rect -100 -10671 100 -10655
rect -100 -10705 -84 -10671
rect 84 -10705 100 -10671
rect -100 -10743 100 -10705
rect -100 -11381 100 -11343
rect -100 -11415 -84 -11381
rect 84 -11415 100 -11381
rect -100 -11431 100 -11415
rect -100 -11489 100 -11473
rect -100 -11523 -84 -11489
rect 84 -11523 100 -11489
rect -100 -11561 100 -11523
rect -100 -12199 100 -12161
rect -100 -12233 -84 -12199
rect 84 -12233 100 -12199
rect -100 -12249 100 -12233
rect -100 -12307 100 -12291
rect -100 -12341 -84 -12307
rect 84 -12341 100 -12307
rect -100 -12379 100 -12341
rect -100 -13017 100 -12979
rect -100 -13051 -84 -13017
rect 84 -13051 100 -13017
rect -100 -13067 100 -13051
rect -100 -13125 100 -13109
rect -100 -13159 -84 -13125
rect 84 -13159 100 -13125
rect -100 -13197 100 -13159
rect -100 -13835 100 -13797
rect -100 -13869 -84 -13835
rect 84 -13869 100 -13835
rect -100 -13885 100 -13869
rect -100 -13943 100 -13927
rect -100 -13977 -84 -13943
rect 84 -13977 100 -13943
rect -100 -14015 100 -13977
rect -100 -14653 100 -14615
rect -100 -14687 -84 -14653
rect 84 -14687 100 -14653
rect -100 -14703 100 -14687
rect -100 -14761 100 -14745
rect -100 -14795 -84 -14761
rect 84 -14795 100 -14761
rect -100 -14833 100 -14795
rect -100 -15471 100 -15433
rect -100 -15505 -84 -15471
rect 84 -15505 100 -15471
rect -100 -15521 100 -15505
rect -100 -15579 100 -15563
rect -100 -15613 -84 -15579
rect 84 -15613 100 -15579
rect -100 -15651 100 -15613
rect -100 -16289 100 -16251
rect -100 -16323 -84 -16289
rect 84 -16323 100 -16289
rect -100 -16339 100 -16323
rect -100 -16397 100 -16381
rect -100 -16431 -84 -16397
rect 84 -16431 100 -16397
rect -100 -16469 100 -16431
rect -100 -17107 100 -17069
rect -100 -17141 -84 -17107
rect 84 -17141 100 -17107
rect -100 -17157 100 -17141
rect -100 -17215 100 -17199
rect -100 -17249 -84 -17215
rect 84 -17249 100 -17215
rect -100 -17287 100 -17249
rect -100 -17925 100 -17887
rect -100 -17959 -84 -17925
rect 84 -17959 100 -17925
rect -100 -17975 100 -17959
rect -100 -18033 100 -18017
rect -100 -18067 -84 -18033
rect 84 -18067 100 -18033
rect -100 -18105 100 -18067
rect -100 -18743 100 -18705
rect -100 -18777 -84 -18743
rect 84 -18777 100 -18743
rect -100 -18793 100 -18777
rect -100 -18851 100 -18835
rect -100 -18885 -84 -18851
rect 84 -18885 100 -18851
rect -100 -18923 100 -18885
rect -100 -19561 100 -19523
rect -100 -19595 -84 -19561
rect 84 -19595 100 -19561
rect -100 -19611 100 -19595
rect -100 -19669 100 -19653
rect -100 -19703 -84 -19669
rect 84 -19703 100 -19669
rect -100 -19741 100 -19703
rect -100 -20379 100 -20341
rect -100 -20413 -84 -20379
rect 84 -20413 100 -20379
rect -100 -20429 100 -20413
rect -100 -20487 100 -20471
rect -100 -20521 -84 -20487
rect 84 -20521 100 -20487
rect -100 -20559 100 -20521
rect -100 -21197 100 -21159
rect -100 -21231 -84 -21197
rect 84 -21231 100 -21197
rect -100 -21247 100 -21231
rect -100 -21305 100 -21289
rect -100 -21339 -84 -21305
rect 84 -21339 100 -21305
rect -100 -21377 100 -21339
rect -100 -22015 100 -21977
rect -100 -22049 -84 -22015
rect 84 -22049 100 -22015
rect -100 -22065 100 -22049
rect -100 -22123 100 -22107
rect -100 -22157 -84 -22123
rect 84 -22157 100 -22123
rect -100 -22195 100 -22157
rect -100 -22833 100 -22795
rect -100 -22867 -84 -22833
rect 84 -22867 100 -22833
rect -100 -22883 100 -22867
rect -100 -22941 100 -22925
rect -100 -22975 -84 -22941
rect 84 -22975 100 -22941
rect -100 -23013 100 -22975
rect -100 -23651 100 -23613
rect -100 -23685 -84 -23651
rect 84 -23685 100 -23651
rect -100 -23701 100 -23685
rect -100 -23759 100 -23743
rect -100 -23793 -84 -23759
rect 84 -23793 100 -23759
rect -100 -23831 100 -23793
rect -100 -24469 100 -24431
rect -100 -24503 -84 -24469
rect 84 -24503 100 -24469
rect -100 -24519 100 -24503
rect -100 -24577 100 -24561
rect -100 -24611 -84 -24577
rect 84 -24611 100 -24577
rect -100 -24649 100 -24611
rect -100 -25287 100 -25249
rect -100 -25321 -84 -25287
rect 84 -25321 100 -25287
rect -100 -25337 100 -25321
rect -100 -25395 100 -25379
rect -100 -25429 -84 -25395
rect 84 -25429 100 -25395
rect -100 -25467 100 -25429
rect -100 -26105 100 -26067
rect -100 -26139 -84 -26105
rect 84 -26139 100 -26105
rect -100 -26155 100 -26139
rect -100 -26213 100 -26197
rect -100 -26247 -84 -26213
rect 84 -26247 100 -26213
rect -100 -26285 100 -26247
rect -100 -26923 100 -26885
rect -100 -26957 -84 -26923
rect 84 -26957 100 -26923
rect -100 -26973 100 -26957
rect -100 -27031 100 -27015
rect -100 -27065 -84 -27031
rect 84 -27065 100 -27031
rect -100 -27103 100 -27065
rect -100 -27741 100 -27703
rect -100 -27775 -84 -27741
rect 84 -27775 100 -27741
rect -100 -27791 100 -27775
rect -100 -27849 100 -27833
rect -100 -27883 -84 -27849
rect 84 -27883 100 -27849
rect -100 -27921 100 -27883
rect -100 -28559 100 -28521
rect -100 -28593 -84 -28559
rect 84 -28593 100 -28559
rect -100 -28609 100 -28593
rect -100 -28667 100 -28651
rect -100 -28701 -84 -28667
rect 84 -28701 100 -28667
rect -100 -28739 100 -28701
rect -100 -29377 100 -29339
rect -100 -29411 -84 -29377
rect 84 -29411 100 -29377
rect -100 -29427 100 -29411
rect -100 -29485 100 -29469
rect -100 -29519 -84 -29485
rect 84 -29519 100 -29485
rect -100 -29557 100 -29519
rect -100 -30195 100 -30157
rect -100 -30229 -84 -30195
rect 84 -30229 100 -30195
rect -100 -30245 100 -30229
rect -100 -30303 100 -30287
rect -100 -30337 -84 -30303
rect 84 -30337 100 -30303
rect -100 -30375 100 -30337
rect -100 -31013 100 -30975
rect -100 -31047 -84 -31013
rect 84 -31047 100 -31013
rect -100 -31063 100 -31047
rect -100 -31121 100 -31105
rect -100 -31155 -84 -31121
rect 84 -31155 100 -31121
rect -100 -31193 100 -31155
rect -100 -31831 100 -31793
rect -100 -31865 -84 -31831
rect 84 -31865 100 -31831
rect -100 -31881 100 -31865
rect -100 -31939 100 -31923
rect -100 -31973 -84 -31939
rect 84 -31973 100 -31939
rect -100 -32011 100 -31973
rect -100 -32649 100 -32611
rect -100 -32683 -84 -32649
rect 84 -32683 100 -32649
rect -100 -32699 100 -32683
rect -100 -32757 100 -32741
rect -100 -32791 -84 -32757
rect 84 -32791 100 -32757
rect -100 -32829 100 -32791
rect -100 -33467 100 -33429
rect -100 -33501 -84 -33467
rect 84 -33501 100 -33467
rect -100 -33517 100 -33501
rect -100 -33575 100 -33559
rect -100 -33609 -84 -33575
rect 84 -33609 100 -33575
rect -100 -33647 100 -33609
rect -100 -34285 100 -34247
rect -100 -34319 -84 -34285
rect 84 -34319 100 -34285
rect -100 -34335 100 -34319
rect -100 -34393 100 -34377
rect -100 -34427 -84 -34393
rect 84 -34427 100 -34393
rect -100 -34465 100 -34427
rect -100 -35103 100 -35065
rect -100 -35137 -84 -35103
rect 84 -35137 100 -35103
rect -100 -35153 100 -35137
rect -100 -35211 100 -35195
rect -100 -35245 -84 -35211
rect 84 -35245 100 -35211
rect -100 -35283 100 -35245
rect -100 -35921 100 -35883
rect -100 -35955 -84 -35921
rect 84 -35955 100 -35921
rect -100 -35971 100 -35955
rect -100 -36029 100 -36013
rect -100 -36063 -84 -36029
rect 84 -36063 100 -36029
rect -100 -36101 100 -36063
rect -100 -36739 100 -36701
rect -100 -36773 -84 -36739
rect 84 -36773 100 -36739
rect -100 -36789 100 -36773
rect -100 -36847 100 -36831
rect -100 -36881 -84 -36847
rect 84 -36881 100 -36847
rect -100 -36919 100 -36881
rect -100 -37557 100 -37519
rect -100 -37591 -84 -37557
rect 84 -37591 100 -37557
rect -100 -37607 100 -37591
rect -100 -37665 100 -37649
rect -100 -37699 -84 -37665
rect 84 -37699 100 -37665
rect -100 -37737 100 -37699
rect -100 -38375 100 -38337
rect -100 -38409 -84 -38375
rect 84 -38409 100 -38375
rect -100 -38425 100 -38409
rect -100 -38483 100 -38467
rect -100 -38517 -84 -38483
rect 84 -38517 100 -38483
rect -100 -38555 100 -38517
rect -100 -39193 100 -39155
rect -100 -39227 -84 -39193
rect 84 -39227 100 -39193
rect -100 -39243 100 -39227
rect -100 -39301 100 -39285
rect -100 -39335 -84 -39301
rect 84 -39335 100 -39301
rect -100 -39373 100 -39335
rect -100 -40011 100 -39973
rect -100 -40045 -84 -40011
rect 84 -40045 100 -40011
rect -100 -40061 100 -40045
rect -100 -40119 100 -40103
rect -100 -40153 -84 -40119
rect 84 -40153 100 -40119
rect -100 -40191 100 -40153
rect -100 -40829 100 -40791
rect -100 -40863 -84 -40829
rect 84 -40863 100 -40829
rect -100 -40879 100 -40863
rect -100 -40937 100 -40921
rect -100 -40971 -84 -40937
rect 84 -40971 100 -40937
rect -100 -41009 100 -40971
rect -100 -41647 100 -41609
rect -100 -41681 -84 -41647
rect 84 -41681 100 -41647
rect -100 -41697 100 -41681
rect -100 -41755 100 -41739
rect -100 -41789 -84 -41755
rect 84 -41789 100 -41755
rect -100 -41827 100 -41789
rect -100 -42465 100 -42427
rect -100 -42499 -84 -42465
rect 84 -42499 100 -42465
rect -100 -42515 100 -42499
rect -100 -42573 100 -42557
rect -100 -42607 -84 -42573
rect 84 -42607 100 -42573
rect -100 -42645 100 -42607
rect -100 -43283 100 -43245
rect -100 -43317 -84 -43283
rect 84 -43317 100 -43283
rect -100 -43333 100 -43317
rect -100 -43391 100 -43375
rect -100 -43425 -84 -43391
rect 84 -43425 100 -43391
rect -100 -43463 100 -43425
rect -100 -44101 100 -44063
rect -100 -44135 -84 -44101
rect 84 -44135 100 -44101
rect -100 -44151 100 -44135
rect -100 -44209 100 -44193
rect -100 -44243 -84 -44209
rect 84 -44243 100 -44209
rect -100 -44281 100 -44243
rect -100 -44919 100 -44881
rect -100 -44953 -84 -44919
rect 84 -44953 100 -44919
rect -100 -44969 100 -44953
rect -100 -45027 100 -45011
rect -100 -45061 -84 -45027
rect 84 -45061 100 -45027
rect -100 -45099 100 -45061
rect -100 -45737 100 -45699
rect -100 -45771 -84 -45737
rect 84 -45771 100 -45737
rect -100 -45787 100 -45771
rect -100 -45845 100 -45829
rect -100 -45879 -84 -45845
rect 84 -45879 100 -45845
rect -100 -45917 100 -45879
rect -100 -46555 100 -46517
rect -100 -46589 -84 -46555
rect 84 -46589 100 -46555
rect -100 -46605 100 -46589
rect -100 -46663 100 -46647
rect -100 -46697 -84 -46663
rect 84 -46697 100 -46663
rect -100 -46735 100 -46697
rect -100 -47373 100 -47335
rect -100 -47407 -84 -47373
rect 84 -47407 100 -47373
rect -100 -47423 100 -47407
rect -100 -47481 100 -47465
rect -100 -47515 -84 -47481
rect 84 -47515 100 -47481
rect -100 -47553 100 -47515
rect -100 -48191 100 -48153
rect -100 -48225 -84 -48191
rect 84 -48225 100 -48191
rect -100 -48241 100 -48225
rect -100 -48299 100 -48283
rect -100 -48333 -84 -48299
rect 84 -48333 100 -48299
rect -100 -48371 100 -48333
rect -100 -49009 100 -48971
rect -100 -49043 -84 -49009
rect 84 -49043 100 -49009
rect -100 -49059 100 -49043
rect -100 -49117 100 -49101
rect -100 -49151 -84 -49117
rect 84 -49151 100 -49117
rect -100 -49189 100 -49151
rect -100 -49827 100 -49789
rect -100 -49861 -84 -49827
rect 84 -49861 100 -49827
rect -100 -49877 100 -49861
rect -100 -49935 100 -49919
rect -100 -49969 -84 -49935
rect 84 -49969 100 -49935
rect -100 -50007 100 -49969
rect -100 -50645 100 -50607
rect -100 -50679 -84 -50645
rect 84 -50679 100 -50645
rect -100 -50695 100 -50679
rect -100 -50753 100 -50737
rect -100 -50787 -84 -50753
rect 84 -50787 100 -50753
rect -100 -50825 100 -50787
rect -100 -51463 100 -51425
rect -100 -51497 -84 -51463
rect 84 -51497 100 -51463
rect -100 -51513 100 -51497
rect -100 -51571 100 -51555
rect -100 -51605 -84 -51571
rect 84 -51605 100 -51571
rect -100 -51643 100 -51605
rect -100 -52281 100 -52243
rect -100 -52315 -84 -52281
rect 84 -52315 100 -52281
rect -100 -52331 100 -52315
rect -100 -52389 100 -52373
rect -100 -52423 -84 -52389
rect 84 -52423 100 -52389
rect -100 -52461 100 -52423
rect -100 -53099 100 -53061
rect -100 -53133 -84 -53099
rect 84 -53133 100 -53099
rect -100 -53149 100 -53133
rect -100 -53207 100 -53191
rect -100 -53241 -84 -53207
rect 84 -53241 100 -53207
rect -100 -53279 100 -53241
rect -100 -53917 100 -53879
rect -100 -53951 -84 -53917
rect 84 -53951 100 -53917
rect -100 -53967 100 -53951
rect -100 -54025 100 -54009
rect -100 -54059 -84 -54025
rect 84 -54059 100 -54025
rect -100 -54097 100 -54059
rect -100 -54735 100 -54697
rect -100 -54769 -84 -54735
rect 84 -54769 100 -54735
rect -100 -54785 100 -54769
rect -100 -54843 100 -54827
rect -100 -54877 -84 -54843
rect 84 -54877 100 -54843
rect -100 -54915 100 -54877
rect -100 -55553 100 -55515
rect -100 -55587 -84 -55553
rect 84 -55587 100 -55553
rect -100 -55603 100 -55587
rect -100 -55661 100 -55645
rect -100 -55695 -84 -55661
rect 84 -55695 100 -55661
rect -100 -55733 100 -55695
rect -100 -56371 100 -56333
rect -100 -56405 -84 -56371
rect 84 -56405 100 -56371
rect -100 -56421 100 -56405
rect -100 -56479 100 -56463
rect -100 -56513 -84 -56479
rect 84 -56513 100 -56479
rect -100 -56551 100 -56513
rect -100 -57189 100 -57151
rect -100 -57223 -84 -57189
rect 84 -57223 100 -57189
rect -100 -57239 100 -57223
rect -100 -57297 100 -57281
rect -100 -57331 -84 -57297
rect 84 -57331 100 -57297
rect -100 -57369 100 -57331
rect -100 -58007 100 -57969
rect -100 -58041 -84 -58007
rect 84 -58041 100 -58007
rect -100 -58057 100 -58041
rect -100 -58115 100 -58099
rect -100 -58149 -84 -58115
rect 84 -58149 100 -58115
rect -100 -58187 100 -58149
rect -100 -58825 100 -58787
rect -100 -58859 -84 -58825
rect 84 -58859 100 -58825
rect -100 -58875 100 -58859
rect -100 -58933 100 -58917
rect -100 -58967 -84 -58933
rect 84 -58967 100 -58933
rect -100 -59005 100 -58967
rect -100 -59643 100 -59605
rect -100 -59677 -84 -59643
rect 84 -59677 100 -59643
rect -100 -59693 100 -59677
rect -100 -59751 100 -59735
rect -100 -59785 -84 -59751
rect 84 -59785 100 -59751
rect -100 -59823 100 -59785
rect -100 -60461 100 -60423
rect -100 -60495 -84 -60461
rect 84 -60495 100 -60461
rect -100 -60511 100 -60495
rect -100 -60569 100 -60553
rect -100 -60603 -84 -60569
rect 84 -60603 100 -60569
rect -100 -60641 100 -60603
rect -100 -61279 100 -61241
rect -100 -61313 -84 -61279
rect 84 -61313 100 -61279
rect -100 -61329 100 -61313
rect -100 -61387 100 -61371
rect -100 -61421 -84 -61387
rect 84 -61421 100 -61387
rect -100 -61459 100 -61421
rect -100 -62097 100 -62059
rect -100 -62131 -84 -62097
rect 84 -62131 100 -62097
rect -100 -62147 100 -62131
rect -100 -62205 100 -62189
rect -100 -62239 -84 -62205
rect 84 -62239 100 -62205
rect -100 -62277 100 -62239
rect -100 -62915 100 -62877
rect -100 -62949 -84 -62915
rect 84 -62949 100 -62915
rect -100 -62965 100 -62949
rect -100 -63023 100 -63007
rect -100 -63057 -84 -63023
rect 84 -63057 100 -63023
rect -100 -63095 100 -63057
rect -100 -63733 100 -63695
rect -100 -63767 -84 -63733
rect 84 -63767 100 -63733
rect -100 -63783 100 -63767
rect -100 -63841 100 -63825
rect -100 -63875 -84 -63841
rect 84 -63875 100 -63841
rect -100 -63913 100 -63875
rect -100 -64551 100 -64513
rect -100 -64585 -84 -64551
rect 84 -64585 100 -64551
rect -100 -64601 100 -64585
rect -100 -64659 100 -64643
rect -100 -64693 -84 -64659
rect 84 -64693 100 -64659
rect -100 -64731 100 -64693
rect -100 -65369 100 -65331
rect -100 -65403 -84 -65369
rect 84 -65403 100 -65369
rect -100 -65419 100 -65403
rect -100 -65477 100 -65461
rect -100 -65511 -84 -65477
rect 84 -65511 100 -65477
rect -100 -65549 100 -65511
rect -100 -66187 100 -66149
rect -100 -66221 -84 -66187
rect 84 -66221 100 -66187
rect -100 -66237 100 -66221
rect -100 -66295 100 -66279
rect -100 -66329 -84 -66295
rect 84 -66329 100 -66295
rect -100 -66367 100 -66329
rect -100 -67005 100 -66967
rect -100 -67039 -84 -67005
rect 84 -67039 100 -67005
rect -100 -67055 100 -67039
rect -100 -67113 100 -67097
rect -100 -67147 -84 -67113
rect 84 -67147 100 -67113
rect -100 -67185 100 -67147
rect -100 -67823 100 -67785
rect -100 -67857 -84 -67823
rect 84 -67857 100 -67823
rect -100 -67873 100 -67857
rect -100 -67931 100 -67915
rect -100 -67965 -84 -67931
rect 84 -67965 100 -67931
rect -100 -68003 100 -67965
rect -100 -68641 100 -68603
rect -100 -68675 -84 -68641
rect 84 -68675 100 -68641
rect -100 -68691 100 -68675
rect -100 -68749 100 -68733
rect -100 -68783 -84 -68749
rect 84 -68783 100 -68749
rect -100 -68821 100 -68783
rect -100 -69459 100 -69421
rect -100 -69493 -84 -69459
rect 84 -69493 100 -69459
rect -100 -69509 100 -69493
rect -100 -69567 100 -69551
rect -100 -69601 -84 -69567
rect 84 -69601 100 -69567
rect -100 -69639 100 -69601
rect -100 -70277 100 -70239
rect -100 -70311 -84 -70277
rect 84 -70311 100 -70277
rect -100 -70327 100 -70311
rect -100 -70385 100 -70369
rect -100 -70419 -84 -70385
rect 84 -70419 100 -70385
rect -100 -70457 100 -70419
rect -100 -71095 100 -71057
rect -100 -71129 -84 -71095
rect 84 -71129 100 -71095
rect -100 -71145 100 -71129
rect -100 -71203 100 -71187
rect -100 -71237 -84 -71203
rect 84 -71237 100 -71203
rect -100 -71275 100 -71237
rect -100 -71913 100 -71875
rect -100 -71947 -84 -71913
rect 84 -71947 100 -71913
rect -100 -71963 100 -71947
rect -100 -72021 100 -72005
rect -100 -72055 -84 -72021
rect 84 -72055 100 -72021
rect -100 -72093 100 -72055
rect -100 -72731 100 -72693
rect -100 -72765 -84 -72731
rect 84 -72765 100 -72731
rect -100 -72781 100 -72765
rect -100 -72839 100 -72823
rect -100 -72873 -84 -72839
rect 84 -72873 100 -72839
rect -100 -72911 100 -72873
rect -100 -73549 100 -73511
rect -100 -73583 -84 -73549
rect 84 -73583 100 -73549
rect -100 -73599 100 -73583
rect -100 -73657 100 -73641
rect -100 -73691 -84 -73657
rect 84 -73691 100 -73657
rect -100 -73729 100 -73691
rect -100 -74367 100 -74329
rect -100 -74401 -84 -74367
rect 84 -74401 100 -74367
rect -100 -74417 100 -74401
rect -100 -74475 100 -74459
rect -100 -74509 -84 -74475
rect 84 -74509 100 -74475
rect -100 -74547 100 -74509
rect -100 -75185 100 -75147
rect -100 -75219 -84 -75185
rect 84 -75219 100 -75185
rect -100 -75235 100 -75219
rect -100 -75293 100 -75277
rect -100 -75327 -84 -75293
rect 84 -75327 100 -75293
rect -100 -75365 100 -75327
rect -100 -76003 100 -75965
rect -100 -76037 -84 -76003
rect 84 -76037 100 -76003
rect -100 -76053 100 -76037
rect -100 -76111 100 -76095
rect -100 -76145 -84 -76111
rect 84 -76145 100 -76111
rect -100 -76183 100 -76145
rect -100 -76821 100 -76783
rect -100 -76855 -84 -76821
rect 84 -76855 100 -76821
rect -100 -76871 100 -76855
rect -100 -76929 100 -76913
rect -100 -76963 -84 -76929
rect 84 -76963 100 -76929
rect -100 -77001 100 -76963
rect -100 -77639 100 -77601
rect -100 -77673 -84 -77639
rect 84 -77673 100 -77639
rect -100 -77689 100 -77673
rect -100 -77747 100 -77731
rect -100 -77781 -84 -77747
rect 84 -77781 100 -77747
rect -100 -77819 100 -77781
rect -100 -78457 100 -78419
rect -100 -78491 -84 -78457
rect 84 -78491 100 -78457
rect -100 -78507 100 -78491
rect -100 -78565 100 -78549
rect -100 -78599 -84 -78565
rect 84 -78599 100 -78565
rect -100 -78637 100 -78599
rect -100 -79275 100 -79237
rect -100 -79309 -84 -79275
rect 84 -79309 100 -79275
rect -100 -79325 100 -79309
rect -100 -79383 100 -79367
rect -100 -79417 -84 -79383
rect 84 -79417 100 -79383
rect -100 -79455 100 -79417
rect -100 -80093 100 -80055
rect -100 -80127 -84 -80093
rect 84 -80127 100 -80093
rect -100 -80143 100 -80127
rect -100 -80201 100 -80185
rect -100 -80235 -84 -80201
rect 84 -80235 100 -80201
rect -100 -80273 100 -80235
rect -100 -80911 100 -80873
rect -100 -80945 -84 -80911
rect 84 -80945 100 -80911
rect -100 -80961 100 -80945
rect -100 -81019 100 -81003
rect -100 -81053 -84 -81019
rect 84 -81053 100 -81019
rect -100 -81091 100 -81053
rect -100 -81729 100 -81691
rect -100 -81763 -84 -81729
rect 84 -81763 100 -81729
rect -100 -81779 100 -81763
rect -100 -81837 100 -81821
rect -100 -81871 -84 -81837
rect 84 -81871 100 -81837
rect -100 -81909 100 -81871
rect -100 -82547 100 -82509
rect -100 -82581 -84 -82547
rect 84 -82581 100 -82547
rect -100 -82597 100 -82581
rect -100 -82655 100 -82639
rect -100 -82689 -84 -82655
rect 84 -82689 100 -82655
rect -100 -82727 100 -82689
rect -100 -83365 100 -83327
rect -100 -83399 -84 -83365
rect 84 -83399 100 -83365
rect -100 -83415 100 -83399
rect -100 -83473 100 -83457
rect -100 -83507 -84 -83473
rect 84 -83507 100 -83473
rect -100 -83545 100 -83507
rect -100 -84183 100 -84145
rect -100 -84217 -84 -84183
rect 84 -84217 100 -84183
rect -100 -84233 100 -84217
rect -100 -84291 100 -84275
rect -100 -84325 -84 -84291
rect 84 -84325 100 -84291
rect -100 -84363 100 -84325
rect -100 -85001 100 -84963
rect -100 -85035 -84 -85001
rect 84 -85035 100 -85001
rect -100 -85051 100 -85035
rect -100 -85109 100 -85093
rect -100 -85143 -84 -85109
rect 84 -85143 100 -85109
rect -100 -85181 100 -85143
rect -100 -85819 100 -85781
rect -100 -85853 -84 -85819
rect 84 -85853 100 -85819
rect -100 -85869 100 -85853
rect -100 -85927 100 -85911
rect -100 -85961 -84 -85927
rect 84 -85961 100 -85927
rect -100 -85999 100 -85961
rect -100 -86637 100 -86599
rect -100 -86671 -84 -86637
rect 84 -86671 100 -86637
rect -100 -86687 100 -86671
rect -100 -86745 100 -86729
rect -100 -86779 -84 -86745
rect 84 -86779 100 -86745
rect -100 -86817 100 -86779
rect -100 -87455 100 -87417
rect -100 -87489 -84 -87455
rect 84 -87489 100 -87455
rect -100 -87505 100 -87489
rect -100 -87563 100 -87547
rect -100 -87597 -84 -87563
rect 84 -87597 100 -87563
rect -100 -87635 100 -87597
rect -100 -88273 100 -88235
rect -100 -88307 -84 -88273
rect 84 -88307 100 -88273
rect -100 -88323 100 -88307
rect -100 -88381 100 -88365
rect -100 -88415 -84 -88381
rect 84 -88415 100 -88381
rect -100 -88453 100 -88415
rect -100 -89091 100 -89053
rect -100 -89125 -84 -89091
rect 84 -89125 100 -89091
rect -100 -89141 100 -89125
rect -100 -89199 100 -89183
rect -100 -89233 -84 -89199
rect 84 -89233 100 -89199
rect -100 -89271 100 -89233
rect -100 -89909 100 -89871
rect -100 -89943 -84 -89909
rect 84 -89943 100 -89909
rect -100 -89959 100 -89943
rect -100 -90017 100 -90001
rect -100 -90051 -84 -90017
rect 84 -90051 100 -90017
rect -100 -90089 100 -90051
rect -100 -90727 100 -90689
rect -100 -90761 -84 -90727
rect 84 -90761 100 -90727
rect -100 -90777 100 -90761
rect -100 -90835 100 -90819
rect -100 -90869 -84 -90835
rect 84 -90869 100 -90835
rect -100 -90907 100 -90869
rect -100 -91545 100 -91507
rect -100 -91579 -84 -91545
rect 84 -91579 100 -91545
rect -100 -91595 100 -91579
rect -100 -91653 100 -91637
rect -100 -91687 -84 -91653
rect 84 -91687 100 -91653
rect -100 -91725 100 -91687
rect -100 -92363 100 -92325
rect -100 -92397 -84 -92363
rect 84 -92397 100 -92363
rect -100 -92413 100 -92397
rect -100 -92471 100 -92455
rect -100 -92505 -84 -92471
rect 84 -92505 100 -92471
rect -100 -92543 100 -92505
rect -100 -93181 100 -93143
rect -100 -93215 -84 -93181
rect 84 -93215 100 -93181
rect -100 -93231 100 -93215
rect -100 -93289 100 -93273
rect -100 -93323 -84 -93289
rect 84 -93323 100 -93289
rect -100 -93361 100 -93323
rect -100 -93999 100 -93961
rect -100 -94033 -84 -93999
rect 84 -94033 100 -93999
rect -100 -94049 100 -94033
rect -100 -94107 100 -94091
rect -100 -94141 -84 -94107
rect 84 -94141 100 -94107
rect -100 -94179 100 -94141
rect -100 -94817 100 -94779
rect -100 -94851 -84 -94817
rect 84 -94851 100 -94817
rect -100 -94867 100 -94851
rect -100 -94925 100 -94909
rect -100 -94959 -84 -94925
rect 84 -94959 100 -94925
rect -100 -94997 100 -94959
rect -100 -95635 100 -95597
rect -100 -95669 -84 -95635
rect 84 -95669 100 -95635
rect -100 -95685 100 -95669
rect -100 -95743 100 -95727
rect -100 -95777 -84 -95743
rect 84 -95777 100 -95743
rect -100 -95815 100 -95777
rect -100 -96453 100 -96415
rect -100 -96487 -84 -96453
rect 84 -96487 100 -96453
rect -100 -96503 100 -96487
rect -100 -96561 100 -96545
rect -100 -96595 -84 -96561
rect 84 -96595 100 -96561
rect -100 -96633 100 -96595
rect -100 -97271 100 -97233
rect -100 -97305 -84 -97271
rect 84 -97305 100 -97271
rect -100 -97321 100 -97305
rect -100 -97379 100 -97363
rect -100 -97413 -84 -97379
rect 84 -97413 100 -97379
rect -100 -97451 100 -97413
rect -100 -98089 100 -98051
rect -100 -98123 -84 -98089
rect 84 -98123 100 -98089
rect -100 -98139 100 -98123
rect -100 -98197 100 -98181
rect -100 -98231 -84 -98197
rect 84 -98231 100 -98197
rect -100 -98269 100 -98231
rect -100 -98907 100 -98869
rect -100 -98941 -84 -98907
rect 84 -98941 100 -98907
rect -100 -98957 100 -98941
rect -100 -99015 100 -98999
rect -100 -99049 -84 -99015
rect 84 -99049 100 -99015
rect -100 -99087 100 -99049
rect -100 -99725 100 -99687
rect -100 -99759 -84 -99725
rect 84 -99759 100 -99725
rect -100 -99775 100 -99759
rect -100 -99833 100 -99817
rect -100 -99867 -84 -99833
rect 84 -99867 100 -99833
rect -100 -99905 100 -99867
rect -100 -100543 100 -100505
rect -100 -100577 -84 -100543
rect 84 -100577 100 -100543
rect -100 -100593 100 -100577
rect -100 -100651 100 -100635
rect -100 -100685 -84 -100651
rect 84 -100685 100 -100651
rect -100 -100723 100 -100685
rect -100 -101361 100 -101323
rect -100 -101395 -84 -101361
rect 84 -101395 100 -101361
rect -100 -101411 100 -101395
rect -100 -101469 100 -101453
rect -100 -101503 -84 -101469
rect 84 -101503 100 -101469
rect -100 -101541 100 -101503
rect -100 -102179 100 -102141
rect -100 -102213 -84 -102179
rect 84 -102213 100 -102179
rect -100 -102229 100 -102213
rect -100 -102287 100 -102271
rect -100 -102321 -84 -102287
rect 84 -102321 100 -102287
rect -100 -102359 100 -102321
rect -100 -102997 100 -102959
rect -100 -103031 -84 -102997
rect 84 -103031 100 -102997
rect -100 -103047 100 -103031
rect -100 -103105 100 -103089
rect -100 -103139 -84 -103105
rect 84 -103139 100 -103105
rect -100 -103177 100 -103139
rect -100 -103815 100 -103777
rect -100 -103849 -84 -103815
rect 84 -103849 100 -103815
rect -100 -103865 100 -103849
rect -100 -103923 100 -103907
rect -100 -103957 -84 -103923
rect 84 -103957 100 -103923
rect -100 -103995 100 -103957
rect -100 -104633 100 -104595
rect -100 -104667 -84 -104633
rect 84 -104667 100 -104633
rect -100 -104683 100 -104667
<< polycont >>
rect -84 104633 84 104667
rect -84 103923 84 103957
rect -84 103815 84 103849
rect -84 103105 84 103139
rect -84 102997 84 103031
rect -84 102287 84 102321
rect -84 102179 84 102213
rect -84 101469 84 101503
rect -84 101361 84 101395
rect -84 100651 84 100685
rect -84 100543 84 100577
rect -84 99833 84 99867
rect -84 99725 84 99759
rect -84 99015 84 99049
rect -84 98907 84 98941
rect -84 98197 84 98231
rect -84 98089 84 98123
rect -84 97379 84 97413
rect -84 97271 84 97305
rect -84 96561 84 96595
rect -84 96453 84 96487
rect -84 95743 84 95777
rect -84 95635 84 95669
rect -84 94925 84 94959
rect -84 94817 84 94851
rect -84 94107 84 94141
rect -84 93999 84 94033
rect -84 93289 84 93323
rect -84 93181 84 93215
rect -84 92471 84 92505
rect -84 92363 84 92397
rect -84 91653 84 91687
rect -84 91545 84 91579
rect -84 90835 84 90869
rect -84 90727 84 90761
rect -84 90017 84 90051
rect -84 89909 84 89943
rect -84 89199 84 89233
rect -84 89091 84 89125
rect -84 88381 84 88415
rect -84 88273 84 88307
rect -84 87563 84 87597
rect -84 87455 84 87489
rect -84 86745 84 86779
rect -84 86637 84 86671
rect -84 85927 84 85961
rect -84 85819 84 85853
rect -84 85109 84 85143
rect -84 85001 84 85035
rect -84 84291 84 84325
rect -84 84183 84 84217
rect -84 83473 84 83507
rect -84 83365 84 83399
rect -84 82655 84 82689
rect -84 82547 84 82581
rect -84 81837 84 81871
rect -84 81729 84 81763
rect -84 81019 84 81053
rect -84 80911 84 80945
rect -84 80201 84 80235
rect -84 80093 84 80127
rect -84 79383 84 79417
rect -84 79275 84 79309
rect -84 78565 84 78599
rect -84 78457 84 78491
rect -84 77747 84 77781
rect -84 77639 84 77673
rect -84 76929 84 76963
rect -84 76821 84 76855
rect -84 76111 84 76145
rect -84 76003 84 76037
rect -84 75293 84 75327
rect -84 75185 84 75219
rect -84 74475 84 74509
rect -84 74367 84 74401
rect -84 73657 84 73691
rect -84 73549 84 73583
rect -84 72839 84 72873
rect -84 72731 84 72765
rect -84 72021 84 72055
rect -84 71913 84 71947
rect -84 71203 84 71237
rect -84 71095 84 71129
rect -84 70385 84 70419
rect -84 70277 84 70311
rect -84 69567 84 69601
rect -84 69459 84 69493
rect -84 68749 84 68783
rect -84 68641 84 68675
rect -84 67931 84 67965
rect -84 67823 84 67857
rect -84 67113 84 67147
rect -84 67005 84 67039
rect -84 66295 84 66329
rect -84 66187 84 66221
rect -84 65477 84 65511
rect -84 65369 84 65403
rect -84 64659 84 64693
rect -84 64551 84 64585
rect -84 63841 84 63875
rect -84 63733 84 63767
rect -84 63023 84 63057
rect -84 62915 84 62949
rect -84 62205 84 62239
rect -84 62097 84 62131
rect -84 61387 84 61421
rect -84 61279 84 61313
rect -84 60569 84 60603
rect -84 60461 84 60495
rect -84 59751 84 59785
rect -84 59643 84 59677
rect -84 58933 84 58967
rect -84 58825 84 58859
rect -84 58115 84 58149
rect -84 58007 84 58041
rect -84 57297 84 57331
rect -84 57189 84 57223
rect -84 56479 84 56513
rect -84 56371 84 56405
rect -84 55661 84 55695
rect -84 55553 84 55587
rect -84 54843 84 54877
rect -84 54735 84 54769
rect -84 54025 84 54059
rect -84 53917 84 53951
rect -84 53207 84 53241
rect -84 53099 84 53133
rect -84 52389 84 52423
rect -84 52281 84 52315
rect -84 51571 84 51605
rect -84 51463 84 51497
rect -84 50753 84 50787
rect -84 50645 84 50679
rect -84 49935 84 49969
rect -84 49827 84 49861
rect -84 49117 84 49151
rect -84 49009 84 49043
rect -84 48299 84 48333
rect -84 48191 84 48225
rect -84 47481 84 47515
rect -84 47373 84 47407
rect -84 46663 84 46697
rect -84 46555 84 46589
rect -84 45845 84 45879
rect -84 45737 84 45771
rect -84 45027 84 45061
rect -84 44919 84 44953
rect -84 44209 84 44243
rect -84 44101 84 44135
rect -84 43391 84 43425
rect -84 43283 84 43317
rect -84 42573 84 42607
rect -84 42465 84 42499
rect -84 41755 84 41789
rect -84 41647 84 41681
rect -84 40937 84 40971
rect -84 40829 84 40863
rect -84 40119 84 40153
rect -84 40011 84 40045
rect -84 39301 84 39335
rect -84 39193 84 39227
rect -84 38483 84 38517
rect -84 38375 84 38409
rect -84 37665 84 37699
rect -84 37557 84 37591
rect -84 36847 84 36881
rect -84 36739 84 36773
rect -84 36029 84 36063
rect -84 35921 84 35955
rect -84 35211 84 35245
rect -84 35103 84 35137
rect -84 34393 84 34427
rect -84 34285 84 34319
rect -84 33575 84 33609
rect -84 33467 84 33501
rect -84 32757 84 32791
rect -84 32649 84 32683
rect -84 31939 84 31973
rect -84 31831 84 31865
rect -84 31121 84 31155
rect -84 31013 84 31047
rect -84 30303 84 30337
rect -84 30195 84 30229
rect -84 29485 84 29519
rect -84 29377 84 29411
rect -84 28667 84 28701
rect -84 28559 84 28593
rect -84 27849 84 27883
rect -84 27741 84 27775
rect -84 27031 84 27065
rect -84 26923 84 26957
rect -84 26213 84 26247
rect -84 26105 84 26139
rect -84 25395 84 25429
rect -84 25287 84 25321
rect -84 24577 84 24611
rect -84 24469 84 24503
rect -84 23759 84 23793
rect -84 23651 84 23685
rect -84 22941 84 22975
rect -84 22833 84 22867
rect -84 22123 84 22157
rect -84 22015 84 22049
rect -84 21305 84 21339
rect -84 21197 84 21231
rect -84 20487 84 20521
rect -84 20379 84 20413
rect -84 19669 84 19703
rect -84 19561 84 19595
rect -84 18851 84 18885
rect -84 18743 84 18777
rect -84 18033 84 18067
rect -84 17925 84 17959
rect -84 17215 84 17249
rect -84 17107 84 17141
rect -84 16397 84 16431
rect -84 16289 84 16323
rect -84 15579 84 15613
rect -84 15471 84 15505
rect -84 14761 84 14795
rect -84 14653 84 14687
rect -84 13943 84 13977
rect -84 13835 84 13869
rect -84 13125 84 13159
rect -84 13017 84 13051
rect -84 12307 84 12341
rect -84 12199 84 12233
rect -84 11489 84 11523
rect -84 11381 84 11415
rect -84 10671 84 10705
rect -84 10563 84 10597
rect -84 9853 84 9887
rect -84 9745 84 9779
rect -84 9035 84 9069
rect -84 8927 84 8961
rect -84 8217 84 8251
rect -84 8109 84 8143
rect -84 7399 84 7433
rect -84 7291 84 7325
rect -84 6581 84 6615
rect -84 6473 84 6507
rect -84 5763 84 5797
rect -84 5655 84 5689
rect -84 4945 84 4979
rect -84 4837 84 4871
rect -84 4127 84 4161
rect -84 4019 84 4053
rect -84 3309 84 3343
rect -84 3201 84 3235
rect -84 2491 84 2525
rect -84 2383 84 2417
rect -84 1673 84 1707
rect -84 1565 84 1599
rect -84 855 84 889
rect -84 747 84 781
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -781 84 -747
rect -84 -889 84 -855
rect -84 -1599 84 -1565
rect -84 -1707 84 -1673
rect -84 -2417 84 -2383
rect -84 -2525 84 -2491
rect -84 -3235 84 -3201
rect -84 -3343 84 -3309
rect -84 -4053 84 -4019
rect -84 -4161 84 -4127
rect -84 -4871 84 -4837
rect -84 -4979 84 -4945
rect -84 -5689 84 -5655
rect -84 -5797 84 -5763
rect -84 -6507 84 -6473
rect -84 -6615 84 -6581
rect -84 -7325 84 -7291
rect -84 -7433 84 -7399
rect -84 -8143 84 -8109
rect -84 -8251 84 -8217
rect -84 -8961 84 -8927
rect -84 -9069 84 -9035
rect -84 -9779 84 -9745
rect -84 -9887 84 -9853
rect -84 -10597 84 -10563
rect -84 -10705 84 -10671
rect -84 -11415 84 -11381
rect -84 -11523 84 -11489
rect -84 -12233 84 -12199
rect -84 -12341 84 -12307
rect -84 -13051 84 -13017
rect -84 -13159 84 -13125
rect -84 -13869 84 -13835
rect -84 -13977 84 -13943
rect -84 -14687 84 -14653
rect -84 -14795 84 -14761
rect -84 -15505 84 -15471
rect -84 -15613 84 -15579
rect -84 -16323 84 -16289
rect -84 -16431 84 -16397
rect -84 -17141 84 -17107
rect -84 -17249 84 -17215
rect -84 -17959 84 -17925
rect -84 -18067 84 -18033
rect -84 -18777 84 -18743
rect -84 -18885 84 -18851
rect -84 -19595 84 -19561
rect -84 -19703 84 -19669
rect -84 -20413 84 -20379
rect -84 -20521 84 -20487
rect -84 -21231 84 -21197
rect -84 -21339 84 -21305
rect -84 -22049 84 -22015
rect -84 -22157 84 -22123
rect -84 -22867 84 -22833
rect -84 -22975 84 -22941
rect -84 -23685 84 -23651
rect -84 -23793 84 -23759
rect -84 -24503 84 -24469
rect -84 -24611 84 -24577
rect -84 -25321 84 -25287
rect -84 -25429 84 -25395
rect -84 -26139 84 -26105
rect -84 -26247 84 -26213
rect -84 -26957 84 -26923
rect -84 -27065 84 -27031
rect -84 -27775 84 -27741
rect -84 -27883 84 -27849
rect -84 -28593 84 -28559
rect -84 -28701 84 -28667
rect -84 -29411 84 -29377
rect -84 -29519 84 -29485
rect -84 -30229 84 -30195
rect -84 -30337 84 -30303
rect -84 -31047 84 -31013
rect -84 -31155 84 -31121
rect -84 -31865 84 -31831
rect -84 -31973 84 -31939
rect -84 -32683 84 -32649
rect -84 -32791 84 -32757
rect -84 -33501 84 -33467
rect -84 -33609 84 -33575
rect -84 -34319 84 -34285
rect -84 -34427 84 -34393
rect -84 -35137 84 -35103
rect -84 -35245 84 -35211
rect -84 -35955 84 -35921
rect -84 -36063 84 -36029
rect -84 -36773 84 -36739
rect -84 -36881 84 -36847
rect -84 -37591 84 -37557
rect -84 -37699 84 -37665
rect -84 -38409 84 -38375
rect -84 -38517 84 -38483
rect -84 -39227 84 -39193
rect -84 -39335 84 -39301
rect -84 -40045 84 -40011
rect -84 -40153 84 -40119
rect -84 -40863 84 -40829
rect -84 -40971 84 -40937
rect -84 -41681 84 -41647
rect -84 -41789 84 -41755
rect -84 -42499 84 -42465
rect -84 -42607 84 -42573
rect -84 -43317 84 -43283
rect -84 -43425 84 -43391
rect -84 -44135 84 -44101
rect -84 -44243 84 -44209
rect -84 -44953 84 -44919
rect -84 -45061 84 -45027
rect -84 -45771 84 -45737
rect -84 -45879 84 -45845
rect -84 -46589 84 -46555
rect -84 -46697 84 -46663
rect -84 -47407 84 -47373
rect -84 -47515 84 -47481
rect -84 -48225 84 -48191
rect -84 -48333 84 -48299
rect -84 -49043 84 -49009
rect -84 -49151 84 -49117
rect -84 -49861 84 -49827
rect -84 -49969 84 -49935
rect -84 -50679 84 -50645
rect -84 -50787 84 -50753
rect -84 -51497 84 -51463
rect -84 -51605 84 -51571
rect -84 -52315 84 -52281
rect -84 -52423 84 -52389
rect -84 -53133 84 -53099
rect -84 -53241 84 -53207
rect -84 -53951 84 -53917
rect -84 -54059 84 -54025
rect -84 -54769 84 -54735
rect -84 -54877 84 -54843
rect -84 -55587 84 -55553
rect -84 -55695 84 -55661
rect -84 -56405 84 -56371
rect -84 -56513 84 -56479
rect -84 -57223 84 -57189
rect -84 -57331 84 -57297
rect -84 -58041 84 -58007
rect -84 -58149 84 -58115
rect -84 -58859 84 -58825
rect -84 -58967 84 -58933
rect -84 -59677 84 -59643
rect -84 -59785 84 -59751
rect -84 -60495 84 -60461
rect -84 -60603 84 -60569
rect -84 -61313 84 -61279
rect -84 -61421 84 -61387
rect -84 -62131 84 -62097
rect -84 -62239 84 -62205
rect -84 -62949 84 -62915
rect -84 -63057 84 -63023
rect -84 -63767 84 -63733
rect -84 -63875 84 -63841
rect -84 -64585 84 -64551
rect -84 -64693 84 -64659
rect -84 -65403 84 -65369
rect -84 -65511 84 -65477
rect -84 -66221 84 -66187
rect -84 -66329 84 -66295
rect -84 -67039 84 -67005
rect -84 -67147 84 -67113
rect -84 -67857 84 -67823
rect -84 -67965 84 -67931
rect -84 -68675 84 -68641
rect -84 -68783 84 -68749
rect -84 -69493 84 -69459
rect -84 -69601 84 -69567
rect -84 -70311 84 -70277
rect -84 -70419 84 -70385
rect -84 -71129 84 -71095
rect -84 -71237 84 -71203
rect -84 -71947 84 -71913
rect -84 -72055 84 -72021
rect -84 -72765 84 -72731
rect -84 -72873 84 -72839
rect -84 -73583 84 -73549
rect -84 -73691 84 -73657
rect -84 -74401 84 -74367
rect -84 -74509 84 -74475
rect -84 -75219 84 -75185
rect -84 -75327 84 -75293
rect -84 -76037 84 -76003
rect -84 -76145 84 -76111
rect -84 -76855 84 -76821
rect -84 -76963 84 -76929
rect -84 -77673 84 -77639
rect -84 -77781 84 -77747
rect -84 -78491 84 -78457
rect -84 -78599 84 -78565
rect -84 -79309 84 -79275
rect -84 -79417 84 -79383
rect -84 -80127 84 -80093
rect -84 -80235 84 -80201
rect -84 -80945 84 -80911
rect -84 -81053 84 -81019
rect -84 -81763 84 -81729
rect -84 -81871 84 -81837
rect -84 -82581 84 -82547
rect -84 -82689 84 -82655
rect -84 -83399 84 -83365
rect -84 -83507 84 -83473
rect -84 -84217 84 -84183
rect -84 -84325 84 -84291
rect -84 -85035 84 -85001
rect -84 -85143 84 -85109
rect -84 -85853 84 -85819
rect -84 -85961 84 -85927
rect -84 -86671 84 -86637
rect -84 -86779 84 -86745
rect -84 -87489 84 -87455
rect -84 -87597 84 -87563
rect -84 -88307 84 -88273
rect -84 -88415 84 -88381
rect -84 -89125 84 -89091
rect -84 -89233 84 -89199
rect -84 -89943 84 -89909
rect -84 -90051 84 -90017
rect -84 -90761 84 -90727
rect -84 -90869 84 -90835
rect -84 -91579 84 -91545
rect -84 -91687 84 -91653
rect -84 -92397 84 -92363
rect -84 -92505 84 -92471
rect -84 -93215 84 -93181
rect -84 -93323 84 -93289
rect -84 -94033 84 -93999
rect -84 -94141 84 -94107
rect -84 -94851 84 -94817
rect -84 -94959 84 -94925
rect -84 -95669 84 -95635
rect -84 -95777 84 -95743
rect -84 -96487 84 -96453
rect -84 -96595 84 -96561
rect -84 -97305 84 -97271
rect -84 -97413 84 -97379
rect -84 -98123 84 -98089
rect -84 -98231 84 -98197
rect -84 -98941 84 -98907
rect -84 -99049 84 -99015
rect -84 -99759 84 -99725
rect -84 -99867 84 -99833
rect -84 -100577 84 -100543
rect -84 -100685 84 -100651
rect -84 -101395 84 -101361
rect -84 -101503 84 -101469
rect -84 -102213 84 -102179
rect -84 -102321 84 -102287
rect -84 -103031 84 -102997
rect -84 -103139 84 -103105
rect -84 -103849 84 -103815
rect -84 -103957 84 -103923
rect -84 -104667 84 -104633
<< locali >>
rect -280 104771 -184 104805
rect 184 104771 280 104805
rect -280 104709 -246 104771
rect 246 104709 280 104771
rect -100 104633 -84 104667
rect 84 104633 100 104667
rect -146 104583 -112 104599
rect -146 103991 -112 104007
rect 112 104583 146 104599
rect 112 103991 146 104007
rect -100 103923 -84 103957
rect 84 103923 100 103957
rect -100 103815 -84 103849
rect 84 103815 100 103849
rect -146 103765 -112 103781
rect -146 103173 -112 103189
rect 112 103765 146 103781
rect 112 103173 146 103189
rect -100 103105 -84 103139
rect 84 103105 100 103139
rect -100 102997 -84 103031
rect 84 102997 100 103031
rect -146 102947 -112 102963
rect -146 102355 -112 102371
rect 112 102947 146 102963
rect 112 102355 146 102371
rect -100 102287 -84 102321
rect 84 102287 100 102321
rect -100 102179 -84 102213
rect 84 102179 100 102213
rect -146 102129 -112 102145
rect -146 101537 -112 101553
rect 112 102129 146 102145
rect 112 101537 146 101553
rect -100 101469 -84 101503
rect 84 101469 100 101503
rect -100 101361 -84 101395
rect 84 101361 100 101395
rect -146 101311 -112 101327
rect -146 100719 -112 100735
rect 112 101311 146 101327
rect 112 100719 146 100735
rect -100 100651 -84 100685
rect 84 100651 100 100685
rect -100 100543 -84 100577
rect 84 100543 100 100577
rect -146 100493 -112 100509
rect -146 99901 -112 99917
rect 112 100493 146 100509
rect 112 99901 146 99917
rect -100 99833 -84 99867
rect 84 99833 100 99867
rect -100 99725 -84 99759
rect 84 99725 100 99759
rect -146 99675 -112 99691
rect -146 99083 -112 99099
rect 112 99675 146 99691
rect 112 99083 146 99099
rect -100 99015 -84 99049
rect 84 99015 100 99049
rect -100 98907 -84 98941
rect 84 98907 100 98941
rect -146 98857 -112 98873
rect -146 98265 -112 98281
rect 112 98857 146 98873
rect 112 98265 146 98281
rect -100 98197 -84 98231
rect 84 98197 100 98231
rect -100 98089 -84 98123
rect 84 98089 100 98123
rect -146 98039 -112 98055
rect -146 97447 -112 97463
rect 112 98039 146 98055
rect 112 97447 146 97463
rect -100 97379 -84 97413
rect 84 97379 100 97413
rect -100 97271 -84 97305
rect 84 97271 100 97305
rect -146 97221 -112 97237
rect -146 96629 -112 96645
rect 112 97221 146 97237
rect 112 96629 146 96645
rect -100 96561 -84 96595
rect 84 96561 100 96595
rect -100 96453 -84 96487
rect 84 96453 100 96487
rect -146 96403 -112 96419
rect -146 95811 -112 95827
rect 112 96403 146 96419
rect 112 95811 146 95827
rect -100 95743 -84 95777
rect 84 95743 100 95777
rect -100 95635 -84 95669
rect 84 95635 100 95669
rect -146 95585 -112 95601
rect -146 94993 -112 95009
rect 112 95585 146 95601
rect 112 94993 146 95009
rect -100 94925 -84 94959
rect 84 94925 100 94959
rect -100 94817 -84 94851
rect 84 94817 100 94851
rect -146 94767 -112 94783
rect -146 94175 -112 94191
rect 112 94767 146 94783
rect 112 94175 146 94191
rect -100 94107 -84 94141
rect 84 94107 100 94141
rect -100 93999 -84 94033
rect 84 93999 100 94033
rect -146 93949 -112 93965
rect -146 93357 -112 93373
rect 112 93949 146 93965
rect 112 93357 146 93373
rect -100 93289 -84 93323
rect 84 93289 100 93323
rect -100 93181 -84 93215
rect 84 93181 100 93215
rect -146 93131 -112 93147
rect -146 92539 -112 92555
rect 112 93131 146 93147
rect 112 92539 146 92555
rect -100 92471 -84 92505
rect 84 92471 100 92505
rect -100 92363 -84 92397
rect 84 92363 100 92397
rect -146 92313 -112 92329
rect -146 91721 -112 91737
rect 112 92313 146 92329
rect 112 91721 146 91737
rect -100 91653 -84 91687
rect 84 91653 100 91687
rect -100 91545 -84 91579
rect 84 91545 100 91579
rect -146 91495 -112 91511
rect -146 90903 -112 90919
rect 112 91495 146 91511
rect 112 90903 146 90919
rect -100 90835 -84 90869
rect 84 90835 100 90869
rect -100 90727 -84 90761
rect 84 90727 100 90761
rect -146 90677 -112 90693
rect -146 90085 -112 90101
rect 112 90677 146 90693
rect 112 90085 146 90101
rect -100 90017 -84 90051
rect 84 90017 100 90051
rect -100 89909 -84 89943
rect 84 89909 100 89943
rect -146 89859 -112 89875
rect -146 89267 -112 89283
rect 112 89859 146 89875
rect 112 89267 146 89283
rect -100 89199 -84 89233
rect 84 89199 100 89233
rect -100 89091 -84 89125
rect 84 89091 100 89125
rect -146 89041 -112 89057
rect -146 88449 -112 88465
rect 112 89041 146 89057
rect 112 88449 146 88465
rect -100 88381 -84 88415
rect 84 88381 100 88415
rect -100 88273 -84 88307
rect 84 88273 100 88307
rect -146 88223 -112 88239
rect -146 87631 -112 87647
rect 112 88223 146 88239
rect 112 87631 146 87647
rect -100 87563 -84 87597
rect 84 87563 100 87597
rect -100 87455 -84 87489
rect 84 87455 100 87489
rect -146 87405 -112 87421
rect -146 86813 -112 86829
rect 112 87405 146 87421
rect 112 86813 146 86829
rect -100 86745 -84 86779
rect 84 86745 100 86779
rect -100 86637 -84 86671
rect 84 86637 100 86671
rect -146 86587 -112 86603
rect -146 85995 -112 86011
rect 112 86587 146 86603
rect 112 85995 146 86011
rect -100 85927 -84 85961
rect 84 85927 100 85961
rect -100 85819 -84 85853
rect 84 85819 100 85853
rect -146 85769 -112 85785
rect -146 85177 -112 85193
rect 112 85769 146 85785
rect 112 85177 146 85193
rect -100 85109 -84 85143
rect 84 85109 100 85143
rect -100 85001 -84 85035
rect 84 85001 100 85035
rect -146 84951 -112 84967
rect -146 84359 -112 84375
rect 112 84951 146 84967
rect 112 84359 146 84375
rect -100 84291 -84 84325
rect 84 84291 100 84325
rect -100 84183 -84 84217
rect 84 84183 100 84217
rect -146 84133 -112 84149
rect -146 83541 -112 83557
rect 112 84133 146 84149
rect 112 83541 146 83557
rect -100 83473 -84 83507
rect 84 83473 100 83507
rect -100 83365 -84 83399
rect 84 83365 100 83399
rect -146 83315 -112 83331
rect -146 82723 -112 82739
rect 112 83315 146 83331
rect 112 82723 146 82739
rect -100 82655 -84 82689
rect 84 82655 100 82689
rect -100 82547 -84 82581
rect 84 82547 100 82581
rect -146 82497 -112 82513
rect -146 81905 -112 81921
rect 112 82497 146 82513
rect 112 81905 146 81921
rect -100 81837 -84 81871
rect 84 81837 100 81871
rect -100 81729 -84 81763
rect 84 81729 100 81763
rect -146 81679 -112 81695
rect -146 81087 -112 81103
rect 112 81679 146 81695
rect 112 81087 146 81103
rect -100 81019 -84 81053
rect 84 81019 100 81053
rect -100 80911 -84 80945
rect 84 80911 100 80945
rect -146 80861 -112 80877
rect -146 80269 -112 80285
rect 112 80861 146 80877
rect 112 80269 146 80285
rect -100 80201 -84 80235
rect 84 80201 100 80235
rect -100 80093 -84 80127
rect 84 80093 100 80127
rect -146 80043 -112 80059
rect -146 79451 -112 79467
rect 112 80043 146 80059
rect 112 79451 146 79467
rect -100 79383 -84 79417
rect 84 79383 100 79417
rect -100 79275 -84 79309
rect 84 79275 100 79309
rect -146 79225 -112 79241
rect -146 78633 -112 78649
rect 112 79225 146 79241
rect 112 78633 146 78649
rect -100 78565 -84 78599
rect 84 78565 100 78599
rect -100 78457 -84 78491
rect 84 78457 100 78491
rect -146 78407 -112 78423
rect -146 77815 -112 77831
rect 112 78407 146 78423
rect 112 77815 146 77831
rect -100 77747 -84 77781
rect 84 77747 100 77781
rect -100 77639 -84 77673
rect 84 77639 100 77673
rect -146 77589 -112 77605
rect -146 76997 -112 77013
rect 112 77589 146 77605
rect 112 76997 146 77013
rect -100 76929 -84 76963
rect 84 76929 100 76963
rect -100 76821 -84 76855
rect 84 76821 100 76855
rect -146 76771 -112 76787
rect -146 76179 -112 76195
rect 112 76771 146 76787
rect 112 76179 146 76195
rect -100 76111 -84 76145
rect 84 76111 100 76145
rect -100 76003 -84 76037
rect 84 76003 100 76037
rect -146 75953 -112 75969
rect -146 75361 -112 75377
rect 112 75953 146 75969
rect 112 75361 146 75377
rect -100 75293 -84 75327
rect 84 75293 100 75327
rect -100 75185 -84 75219
rect 84 75185 100 75219
rect -146 75135 -112 75151
rect -146 74543 -112 74559
rect 112 75135 146 75151
rect 112 74543 146 74559
rect -100 74475 -84 74509
rect 84 74475 100 74509
rect -100 74367 -84 74401
rect 84 74367 100 74401
rect -146 74317 -112 74333
rect -146 73725 -112 73741
rect 112 74317 146 74333
rect 112 73725 146 73741
rect -100 73657 -84 73691
rect 84 73657 100 73691
rect -100 73549 -84 73583
rect 84 73549 100 73583
rect -146 73499 -112 73515
rect -146 72907 -112 72923
rect 112 73499 146 73515
rect 112 72907 146 72923
rect -100 72839 -84 72873
rect 84 72839 100 72873
rect -100 72731 -84 72765
rect 84 72731 100 72765
rect -146 72681 -112 72697
rect -146 72089 -112 72105
rect 112 72681 146 72697
rect 112 72089 146 72105
rect -100 72021 -84 72055
rect 84 72021 100 72055
rect -100 71913 -84 71947
rect 84 71913 100 71947
rect -146 71863 -112 71879
rect -146 71271 -112 71287
rect 112 71863 146 71879
rect 112 71271 146 71287
rect -100 71203 -84 71237
rect 84 71203 100 71237
rect -100 71095 -84 71129
rect 84 71095 100 71129
rect -146 71045 -112 71061
rect -146 70453 -112 70469
rect 112 71045 146 71061
rect 112 70453 146 70469
rect -100 70385 -84 70419
rect 84 70385 100 70419
rect -100 70277 -84 70311
rect 84 70277 100 70311
rect -146 70227 -112 70243
rect -146 69635 -112 69651
rect 112 70227 146 70243
rect 112 69635 146 69651
rect -100 69567 -84 69601
rect 84 69567 100 69601
rect -100 69459 -84 69493
rect 84 69459 100 69493
rect -146 69409 -112 69425
rect -146 68817 -112 68833
rect 112 69409 146 69425
rect 112 68817 146 68833
rect -100 68749 -84 68783
rect 84 68749 100 68783
rect -100 68641 -84 68675
rect 84 68641 100 68675
rect -146 68591 -112 68607
rect -146 67999 -112 68015
rect 112 68591 146 68607
rect 112 67999 146 68015
rect -100 67931 -84 67965
rect 84 67931 100 67965
rect -100 67823 -84 67857
rect 84 67823 100 67857
rect -146 67773 -112 67789
rect -146 67181 -112 67197
rect 112 67773 146 67789
rect 112 67181 146 67197
rect -100 67113 -84 67147
rect 84 67113 100 67147
rect -100 67005 -84 67039
rect 84 67005 100 67039
rect -146 66955 -112 66971
rect -146 66363 -112 66379
rect 112 66955 146 66971
rect 112 66363 146 66379
rect -100 66295 -84 66329
rect 84 66295 100 66329
rect -100 66187 -84 66221
rect 84 66187 100 66221
rect -146 66137 -112 66153
rect -146 65545 -112 65561
rect 112 66137 146 66153
rect 112 65545 146 65561
rect -100 65477 -84 65511
rect 84 65477 100 65511
rect -100 65369 -84 65403
rect 84 65369 100 65403
rect -146 65319 -112 65335
rect -146 64727 -112 64743
rect 112 65319 146 65335
rect 112 64727 146 64743
rect -100 64659 -84 64693
rect 84 64659 100 64693
rect -100 64551 -84 64585
rect 84 64551 100 64585
rect -146 64501 -112 64517
rect -146 63909 -112 63925
rect 112 64501 146 64517
rect 112 63909 146 63925
rect -100 63841 -84 63875
rect 84 63841 100 63875
rect -100 63733 -84 63767
rect 84 63733 100 63767
rect -146 63683 -112 63699
rect -146 63091 -112 63107
rect 112 63683 146 63699
rect 112 63091 146 63107
rect -100 63023 -84 63057
rect 84 63023 100 63057
rect -100 62915 -84 62949
rect 84 62915 100 62949
rect -146 62865 -112 62881
rect -146 62273 -112 62289
rect 112 62865 146 62881
rect 112 62273 146 62289
rect -100 62205 -84 62239
rect 84 62205 100 62239
rect -100 62097 -84 62131
rect 84 62097 100 62131
rect -146 62047 -112 62063
rect -146 61455 -112 61471
rect 112 62047 146 62063
rect 112 61455 146 61471
rect -100 61387 -84 61421
rect 84 61387 100 61421
rect -100 61279 -84 61313
rect 84 61279 100 61313
rect -146 61229 -112 61245
rect -146 60637 -112 60653
rect 112 61229 146 61245
rect 112 60637 146 60653
rect -100 60569 -84 60603
rect 84 60569 100 60603
rect -100 60461 -84 60495
rect 84 60461 100 60495
rect -146 60411 -112 60427
rect -146 59819 -112 59835
rect 112 60411 146 60427
rect 112 59819 146 59835
rect -100 59751 -84 59785
rect 84 59751 100 59785
rect -100 59643 -84 59677
rect 84 59643 100 59677
rect -146 59593 -112 59609
rect -146 59001 -112 59017
rect 112 59593 146 59609
rect 112 59001 146 59017
rect -100 58933 -84 58967
rect 84 58933 100 58967
rect -100 58825 -84 58859
rect 84 58825 100 58859
rect -146 58775 -112 58791
rect -146 58183 -112 58199
rect 112 58775 146 58791
rect 112 58183 146 58199
rect -100 58115 -84 58149
rect 84 58115 100 58149
rect -100 58007 -84 58041
rect 84 58007 100 58041
rect -146 57957 -112 57973
rect -146 57365 -112 57381
rect 112 57957 146 57973
rect 112 57365 146 57381
rect -100 57297 -84 57331
rect 84 57297 100 57331
rect -100 57189 -84 57223
rect 84 57189 100 57223
rect -146 57139 -112 57155
rect -146 56547 -112 56563
rect 112 57139 146 57155
rect 112 56547 146 56563
rect -100 56479 -84 56513
rect 84 56479 100 56513
rect -100 56371 -84 56405
rect 84 56371 100 56405
rect -146 56321 -112 56337
rect -146 55729 -112 55745
rect 112 56321 146 56337
rect 112 55729 146 55745
rect -100 55661 -84 55695
rect 84 55661 100 55695
rect -100 55553 -84 55587
rect 84 55553 100 55587
rect -146 55503 -112 55519
rect -146 54911 -112 54927
rect 112 55503 146 55519
rect 112 54911 146 54927
rect -100 54843 -84 54877
rect 84 54843 100 54877
rect -100 54735 -84 54769
rect 84 54735 100 54769
rect -146 54685 -112 54701
rect -146 54093 -112 54109
rect 112 54685 146 54701
rect 112 54093 146 54109
rect -100 54025 -84 54059
rect 84 54025 100 54059
rect -100 53917 -84 53951
rect 84 53917 100 53951
rect -146 53867 -112 53883
rect -146 53275 -112 53291
rect 112 53867 146 53883
rect 112 53275 146 53291
rect -100 53207 -84 53241
rect 84 53207 100 53241
rect -100 53099 -84 53133
rect 84 53099 100 53133
rect -146 53049 -112 53065
rect -146 52457 -112 52473
rect 112 53049 146 53065
rect 112 52457 146 52473
rect -100 52389 -84 52423
rect 84 52389 100 52423
rect -100 52281 -84 52315
rect 84 52281 100 52315
rect -146 52231 -112 52247
rect -146 51639 -112 51655
rect 112 52231 146 52247
rect 112 51639 146 51655
rect -100 51571 -84 51605
rect 84 51571 100 51605
rect -100 51463 -84 51497
rect 84 51463 100 51497
rect -146 51413 -112 51429
rect -146 50821 -112 50837
rect 112 51413 146 51429
rect 112 50821 146 50837
rect -100 50753 -84 50787
rect 84 50753 100 50787
rect -100 50645 -84 50679
rect 84 50645 100 50679
rect -146 50595 -112 50611
rect -146 50003 -112 50019
rect 112 50595 146 50611
rect 112 50003 146 50019
rect -100 49935 -84 49969
rect 84 49935 100 49969
rect -100 49827 -84 49861
rect 84 49827 100 49861
rect -146 49777 -112 49793
rect -146 49185 -112 49201
rect 112 49777 146 49793
rect 112 49185 146 49201
rect -100 49117 -84 49151
rect 84 49117 100 49151
rect -100 49009 -84 49043
rect 84 49009 100 49043
rect -146 48959 -112 48975
rect -146 48367 -112 48383
rect 112 48959 146 48975
rect 112 48367 146 48383
rect -100 48299 -84 48333
rect 84 48299 100 48333
rect -100 48191 -84 48225
rect 84 48191 100 48225
rect -146 48141 -112 48157
rect -146 47549 -112 47565
rect 112 48141 146 48157
rect 112 47549 146 47565
rect -100 47481 -84 47515
rect 84 47481 100 47515
rect -100 47373 -84 47407
rect 84 47373 100 47407
rect -146 47323 -112 47339
rect -146 46731 -112 46747
rect 112 47323 146 47339
rect 112 46731 146 46747
rect -100 46663 -84 46697
rect 84 46663 100 46697
rect -100 46555 -84 46589
rect 84 46555 100 46589
rect -146 46505 -112 46521
rect -146 45913 -112 45929
rect 112 46505 146 46521
rect 112 45913 146 45929
rect -100 45845 -84 45879
rect 84 45845 100 45879
rect -100 45737 -84 45771
rect 84 45737 100 45771
rect -146 45687 -112 45703
rect -146 45095 -112 45111
rect 112 45687 146 45703
rect 112 45095 146 45111
rect -100 45027 -84 45061
rect 84 45027 100 45061
rect -100 44919 -84 44953
rect 84 44919 100 44953
rect -146 44869 -112 44885
rect -146 44277 -112 44293
rect 112 44869 146 44885
rect 112 44277 146 44293
rect -100 44209 -84 44243
rect 84 44209 100 44243
rect -100 44101 -84 44135
rect 84 44101 100 44135
rect -146 44051 -112 44067
rect -146 43459 -112 43475
rect 112 44051 146 44067
rect 112 43459 146 43475
rect -100 43391 -84 43425
rect 84 43391 100 43425
rect -100 43283 -84 43317
rect 84 43283 100 43317
rect -146 43233 -112 43249
rect -146 42641 -112 42657
rect 112 43233 146 43249
rect 112 42641 146 42657
rect -100 42573 -84 42607
rect 84 42573 100 42607
rect -100 42465 -84 42499
rect 84 42465 100 42499
rect -146 42415 -112 42431
rect -146 41823 -112 41839
rect 112 42415 146 42431
rect 112 41823 146 41839
rect -100 41755 -84 41789
rect 84 41755 100 41789
rect -100 41647 -84 41681
rect 84 41647 100 41681
rect -146 41597 -112 41613
rect -146 41005 -112 41021
rect 112 41597 146 41613
rect 112 41005 146 41021
rect -100 40937 -84 40971
rect 84 40937 100 40971
rect -100 40829 -84 40863
rect 84 40829 100 40863
rect -146 40779 -112 40795
rect -146 40187 -112 40203
rect 112 40779 146 40795
rect 112 40187 146 40203
rect -100 40119 -84 40153
rect 84 40119 100 40153
rect -100 40011 -84 40045
rect 84 40011 100 40045
rect -146 39961 -112 39977
rect -146 39369 -112 39385
rect 112 39961 146 39977
rect 112 39369 146 39385
rect -100 39301 -84 39335
rect 84 39301 100 39335
rect -100 39193 -84 39227
rect 84 39193 100 39227
rect -146 39143 -112 39159
rect -146 38551 -112 38567
rect 112 39143 146 39159
rect 112 38551 146 38567
rect -100 38483 -84 38517
rect 84 38483 100 38517
rect -100 38375 -84 38409
rect 84 38375 100 38409
rect -146 38325 -112 38341
rect -146 37733 -112 37749
rect 112 38325 146 38341
rect 112 37733 146 37749
rect -100 37665 -84 37699
rect 84 37665 100 37699
rect -100 37557 -84 37591
rect 84 37557 100 37591
rect -146 37507 -112 37523
rect -146 36915 -112 36931
rect 112 37507 146 37523
rect 112 36915 146 36931
rect -100 36847 -84 36881
rect 84 36847 100 36881
rect -100 36739 -84 36773
rect 84 36739 100 36773
rect -146 36689 -112 36705
rect -146 36097 -112 36113
rect 112 36689 146 36705
rect 112 36097 146 36113
rect -100 36029 -84 36063
rect 84 36029 100 36063
rect -100 35921 -84 35955
rect 84 35921 100 35955
rect -146 35871 -112 35887
rect -146 35279 -112 35295
rect 112 35871 146 35887
rect 112 35279 146 35295
rect -100 35211 -84 35245
rect 84 35211 100 35245
rect -100 35103 -84 35137
rect 84 35103 100 35137
rect -146 35053 -112 35069
rect -146 34461 -112 34477
rect 112 35053 146 35069
rect 112 34461 146 34477
rect -100 34393 -84 34427
rect 84 34393 100 34427
rect -100 34285 -84 34319
rect 84 34285 100 34319
rect -146 34235 -112 34251
rect -146 33643 -112 33659
rect 112 34235 146 34251
rect 112 33643 146 33659
rect -100 33575 -84 33609
rect 84 33575 100 33609
rect -100 33467 -84 33501
rect 84 33467 100 33501
rect -146 33417 -112 33433
rect -146 32825 -112 32841
rect 112 33417 146 33433
rect 112 32825 146 32841
rect -100 32757 -84 32791
rect 84 32757 100 32791
rect -100 32649 -84 32683
rect 84 32649 100 32683
rect -146 32599 -112 32615
rect -146 32007 -112 32023
rect 112 32599 146 32615
rect 112 32007 146 32023
rect -100 31939 -84 31973
rect 84 31939 100 31973
rect -100 31831 -84 31865
rect 84 31831 100 31865
rect -146 31781 -112 31797
rect -146 31189 -112 31205
rect 112 31781 146 31797
rect 112 31189 146 31205
rect -100 31121 -84 31155
rect 84 31121 100 31155
rect -100 31013 -84 31047
rect 84 31013 100 31047
rect -146 30963 -112 30979
rect -146 30371 -112 30387
rect 112 30963 146 30979
rect 112 30371 146 30387
rect -100 30303 -84 30337
rect 84 30303 100 30337
rect -100 30195 -84 30229
rect 84 30195 100 30229
rect -146 30145 -112 30161
rect -146 29553 -112 29569
rect 112 30145 146 30161
rect 112 29553 146 29569
rect -100 29485 -84 29519
rect 84 29485 100 29519
rect -100 29377 -84 29411
rect 84 29377 100 29411
rect -146 29327 -112 29343
rect -146 28735 -112 28751
rect 112 29327 146 29343
rect 112 28735 146 28751
rect -100 28667 -84 28701
rect 84 28667 100 28701
rect -100 28559 -84 28593
rect 84 28559 100 28593
rect -146 28509 -112 28525
rect -146 27917 -112 27933
rect 112 28509 146 28525
rect 112 27917 146 27933
rect -100 27849 -84 27883
rect 84 27849 100 27883
rect -100 27741 -84 27775
rect 84 27741 100 27775
rect -146 27691 -112 27707
rect -146 27099 -112 27115
rect 112 27691 146 27707
rect 112 27099 146 27115
rect -100 27031 -84 27065
rect 84 27031 100 27065
rect -100 26923 -84 26957
rect 84 26923 100 26957
rect -146 26873 -112 26889
rect -146 26281 -112 26297
rect 112 26873 146 26889
rect 112 26281 146 26297
rect -100 26213 -84 26247
rect 84 26213 100 26247
rect -100 26105 -84 26139
rect 84 26105 100 26139
rect -146 26055 -112 26071
rect -146 25463 -112 25479
rect 112 26055 146 26071
rect 112 25463 146 25479
rect -100 25395 -84 25429
rect 84 25395 100 25429
rect -100 25287 -84 25321
rect 84 25287 100 25321
rect -146 25237 -112 25253
rect -146 24645 -112 24661
rect 112 25237 146 25253
rect 112 24645 146 24661
rect -100 24577 -84 24611
rect 84 24577 100 24611
rect -100 24469 -84 24503
rect 84 24469 100 24503
rect -146 24419 -112 24435
rect -146 23827 -112 23843
rect 112 24419 146 24435
rect 112 23827 146 23843
rect -100 23759 -84 23793
rect 84 23759 100 23793
rect -100 23651 -84 23685
rect 84 23651 100 23685
rect -146 23601 -112 23617
rect -146 23009 -112 23025
rect 112 23601 146 23617
rect 112 23009 146 23025
rect -100 22941 -84 22975
rect 84 22941 100 22975
rect -100 22833 -84 22867
rect 84 22833 100 22867
rect -146 22783 -112 22799
rect -146 22191 -112 22207
rect 112 22783 146 22799
rect 112 22191 146 22207
rect -100 22123 -84 22157
rect 84 22123 100 22157
rect -100 22015 -84 22049
rect 84 22015 100 22049
rect -146 21965 -112 21981
rect -146 21373 -112 21389
rect 112 21965 146 21981
rect 112 21373 146 21389
rect -100 21305 -84 21339
rect 84 21305 100 21339
rect -100 21197 -84 21231
rect 84 21197 100 21231
rect -146 21147 -112 21163
rect -146 20555 -112 20571
rect 112 21147 146 21163
rect 112 20555 146 20571
rect -100 20487 -84 20521
rect 84 20487 100 20521
rect -100 20379 -84 20413
rect 84 20379 100 20413
rect -146 20329 -112 20345
rect -146 19737 -112 19753
rect 112 20329 146 20345
rect 112 19737 146 19753
rect -100 19669 -84 19703
rect 84 19669 100 19703
rect -100 19561 -84 19595
rect 84 19561 100 19595
rect -146 19511 -112 19527
rect -146 18919 -112 18935
rect 112 19511 146 19527
rect 112 18919 146 18935
rect -100 18851 -84 18885
rect 84 18851 100 18885
rect -100 18743 -84 18777
rect 84 18743 100 18777
rect -146 18693 -112 18709
rect -146 18101 -112 18117
rect 112 18693 146 18709
rect 112 18101 146 18117
rect -100 18033 -84 18067
rect 84 18033 100 18067
rect -100 17925 -84 17959
rect 84 17925 100 17959
rect -146 17875 -112 17891
rect -146 17283 -112 17299
rect 112 17875 146 17891
rect 112 17283 146 17299
rect -100 17215 -84 17249
rect 84 17215 100 17249
rect -100 17107 -84 17141
rect 84 17107 100 17141
rect -146 17057 -112 17073
rect -146 16465 -112 16481
rect 112 17057 146 17073
rect 112 16465 146 16481
rect -100 16397 -84 16431
rect 84 16397 100 16431
rect -100 16289 -84 16323
rect 84 16289 100 16323
rect -146 16239 -112 16255
rect -146 15647 -112 15663
rect 112 16239 146 16255
rect 112 15647 146 15663
rect -100 15579 -84 15613
rect 84 15579 100 15613
rect -100 15471 -84 15505
rect 84 15471 100 15505
rect -146 15421 -112 15437
rect -146 14829 -112 14845
rect 112 15421 146 15437
rect 112 14829 146 14845
rect -100 14761 -84 14795
rect 84 14761 100 14795
rect -100 14653 -84 14687
rect 84 14653 100 14687
rect -146 14603 -112 14619
rect -146 14011 -112 14027
rect 112 14603 146 14619
rect 112 14011 146 14027
rect -100 13943 -84 13977
rect 84 13943 100 13977
rect -100 13835 -84 13869
rect 84 13835 100 13869
rect -146 13785 -112 13801
rect -146 13193 -112 13209
rect 112 13785 146 13801
rect 112 13193 146 13209
rect -100 13125 -84 13159
rect 84 13125 100 13159
rect -100 13017 -84 13051
rect 84 13017 100 13051
rect -146 12967 -112 12983
rect -146 12375 -112 12391
rect 112 12967 146 12983
rect 112 12375 146 12391
rect -100 12307 -84 12341
rect 84 12307 100 12341
rect -100 12199 -84 12233
rect 84 12199 100 12233
rect -146 12149 -112 12165
rect -146 11557 -112 11573
rect 112 12149 146 12165
rect 112 11557 146 11573
rect -100 11489 -84 11523
rect 84 11489 100 11523
rect -100 11381 -84 11415
rect 84 11381 100 11415
rect -146 11331 -112 11347
rect -146 10739 -112 10755
rect 112 11331 146 11347
rect 112 10739 146 10755
rect -100 10671 -84 10705
rect 84 10671 100 10705
rect -100 10563 -84 10597
rect 84 10563 100 10597
rect -146 10513 -112 10529
rect -146 9921 -112 9937
rect 112 10513 146 10529
rect 112 9921 146 9937
rect -100 9853 -84 9887
rect 84 9853 100 9887
rect -100 9745 -84 9779
rect 84 9745 100 9779
rect -146 9695 -112 9711
rect -146 9103 -112 9119
rect 112 9695 146 9711
rect 112 9103 146 9119
rect -100 9035 -84 9069
rect 84 9035 100 9069
rect -100 8927 -84 8961
rect 84 8927 100 8961
rect -146 8877 -112 8893
rect -146 8285 -112 8301
rect 112 8877 146 8893
rect 112 8285 146 8301
rect -100 8217 -84 8251
rect 84 8217 100 8251
rect -100 8109 -84 8143
rect 84 8109 100 8143
rect -146 8059 -112 8075
rect -146 7467 -112 7483
rect 112 8059 146 8075
rect 112 7467 146 7483
rect -100 7399 -84 7433
rect 84 7399 100 7433
rect -100 7291 -84 7325
rect 84 7291 100 7325
rect -146 7241 -112 7257
rect -146 6649 -112 6665
rect 112 7241 146 7257
rect 112 6649 146 6665
rect -100 6581 -84 6615
rect 84 6581 100 6615
rect -100 6473 -84 6507
rect 84 6473 100 6507
rect -146 6423 -112 6439
rect -146 5831 -112 5847
rect 112 6423 146 6439
rect 112 5831 146 5847
rect -100 5763 -84 5797
rect 84 5763 100 5797
rect -100 5655 -84 5689
rect 84 5655 100 5689
rect -146 5605 -112 5621
rect -146 5013 -112 5029
rect 112 5605 146 5621
rect 112 5013 146 5029
rect -100 4945 -84 4979
rect 84 4945 100 4979
rect -100 4837 -84 4871
rect 84 4837 100 4871
rect -146 4787 -112 4803
rect -146 4195 -112 4211
rect 112 4787 146 4803
rect 112 4195 146 4211
rect -100 4127 -84 4161
rect 84 4127 100 4161
rect -100 4019 -84 4053
rect 84 4019 100 4053
rect -146 3969 -112 3985
rect -146 3377 -112 3393
rect 112 3969 146 3985
rect 112 3377 146 3393
rect -100 3309 -84 3343
rect 84 3309 100 3343
rect -100 3201 -84 3235
rect 84 3201 100 3235
rect -146 3151 -112 3167
rect -146 2559 -112 2575
rect 112 3151 146 3167
rect 112 2559 146 2575
rect -100 2491 -84 2525
rect 84 2491 100 2525
rect -100 2383 -84 2417
rect 84 2383 100 2417
rect -146 2333 -112 2349
rect -146 1741 -112 1757
rect 112 2333 146 2349
rect 112 1741 146 1757
rect -100 1673 -84 1707
rect 84 1673 100 1707
rect -100 1565 -84 1599
rect 84 1565 100 1599
rect -146 1515 -112 1531
rect -146 923 -112 939
rect 112 1515 146 1531
rect 112 923 146 939
rect -100 855 -84 889
rect 84 855 100 889
rect -100 747 -84 781
rect 84 747 100 781
rect -146 697 -112 713
rect -146 105 -112 121
rect 112 697 146 713
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -713 -112 -697
rect 112 -121 146 -105
rect 112 -713 146 -697
rect -100 -781 -84 -747
rect 84 -781 100 -747
rect -100 -889 -84 -855
rect 84 -889 100 -855
rect -146 -939 -112 -923
rect -146 -1531 -112 -1515
rect 112 -939 146 -923
rect 112 -1531 146 -1515
rect -100 -1599 -84 -1565
rect 84 -1599 100 -1565
rect -100 -1707 -84 -1673
rect 84 -1707 100 -1673
rect -146 -1757 -112 -1741
rect -146 -2349 -112 -2333
rect 112 -1757 146 -1741
rect 112 -2349 146 -2333
rect -100 -2417 -84 -2383
rect 84 -2417 100 -2383
rect -100 -2525 -84 -2491
rect 84 -2525 100 -2491
rect -146 -2575 -112 -2559
rect -146 -3167 -112 -3151
rect 112 -2575 146 -2559
rect 112 -3167 146 -3151
rect -100 -3235 -84 -3201
rect 84 -3235 100 -3201
rect -100 -3343 -84 -3309
rect 84 -3343 100 -3309
rect -146 -3393 -112 -3377
rect -146 -3985 -112 -3969
rect 112 -3393 146 -3377
rect 112 -3985 146 -3969
rect -100 -4053 -84 -4019
rect 84 -4053 100 -4019
rect -100 -4161 -84 -4127
rect 84 -4161 100 -4127
rect -146 -4211 -112 -4195
rect -146 -4803 -112 -4787
rect 112 -4211 146 -4195
rect 112 -4803 146 -4787
rect -100 -4871 -84 -4837
rect 84 -4871 100 -4837
rect -100 -4979 -84 -4945
rect 84 -4979 100 -4945
rect -146 -5029 -112 -5013
rect -146 -5621 -112 -5605
rect 112 -5029 146 -5013
rect 112 -5621 146 -5605
rect -100 -5689 -84 -5655
rect 84 -5689 100 -5655
rect -100 -5797 -84 -5763
rect 84 -5797 100 -5763
rect -146 -5847 -112 -5831
rect -146 -6439 -112 -6423
rect 112 -5847 146 -5831
rect 112 -6439 146 -6423
rect -100 -6507 -84 -6473
rect 84 -6507 100 -6473
rect -100 -6615 -84 -6581
rect 84 -6615 100 -6581
rect -146 -6665 -112 -6649
rect -146 -7257 -112 -7241
rect 112 -6665 146 -6649
rect 112 -7257 146 -7241
rect -100 -7325 -84 -7291
rect 84 -7325 100 -7291
rect -100 -7433 -84 -7399
rect 84 -7433 100 -7399
rect -146 -7483 -112 -7467
rect -146 -8075 -112 -8059
rect 112 -7483 146 -7467
rect 112 -8075 146 -8059
rect -100 -8143 -84 -8109
rect 84 -8143 100 -8109
rect -100 -8251 -84 -8217
rect 84 -8251 100 -8217
rect -146 -8301 -112 -8285
rect -146 -8893 -112 -8877
rect 112 -8301 146 -8285
rect 112 -8893 146 -8877
rect -100 -8961 -84 -8927
rect 84 -8961 100 -8927
rect -100 -9069 -84 -9035
rect 84 -9069 100 -9035
rect -146 -9119 -112 -9103
rect -146 -9711 -112 -9695
rect 112 -9119 146 -9103
rect 112 -9711 146 -9695
rect -100 -9779 -84 -9745
rect 84 -9779 100 -9745
rect -100 -9887 -84 -9853
rect 84 -9887 100 -9853
rect -146 -9937 -112 -9921
rect -146 -10529 -112 -10513
rect 112 -9937 146 -9921
rect 112 -10529 146 -10513
rect -100 -10597 -84 -10563
rect 84 -10597 100 -10563
rect -100 -10705 -84 -10671
rect 84 -10705 100 -10671
rect -146 -10755 -112 -10739
rect -146 -11347 -112 -11331
rect 112 -10755 146 -10739
rect 112 -11347 146 -11331
rect -100 -11415 -84 -11381
rect 84 -11415 100 -11381
rect -100 -11523 -84 -11489
rect 84 -11523 100 -11489
rect -146 -11573 -112 -11557
rect -146 -12165 -112 -12149
rect 112 -11573 146 -11557
rect 112 -12165 146 -12149
rect -100 -12233 -84 -12199
rect 84 -12233 100 -12199
rect -100 -12341 -84 -12307
rect 84 -12341 100 -12307
rect -146 -12391 -112 -12375
rect -146 -12983 -112 -12967
rect 112 -12391 146 -12375
rect 112 -12983 146 -12967
rect -100 -13051 -84 -13017
rect 84 -13051 100 -13017
rect -100 -13159 -84 -13125
rect 84 -13159 100 -13125
rect -146 -13209 -112 -13193
rect -146 -13801 -112 -13785
rect 112 -13209 146 -13193
rect 112 -13801 146 -13785
rect -100 -13869 -84 -13835
rect 84 -13869 100 -13835
rect -100 -13977 -84 -13943
rect 84 -13977 100 -13943
rect -146 -14027 -112 -14011
rect -146 -14619 -112 -14603
rect 112 -14027 146 -14011
rect 112 -14619 146 -14603
rect -100 -14687 -84 -14653
rect 84 -14687 100 -14653
rect -100 -14795 -84 -14761
rect 84 -14795 100 -14761
rect -146 -14845 -112 -14829
rect -146 -15437 -112 -15421
rect 112 -14845 146 -14829
rect 112 -15437 146 -15421
rect -100 -15505 -84 -15471
rect 84 -15505 100 -15471
rect -100 -15613 -84 -15579
rect 84 -15613 100 -15579
rect -146 -15663 -112 -15647
rect -146 -16255 -112 -16239
rect 112 -15663 146 -15647
rect 112 -16255 146 -16239
rect -100 -16323 -84 -16289
rect 84 -16323 100 -16289
rect -100 -16431 -84 -16397
rect 84 -16431 100 -16397
rect -146 -16481 -112 -16465
rect -146 -17073 -112 -17057
rect 112 -16481 146 -16465
rect 112 -17073 146 -17057
rect -100 -17141 -84 -17107
rect 84 -17141 100 -17107
rect -100 -17249 -84 -17215
rect 84 -17249 100 -17215
rect -146 -17299 -112 -17283
rect -146 -17891 -112 -17875
rect 112 -17299 146 -17283
rect 112 -17891 146 -17875
rect -100 -17959 -84 -17925
rect 84 -17959 100 -17925
rect -100 -18067 -84 -18033
rect 84 -18067 100 -18033
rect -146 -18117 -112 -18101
rect -146 -18709 -112 -18693
rect 112 -18117 146 -18101
rect 112 -18709 146 -18693
rect -100 -18777 -84 -18743
rect 84 -18777 100 -18743
rect -100 -18885 -84 -18851
rect 84 -18885 100 -18851
rect -146 -18935 -112 -18919
rect -146 -19527 -112 -19511
rect 112 -18935 146 -18919
rect 112 -19527 146 -19511
rect -100 -19595 -84 -19561
rect 84 -19595 100 -19561
rect -100 -19703 -84 -19669
rect 84 -19703 100 -19669
rect -146 -19753 -112 -19737
rect -146 -20345 -112 -20329
rect 112 -19753 146 -19737
rect 112 -20345 146 -20329
rect -100 -20413 -84 -20379
rect 84 -20413 100 -20379
rect -100 -20521 -84 -20487
rect 84 -20521 100 -20487
rect -146 -20571 -112 -20555
rect -146 -21163 -112 -21147
rect 112 -20571 146 -20555
rect 112 -21163 146 -21147
rect -100 -21231 -84 -21197
rect 84 -21231 100 -21197
rect -100 -21339 -84 -21305
rect 84 -21339 100 -21305
rect -146 -21389 -112 -21373
rect -146 -21981 -112 -21965
rect 112 -21389 146 -21373
rect 112 -21981 146 -21965
rect -100 -22049 -84 -22015
rect 84 -22049 100 -22015
rect -100 -22157 -84 -22123
rect 84 -22157 100 -22123
rect -146 -22207 -112 -22191
rect -146 -22799 -112 -22783
rect 112 -22207 146 -22191
rect 112 -22799 146 -22783
rect -100 -22867 -84 -22833
rect 84 -22867 100 -22833
rect -100 -22975 -84 -22941
rect 84 -22975 100 -22941
rect -146 -23025 -112 -23009
rect -146 -23617 -112 -23601
rect 112 -23025 146 -23009
rect 112 -23617 146 -23601
rect -100 -23685 -84 -23651
rect 84 -23685 100 -23651
rect -100 -23793 -84 -23759
rect 84 -23793 100 -23759
rect -146 -23843 -112 -23827
rect -146 -24435 -112 -24419
rect 112 -23843 146 -23827
rect 112 -24435 146 -24419
rect -100 -24503 -84 -24469
rect 84 -24503 100 -24469
rect -100 -24611 -84 -24577
rect 84 -24611 100 -24577
rect -146 -24661 -112 -24645
rect -146 -25253 -112 -25237
rect 112 -24661 146 -24645
rect 112 -25253 146 -25237
rect -100 -25321 -84 -25287
rect 84 -25321 100 -25287
rect -100 -25429 -84 -25395
rect 84 -25429 100 -25395
rect -146 -25479 -112 -25463
rect -146 -26071 -112 -26055
rect 112 -25479 146 -25463
rect 112 -26071 146 -26055
rect -100 -26139 -84 -26105
rect 84 -26139 100 -26105
rect -100 -26247 -84 -26213
rect 84 -26247 100 -26213
rect -146 -26297 -112 -26281
rect -146 -26889 -112 -26873
rect 112 -26297 146 -26281
rect 112 -26889 146 -26873
rect -100 -26957 -84 -26923
rect 84 -26957 100 -26923
rect -100 -27065 -84 -27031
rect 84 -27065 100 -27031
rect -146 -27115 -112 -27099
rect -146 -27707 -112 -27691
rect 112 -27115 146 -27099
rect 112 -27707 146 -27691
rect -100 -27775 -84 -27741
rect 84 -27775 100 -27741
rect -100 -27883 -84 -27849
rect 84 -27883 100 -27849
rect -146 -27933 -112 -27917
rect -146 -28525 -112 -28509
rect 112 -27933 146 -27917
rect 112 -28525 146 -28509
rect -100 -28593 -84 -28559
rect 84 -28593 100 -28559
rect -100 -28701 -84 -28667
rect 84 -28701 100 -28667
rect -146 -28751 -112 -28735
rect -146 -29343 -112 -29327
rect 112 -28751 146 -28735
rect 112 -29343 146 -29327
rect -100 -29411 -84 -29377
rect 84 -29411 100 -29377
rect -100 -29519 -84 -29485
rect 84 -29519 100 -29485
rect -146 -29569 -112 -29553
rect -146 -30161 -112 -30145
rect 112 -29569 146 -29553
rect 112 -30161 146 -30145
rect -100 -30229 -84 -30195
rect 84 -30229 100 -30195
rect -100 -30337 -84 -30303
rect 84 -30337 100 -30303
rect -146 -30387 -112 -30371
rect -146 -30979 -112 -30963
rect 112 -30387 146 -30371
rect 112 -30979 146 -30963
rect -100 -31047 -84 -31013
rect 84 -31047 100 -31013
rect -100 -31155 -84 -31121
rect 84 -31155 100 -31121
rect -146 -31205 -112 -31189
rect -146 -31797 -112 -31781
rect 112 -31205 146 -31189
rect 112 -31797 146 -31781
rect -100 -31865 -84 -31831
rect 84 -31865 100 -31831
rect -100 -31973 -84 -31939
rect 84 -31973 100 -31939
rect -146 -32023 -112 -32007
rect -146 -32615 -112 -32599
rect 112 -32023 146 -32007
rect 112 -32615 146 -32599
rect -100 -32683 -84 -32649
rect 84 -32683 100 -32649
rect -100 -32791 -84 -32757
rect 84 -32791 100 -32757
rect -146 -32841 -112 -32825
rect -146 -33433 -112 -33417
rect 112 -32841 146 -32825
rect 112 -33433 146 -33417
rect -100 -33501 -84 -33467
rect 84 -33501 100 -33467
rect -100 -33609 -84 -33575
rect 84 -33609 100 -33575
rect -146 -33659 -112 -33643
rect -146 -34251 -112 -34235
rect 112 -33659 146 -33643
rect 112 -34251 146 -34235
rect -100 -34319 -84 -34285
rect 84 -34319 100 -34285
rect -100 -34427 -84 -34393
rect 84 -34427 100 -34393
rect -146 -34477 -112 -34461
rect -146 -35069 -112 -35053
rect 112 -34477 146 -34461
rect 112 -35069 146 -35053
rect -100 -35137 -84 -35103
rect 84 -35137 100 -35103
rect -100 -35245 -84 -35211
rect 84 -35245 100 -35211
rect -146 -35295 -112 -35279
rect -146 -35887 -112 -35871
rect 112 -35295 146 -35279
rect 112 -35887 146 -35871
rect -100 -35955 -84 -35921
rect 84 -35955 100 -35921
rect -100 -36063 -84 -36029
rect 84 -36063 100 -36029
rect -146 -36113 -112 -36097
rect -146 -36705 -112 -36689
rect 112 -36113 146 -36097
rect 112 -36705 146 -36689
rect -100 -36773 -84 -36739
rect 84 -36773 100 -36739
rect -100 -36881 -84 -36847
rect 84 -36881 100 -36847
rect -146 -36931 -112 -36915
rect -146 -37523 -112 -37507
rect 112 -36931 146 -36915
rect 112 -37523 146 -37507
rect -100 -37591 -84 -37557
rect 84 -37591 100 -37557
rect -100 -37699 -84 -37665
rect 84 -37699 100 -37665
rect -146 -37749 -112 -37733
rect -146 -38341 -112 -38325
rect 112 -37749 146 -37733
rect 112 -38341 146 -38325
rect -100 -38409 -84 -38375
rect 84 -38409 100 -38375
rect -100 -38517 -84 -38483
rect 84 -38517 100 -38483
rect -146 -38567 -112 -38551
rect -146 -39159 -112 -39143
rect 112 -38567 146 -38551
rect 112 -39159 146 -39143
rect -100 -39227 -84 -39193
rect 84 -39227 100 -39193
rect -100 -39335 -84 -39301
rect 84 -39335 100 -39301
rect -146 -39385 -112 -39369
rect -146 -39977 -112 -39961
rect 112 -39385 146 -39369
rect 112 -39977 146 -39961
rect -100 -40045 -84 -40011
rect 84 -40045 100 -40011
rect -100 -40153 -84 -40119
rect 84 -40153 100 -40119
rect -146 -40203 -112 -40187
rect -146 -40795 -112 -40779
rect 112 -40203 146 -40187
rect 112 -40795 146 -40779
rect -100 -40863 -84 -40829
rect 84 -40863 100 -40829
rect -100 -40971 -84 -40937
rect 84 -40971 100 -40937
rect -146 -41021 -112 -41005
rect -146 -41613 -112 -41597
rect 112 -41021 146 -41005
rect 112 -41613 146 -41597
rect -100 -41681 -84 -41647
rect 84 -41681 100 -41647
rect -100 -41789 -84 -41755
rect 84 -41789 100 -41755
rect -146 -41839 -112 -41823
rect -146 -42431 -112 -42415
rect 112 -41839 146 -41823
rect 112 -42431 146 -42415
rect -100 -42499 -84 -42465
rect 84 -42499 100 -42465
rect -100 -42607 -84 -42573
rect 84 -42607 100 -42573
rect -146 -42657 -112 -42641
rect -146 -43249 -112 -43233
rect 112 -42657 146 -42641
rect 112 -43249 146 -43233
rect -100 -43317 -84 -43283
rect 84 -43317 100 -43283
rect -100 -43425 -84 -43391
rect 84 -43425 100 -43391
rect -146 -43475 -112 -43459
rect -146 -44067 -112 -44051
rect 112 -43475 146 -43459
rect 112 -44067 146 -44051
rect -100 -44135 -84 -44101
rect 84 -44135 100 -44101
rect -100 -44243 -84 -44209
rect 84 -44243 100 -44209
rect -146 -44293 -112 -44277
rect -146 -44885 -112 -44869
rect 112 -44293 146 -44277
rect 112 -44885 146 -44869
rect -100 -44953 -84 -44919
rect 84 -44953 100 -44919
rect -100 -45061 -84 -45027
rect 84 -45061 100 -45027
rect -146 -45111 -112 -45095
rect -146 -45703 -112 -45687
rect 112 -45111 146 -45095
rect 112 -45703 146 -45687
rect -100 -45771 -84 -45737
rect 84 -45771 100 -45737
rect -100 -45879 -84 -45845
rect 84 -45879 100 -45845
rect -146 -45929 -112 -45913
rect -146 -46521 -112 -46505
rect 112 -45929 146 -45913
rect 112 -46521 146 -46505
rect -100 -46589 -84 -46555
rect 84 -46589 100 -46555
rect -100 -46697 -84 -46663
rect 84 -46697 100 -46663
rect -146 -46747 -112 -46731
rect -146 -47339 -112 -47323
rect 112 -46747 146 -46731
rect 112 -47339 146 -47323
rect -100 -47407 -84 -47373
rect 84 -47407 100 -47373
rect -100 -47515 -84 -47481
rect 84 -47515 100 -47481
rect -146 -47565 -112 -47549
rect -146 -48157 -112 -48141
rect 112 -47565 146 -47549
rect 112 -48157 146 -48141
rect -100 -48225 -84 -48191
rect 84 -48225 100 -48191
rect -100 -48333 -84 -48299
rect 84 -48333 100 -48299
rect -146 -48383 -112 -48367
rect -146 -48975 -112 -48959
rect 112 -48383 146 -48367
rect 112 -48975 146 -48959
rect -100 -49043 -84 -49009
rect 84 -49043 100 -49009
rect -100 -49151 -84 -49117
rect 84 -49151 100 -49117
rect -146 -49201 -112 -49185
rect -146 -49793 -112 -49777
rect 112 -49201 146 -49185
rect 112 -49793 146 -49777
rect -100 -49861 -84 -49827
rect 84 -49861 100 -49827
rect -100 -49969 -84 -49935
rect 84 -49969 100 -49935
rect -146 -50019 -112 -50003
rect -146 -50611 -112 -50595
rect 112 -50019 146 -50003
rect 112 -50611 146 -50595
rect -100 -50679 -84 -50645
rect 84 -50679 100 -50645
rect -100 -50787 -84 -50753
rect 84 -50787 100 -50753
rect -146 -50837 -112 -50821
rect -146 -51429 -112 -51413
rect 112 -50837 146 -50821
rect 112 -51429 146 -51413
rect -100 -51497 -84 -51463
rect 84 -51497 100 -51463
rect -100 -51605 -84 -51571
rect 84 -51605 100 -51571
rect -146 -51655 -112 -51639
rect -146 -52247 -112 -52231
rect 112 -51655 146 -51639
rect 112 -52247 146 -52231
rect -100 -52315 -84 -52281
rect 84 -52315 100 -52281
rect -100 -52423 -84 -52389
rect 84 -52423 100 -52389
rect -146 -52473 -112 -52457
rect -146 -53065 -112 -53049
rect 112 -52473 146 -52457
rect 112 -53065 146 -53049
rect -100 -53133 -84 -53099
rect 84 -53133 100 -53099
rect -100 -53241 -84 -53207
rect 84 -53241 100 -53207
rect -146 -53291 -112 -53275
rect -146 -53883 -112 -53867
rect 112 -53291 146 -53275
rect 112 -53883 146 -53867
rect -100 -53951 -84 -53917
rect 84 -53951 100 -53917
rect -100 -54059 -84 -54025
rect 84 -54059 100 -54025
rect -146 -54109 -112 -54093
rect -146 -54701 -112 -54685
rect 112 -54109 146 -54093
rect 112 -54701 146 -54685
rect -100 -54769 -84 -54735
rect 84 -54769 100 -54735
rect -100 -54877 -84 -54843
rect 84 -54877 100 -54843
rect -146 -54927 -112 -54911
rect -146 -55519 -112 -55503
rect 112 -54927 146 -54911
rect 112 -55519 146 -55503
rect -100 -55587 -84 -55553
rect 84 -55587 100 -55553
rect -100 -55695 -84 -55661
rect 84 -55695 100 -55661
rect -146 -55745 -112 -55729
rect -146 -56337 -112 -56321
rect 112 -55745 146 -55729
rect 112 -56337 146 -56321
rect -100 -56405 -84 -56371
rect 84 -56405 100 -56371
rect -100 -56513 -84 -56479
rect 84 -56513 100 -56479
rect -146 -56563 -112 -56547
rect -146 -57155 -112 -57139
rect 112 -56563 146 -56547
rect 112 -57155 146 -57139
rect -100 -57223 -84 -57189
rect 84 -57223 100 -57189
rect -100 -57331 -84 -57297
rect 84 -57331 100 -57297
rect -146 -57381 -112 -57365
rect -146 -57973 -112 -57957
rect 112 -57381 146 -57365
rect 112 -57973 146 -57957
rect -100 -58041 -84 -58007
rect 84 -58041 100 -58007
rect -100 -58149 -84 -58115
rect 84 -58149 100 -58115
rect -146 -58199 -112 -58183
rect -146 -58791 -112 -58775
rect 112 -58199 146 -58183
rect 112 -58791 146 -58775
rect -100 -58859 -84 -58825
rect 84 -58859 100 -58825
rect -100 -58967 -84 -58933
rect 84 -58967 100 -58933
rect -146 -59017 -112 -59001
rect -146 -59609 -112 -59593
rect 112 -59017 146 -59001
rect 112 -59609 146 -59593
rect -100 -59677 -84 -59643
rect 84 -59677 100 -59643
rect -100 -59785 -84 -59751
rect 84 -59785 100 -59751
rect -146 -59835 -112 -59819
rect -146 -60427 -112 -60411
rect 112 -59835 146 -59819
rect 112 -60427 146 -60411
rect -100 -60495 -84 -60461
rect 84 -60495 100 -60461
rect -100 -60603 -84 -60569
rect 84 -60603 100 -60569
rect -146 -60653 -112 -60637
rect -146 -61245 -112 -61229
rect 112 -60653 146 -60637
rect 112 -61245 146 -61229
rect -100 -61313 -84 -61279
rect 84 -61313 100 -61279
rect -100 -61421 -84 -61387
rect 84 -61421 100 -61387
rect -146 -61471 -112 -61455
rect -146 -62063 -112 -62047
rect 112 -61471 146 -61455
rect 112 -62063 146 -62047
rect -100 -62131 -84 -62097
rect 84 -62131 100 -62097
rect -100 -62239 -84 -62205
rect 84 -62239 100 -62205
rect -146 -62289 -112 -62273
rect -146 -62881 -112 -62865
rect 112 -62289 146 -62273
rect 112 -62881 146 -62865
rect -100 -62949 -84 -62915
rect 84 -62949 100 -62915
rect -100 -63057 -84 -63023
rect 84 -63057 100 -63023
rect -146 -63107 -112 -63091
rect -146 -63699 -112 -63683
rect 112 -63107 146 -63091
rect 112 -63699 146 -63683
rect -100 -63767 -84 -63733
rect 84 -63767 100 -63733
rect -100 -63875 -84 -63841
rect 84 -63875 100 -63841
rect -146 -63925 -112 -63909
rect -146 -64517 -112 -64501
rect 112 -63925 146 -63909
rect 112 -64517 146 -64501
rect -100 -64585 -84 -64551
rect 84 -64585 100 -64551
rect -100 -64693 -84 -64659
rect 84 -64693 100 -64659
rect -146 -64743 -112 -64727
rect -146 -65335 -112 -65319
rect 112 -64743 146 -64727
rect 112 -65335 146 -65319
rect -100 -65403 -84 -65369
rect 84 -65403 100 -65369
rect -100 -65511 -84 -65477
rect 84 -65511 100 -65477
rect -146 -65561 -112 -65545
rect -146 -66153 -112 -66137
rect 112 -65561 146 -65545
rect 112 -66153 146 -66137
rect -100 -66221 -84 -66187
rect 84 -66221 100 -66187
rect -100 -66329 -84 -66295
rect 84 -66329 100 -66295
rect -146 -66379 -112 -66363
rect -146 -66971 -112 -66955
rect 112 -66379 146 -66363
rect 112 -66971 146 -66955
rect -100 -67039 -84 -67005
rect 84 -67039 100 -67005
rect -100 -67147 -84 -67113
rect 84 -67147 100 -67113
rect -146 -67197 -112 -67181
rect -146 -67789 -112 -67773
rect 112 -67197 146 -67181
rect 112 -67789 146 -67773
rect -100 -67857 -84 -67823
rect 84 -67857 100 -67823
rect -100 -67965 -84 -67931
rect 84 -67965 100 -67931
rect -146 -68015 -112 -67999
rect -146 -68607 -112 -68591
rect 112 -68015 146 -67999
rect 112 -68607 146 -68591
rect -100 -68675 -84 -68641
rect 84 -68675 100 -68641
rect -100 -68783 -84 -68749
rect 84 -68783 100 -68749
rect -146 -68833 -112 -68817
rect -146 -69425 -112 -69409
rect 112 -68833 146 -68817
rect 112 -69425 146 -69409
rect -100 -69493 -84 -69459
rect 84 -69493 100 -69459
rect -100 -69601 -84 -69567
rect 84 -69601 100 -69567
rect -146 -69651 -112 -69635
rect -146 -70243 -112 -70227
rect 112 -69651 146 -69635
rect 112 -70243 146 -70227
rect -100 -70311 -84 -70277
rect 84 -70311 100 -70277
rect -100 -70419 -84 -70385
rect 84 -70419 100 -70385
rect -146 -70469 -112 -70453
rect -146 -71061 -112 -71045
rect 112 -70469 146 -70453
rect 112 -71061 146 -71045
rect -100 -71129 -84 -71095
rect 84 -71129 100 -71095
rect -100 -71237 -84 -71203
rect 84 -71237 100 -71203
rect -146 -71287 -112 -71271
rect -146 -71879 -112 -71863
rect 112 -71287 146 -71271
rect 112 -71879 146 -71863
rect -100 -71947 -84 -71913
rect 84 -71947 100 -71913
rect -100 -72055 -84 -72021
rect 84 -72055 100 -72021
rect -146 -72105 -112 -72089
rect -146 -72697 -112 -72681
rect 112 -72105 146 -72089
rect 112 -72697 146 -72681
rect -100 -72765 -84 -72731
rect 84 -72765 100 -72731
rect -100 -72873 -84 -72839
rect 84 -72873 100 -72839
rect -146 -72923 -112 -72907
rect -146 -73515 -112 -73499
rect 112 -72923 146 -72907
rect 112 -73515 146 -73499
rect -100 -73583 -84 -73549
rect 84 -73583 100 -73549
rect -100 -73691 -84 -73657
rect 84 -73691 100 -73657
rect -146 -73741 -112 -73725
rect -146 -74333 -112 -74317
rect 112 -73741 146 -73725
rect 112 -74333 146 -74317
rect -100 -74401 -84 -74367
rect 84 -74401 100 -74367
rect -100 -74509 -84 -74475
rect 84 -74509 100 -74475
rect -146 -74559 -112 -74543
rect -146 -75151 -112 -75135
rect 112 -74559 146 -74543
rect 112 -75151 146 -75135
rect -100 -75219 -84 -75185
rect 84 -75219 100 -75185
rect -100 -75327 -84 -75293
rect 84 -75327 100 -75293
rect -146 -75377 -112 -75361
rect -146 -75969 -112 -75953
rect 112 -75377 146 -75361
rect 112 -75969 146 -75953
rect -100 -76037 -84 -76003
rect 84 -76037 100 -76003
rect -100 -76145 -84 -76111
rect 84 -76145 100 -76111
rect -146 -76195 -112 -76179
rect -146 -76787 -112 -76771
rect 112 -76195 146 -76179
rect 112 -76787 146 -76771
rect -100 -76855 -84 -76821
rect 84 -76855 100 -76821
rect -100 -76963 -84 -76929
rect 84 -76963 100 -76929
rect -146 -77013 -112 -76997
rect -146 -77605 -112 -77589
rect 112 -77013 146 -76997
rect 112 -77605 146 -77589
rect -100 -77673 -84 -77639
rect 84 -77673 100 -77639
rect -100 -77781 -84 -77747
rect 84 -77781 100 -77747
rect -146 -77831 -112 -77815
rect -146 -78423 -112 -78407
rect 112 -77831 146 -77815
rect 112 -78423 146 -78407
rect -100 -78491 -84 -78457
rect 84 -78491 100 -78457
rect -100 -78599 -84 -78565
rect 84 -78599 100 -78565
rect -146 -78649 -112 -78633
rect -146 -79241 -112 -79225
rect 112 -78649 146 -78633
rect 112 -79241 146 -79225
rect -100 -79309 -84 -79275
rect 84 -79309 100 -79275
rect -100 -79417 -84 -79383
rect 84 -79417 100 -79383
rect -146 -79467 -112 -79451
rect -146 -80059 -112 -80043
rect 112 -79467 146 -79451
rect 112 -80059 146 -80043
rect -100 -80127 -84 -80093
rect 84 -80127 100 -80093
rect -100 -80235 -84 -80201
rect 84 -80235 100 -80201
rect -146 -80285 -112 -80269
rect -146 -80877 -112 -80861
rect 112 -80285 146 -80269
rect 112 -80877 146 -80861
rect -100 -80945 -84 -80911
rect 84 -80945 100 -80911
rect -100 -81053 -84 -81019
rect 84 -81053 100 -81019
rect -146 -81103 -112 -81087
rect -146 -81695 -112 -81679
rect 112 -81103 146 -81087
rect 112 -81695 146 -81679
rect -100 -81763 -84 -81729
rect 84 -81763 100 -81729
rect -100 -81871 -84 -81837
rect 84 -81871 100 -81837
rect -146 -81921 -112 -81905
rect -146 -82513 -112 -82497
rect 112 -81921 146 -81905
rect 112 -82513 146 -82497
rect -100 -82581 -84 -82547
rect 84 -82581 100 -82547
rect -100 -82689 -84 -82655
rect 84 -82689 100 -82655
rect -146 -82739 -112 -82723
rect -146 -83331 -112 -83315
rect 112 -82739 146 -82723
rect 112 -83331 146 -83315
rect -100 -83399 -84 -83365
rect 84 -83399 100 -83365
rect -100 -83507 -84 -83473
rect 84 -83507 100 -83473
rect -146 -83557 -112 -83541
rect -146 -84149 -112 -84133
rect 112 -83557 146 -83541
rect 112 -84149 146 -84133
rect -100 -84217 -84 -84183
rect 84 -84217 100 -84183
rect -100 -84325 -84 -84291
rect 84 -84325 100 -84291
rect -146 -84375 -112 -84359
rect -146 -84967 -112 -84951
rect 112 -84375 146 -84359
rect 112 -84967 146 -84951
rect -100 -85035 -84 -85001
rect 84 -85035 100 -85001
rect -100 -85143 -84 -85109
rect 84 -85143 100 -85109
rect -146 -85193 -112 -85177
rect -146 -85785 -112 -85769
rect 112 -85193 146 -85177
rect 112 -85785 146 -85769
rect -100 -85853 -84 -85819
rect 84 -85853 100 -85819
rect -100 -85961 -84 -85927
rect 84 -85961 100 -85927
rect -146 -86011 -112 -85995
rect -146 -86603 -112 -86587
rect 112 -86011 146 -85995
rect 112 -86603 146 -86587
rect -100 -86671 -84 -86637
rect 84 -86671 100 -86637
rect -100 -86779 -84 -86745
rect 84 -86779 100 -86745
rect -146 -86829 -112 -86813
rect -146 -87421 -112 -87405
rect 112 -86829 146 -86813
rect 112 -87421 146 -87405
rect -100 -87489 -84 -87455
rect 84 -87489 100 -87455
rect -100 -87597 -84 -87563
rect 84 -87597 100 -87563
rect -146 -87647 -112 -87631
rect -146 -88239 -112 -88223
rect 112 -87647 146 -87631
rect 112 -88239 146 -88223
rect -100 -88307 -84 -88273
rect 84 -88307 100 -88273
rect -100 -88415 -84 -88381
rect 84 -88415 100 -88381
rect -146 -88465 -112 -88449
rect -146 -89057 -112 -89041
rect 112 -88465 146 -88449
rect 112 -89057 146 -89041
rect -100 -89125 -84 -89091
rect 84 -89125 100 -89091
rect -100 -89233 -84 -89199
rect 84 -89233 100 -89199
rect -146 -89283 -112 -89267
rect -146 -89875 -112 -89859
rect 112 -89283 146 -89267
rect 112 -89875 146 -89859
rect -100 -89943 -84 -89909
rect 84 -89943 100 -89909
rect -100 -90051 -84 -90017
rect 84 -90051 100 -90017
rect -146 -90101 -112 -90085
rect -146 -90693 -112 -90677
rect 112 -90101 146 -90085
rect 112 -90693 146 -90677
rect -100 -90761 -84 -90727
rect 84 -90761 100 -90727
rect -100 -90869 -84 -90835
rect 84 -90869 100 -90835
rect -146 -90919 -112 -90903
rect -146 -91511 -112 -91495
rect 112 -90919 146 -90903
rect 112 -91511 146 -91495
rect -100 -91579 -84 -91545
rect 84 -91579 100 -91545
rect -100 -91687 -84 -91653
rect 84 -91687 100 -91653
rect -146 -91737 -112 -91721
rect -146 -92329 -112 -92313
rect 112 -91737 146 -91721
rect 112 -92329 146 -92313
rect -100 -92397 -84 -92363
rect 84 -92397 100 -92363
rect -100 -92505 -84 -92471
rect 84 -92505 100 -92471
rect -146 -92555 -112 -92539
rect -146 -93147 -112 -93131
rect 112 -92555 146 -92539
rect 112 -93147 146 -93131
rect -100 -93215 -84 -93181
rect 84 -93215 100 -93181
rect -100 -93323 -84 -93289
rect 84 -93323 100 -93289
rect -146 -93373 -112 -93357
rect -146 -93965 -112 -93949
rect 112 -93373 146 -93357
rect 112 -93965 146 -93949
rect -100 -94033 -84 -93999
rect 84 -94033 100 -93999
rect -100 -94141 -84 -94107
rect 84 -94141 100 -94107
rect -146 -94191 -112 -94175
rect -146 -94783 -112 -94767
rect 112 -94191 146 -94175
rect 112 -94783 146 -94767
rect -100 -94851 -84 -94817
rect 84 -94851 100 -94817
rect -100 -94959 -84 -94925
rect 84 -94959 100 -94925
rect -146 -95009 -112 -94993
rect -146 -95601 -112 -95585
rect 112 -95009 146 -94993
rect 112 -95601 146 -95585
rect -100 -95669 -84 -95635
rect 84 -95669 100 -95635
rect -100 -95777 -84 -95743
rect 84 -95777 100 -95743
rect -146 -95827 -112 -95811
rect -146 -96419 -112 -96403
rect 112 -95827 146 -95811
rect 112 -96419 146 -96403
rect -100 -96487 -84 -96453
rect 84 -96487 100 -96453
rect -100 -96595 -84 -96561
rect 84 -96595 100 -96561
rect -146 -96645 -112 -96629
rect -146 -97237 -112 -97221
rect 112 -96645 146 -96629
rect 112 -97237 146 -97221
rect -100 -97305 -84 -97271
rect 84 -97305 100 -97271
rect -100 -97413 -84 -97379
rect 84 -97413 100 -97379
rect -146 -97463 -112 -97447
rect -146 -98055 -112 -98039
rect 112 -97463 146 -97447
rect 112 -98055 146 -98039
rect -100 -98123 -84 -98089
rect 84 -98123 100 -98089
rect -100 -98231 -84 -98197
rect 84 -98231 100 -98197
rect -146 -98281 -112 -98265
rect -146 -98873 -112 -98857
rect 112 -98281 146 -98265
rect 112 -98873 146 -98857
rect -100 -98941 -84 -98907
rect 84 -98941 100 -98907
rect -100 -99049 -84 -99015
rect 84 -99049 100 -99015
rect -146 -99099 -112 -99083
rect -146 -99691 -112 -99675
rect 112 -99099 146 -99083
rect 112 -99691 146 -99675
rect -100 -99759 -84 -99725
rect 84 -99759 100 -99725
rect -100 -99867 -84 -99833
rect 84 -99867 100 -99833
rect -146 -99917 -112 -99901
rect -146 -100509 -112 -100493
rect 112 -99917 146 -99901
rect 112 -100509 146 -100493
rect -100 -100577 -84 -100543
rect 84 -100577 100 -100543
rect -100 -100685 -84 -100651
rect 84 -100685 100 -100651
rect -146 -100735 -112 -100719
rect -146 -101327 -112 -101311
rect 112 -100735 146 -100719
rect 112 -101327 146 -101311
rect -100 -101395 -84 -101361
rect 84 -101395 100 -101361
rect -100 -101503 -84 -101469
rect 84 -101503 100 -101469
rect -146 -101553 -112 -101537
rect -146 -102145 -112 -102129
rect 112 -101553 146 -101537
rect 112 -102145 146 -102129
rect -100 -102213 -84 -102179
rect 84 -102213 100 -102179
rect -100 -102321 -84 -102287
rect 84 -102321 100 -102287
rect -146 -102371 -112 -102355
rect -146 -102963 -112 -102947
rect 112 -102371 146 -102355
rect 112 -102963 146 -102947
rect -100 -103031 -84 -102997
rect 84 -103031 100 -102997
rect -100 -103139 -84 -103105
rect 84 -103139 100 -103105
rect -146 -103189 -112 -103173
rect -146 -103781 -112 -103765
rect 112 -103189 146 -103173
rect 112 -103781 146 -103765
rect -100 -103849 -84 -103815
rect 84 -103849 100 -103815
rect -100 -103957 -84 -103923
rect 84 -103957 100 -103923
rect -146 -104007 -112 -103991
rect -146 -104599 -112 -104583
rect 112 -104007 146 -103991
rect 112 -104599 146 -104583
rect -100 -104667 -84 -104633
rect 84 -104667 100 -104633
rect -280 -104771 -246 -104709
rect 246 -104771 280 -104709
rect -280 -104805 -184 -104771
rect 184 -104805 280 -104771
<< viali >>
rect -84 104633 84 104667
rect -146 104007 -112 104583
rect 112 104007 146 104583
rect -84 103923 84 103957
rect -84 103815 84 103849
rect -146 103189 -112 103765
rect 112 103189 146 103765
rect -84 103105 84 103139
rect -84 102997 84 103031
rect -146 102371 -112 102947
rect 112 102371 146 102947
rect -84 102287 84 102321
rect -84 102179 84 102213
rect -146 101553 -112 102129
rect 112 101553 146 102129
rect -84 101469 84 101503
rect -84 101361 84 101395
rect -146 100735 -112 101311
rect 112 100735 146 101311
rect -84 100651 84 100685
rect -84 100543 84 100577
rect -146 99917 -112 100493
rect 112 99917 146 100493
rect -84 99833 84 99867
rect -84 99725 84 99759
rect -146 99099 -112 99675
rect 112 99099 146 99675
rect -84 99015 84 99049
rect -84 98907 84 98941
rect -146 98281 -112 98857
rect 112 98281 146 98857
rect -84 98197 84 98231
rect -84 98089 84 98123
rect -146 97463 -112 98039
rect 112 97463 146 98039
rect -84 97379 84 97413
rect -84 97271 84 97305
rect -146 96645 -112 97221
rect 112 96645 146 97221
rect -84 96561 84 96595
rect -84 96453 84 96487
rect -146 95827 -112 96403
rect 112 95827 146 96403
rect -84 95743 84 95777
rect -84 95635 84 95669
rect -146 95009 -112 95585
rect 112 95009 146 95585
rect -84 94925 84 94959
rect -84 94817 84 94851
rect -146 94191 -112 94767
rect 112 94191 146 94767
rect -84 94107 84 94141
rect -84 93999 84 94033
rect -146 93373 -112 93949
rect 112 93373 146 93949
rect -84 93289 84 93323
rect -84 93181 84 93215
rect -146 92555 -112 93131
rect 112 92555 146 93131
rect -84 92471 84 92505
rect -84 92363 84 92397
rect -146 91737 -112 92313
rect 112 91737 146 92313
rect -84 91653 84 91687
rect -84 91545 84 91579
rect -146 90919 -112 91495
rect 112 90919 146 91495
rect -84 90835 84 90869
rect -84 90727 84 90761
rect -146 90101 -112 90677
rect 112 90101 146 90677
rect -84 90017 84 90051
rect -84 89909 84 89943
rect -146 89283 -112 89859
rect 112 89283 146 89859
rect -84 89199 84 89233
rect -84 89091 84 89125
rect -146 88465 -112 89041
rect 112 88465 146 89041
rect -84 88381 84 88415
rect -84 88273 84 88307
rect -146 87647 -112 88223
rect 112 87647 146 88223
rect -84 87563 84 87597
rect -84 87455 84 87489
rect -146 86829 -112 87405
rect 112 86829 146 87405
rect -84 86745 84 86779
rect -84 86637 84 86671
rect -146 86011 -112 86587
rect 112 86011 146 86587
rect -84 85927 84 85961
rect -84 85819 84 85853
rect -146 85193 -112 85769
rect 112 85193 146 85769
rect -84 85109 84 85143
rect -84 85001 84 85035
rect -146 84375 -112 84951
rect 112 84375 146 84951
rect -84 84291 84 84325
rect -84 84183 84 84217
rect -146 83557 -112 84133
rect 112 83557 146 84133
rect -84 83473 84 83507
rect -84 83365 84 83399
rect -146 82739 -112 83315
rect 112 82739 146 83315
rect -84 82655 84 82689
rect -84 82547 84 82581
rect -146 81921 -112 82497
rect 112 81921 146 82497
rect -84 81837 84 81871
rect -84 81729 84 81763
rect -146 81103 -112 81679
rect 112 81103 146 81679
rect -84 81019 84 81053
rect -84 80911 84 80945
rect -146 80285 -112 80861
rect 112 80285 146 80861
rect -84 80201 84 80235
rect -84 80093 84 80127
rect -146 79467 -112 80043
rect 112 79467 146 80043
rect -84 79383 84 79417
rect -84 79275 84 79309
rect -146 78649 -112 79225
rect 112 78649 146 79225
rect -84 78565 84 78599
rect -84 78457 84 78491
rect -146 77831 -112 78407
rect 112 77831 146 78407
rect -84 77747 84 77781
rect -84 77639 84 77673
rect -146 77013 -112 77589
rect 112 77013 146 77589
rect -84 76929 84 76963
rect -84 76821 84 76855
rect -146 76195 -112 76771
rect 112 76195 146 76771
rect -84 76111 84 76145
rect -84 76003 84 76037
rect -146 75377 -112 75953
rect 112 75377 146 75953
rect -84 75293 84 75327
rect -84 75185 84 75219
rect -146 74559 -112 75135
rect 112 74559 146 75135
rect -84 74475 84 74509
rect -84 74367 84 74401
rect -146 73741 -112 74317
rect 112 73741 146 74317
rect -84 73657 84 73691
rect -84 73549 84 73583
rect -146 72923 -112 73499
rect 112 72923 146 73499
rect -84 72839 84 72873
rect -84 72731 84 72765
rect -146 72105 -112 72681
rect 112 72105 146 72681
rect -84 72021 84 72055
rect -84 71913 84 71947
rect -146 71287 -112 71863
rect 112 71287 146 71863
rect -84 71203 84 71237
rect -84 71095 84 71129
rect -146 70469 -112 71045
rect 112 70469 146 71045
rect -84 70385 84 70419
rect -84 70277 84 70311
rect -146 69651 -112 70227
rect 112 69651 146 70227
rect -84 69567 84 69601
rect -84 69459 84 69493
rect -146 68833 -112 69409
rect 112 68833 146 69409
rect -84 68749 84 68783
rect -84 68641 84 68675
rect -146 68015 -112 68591
rect 112 68015 146 68591
rect -84 67931 84 67965
rect -84 67823 84 67857
rect -146 67197 -112 67773
rect 112 67197 146 67773
rect -84 67113 84 67147
rect -84 67005 84 67039
rect -146 66379 -112 66955
rect 112 66379 146 66955
rect -84 66295 84 66329
rect -84 66187 84 66221
rect -146 65561 -112 66137
rect 112 65561 146 66137
rect -84 65477 84 65511
rect -84 65369 84 65403
rect -146 64743 -112 65319
rect 112 64743 146 65319
rect -84 64659 84 64693
rect -84 64551 84 64585
rect -146 63925 -112 64501
rect 112 63925 146 64501
rect -84 63841 84 63875
rect -84 63733 84 63767
rect -146 63107 -112 63683
rect 112 63107 146 63683
rect -84 63023 84 63057
rect -84 62915 84 62949
rect -146 62289 -112 62865
rect 112 62289 146 62865
rect -84 62205 84 62239
rect -84 62097 84 62131
rect -146 61471 -112 62047
rect 112 61471 146 62047
rect -84 61387 84 61421
rect -84 61279 84 61313
rect -146 60653 -112 61229
rect 112 60653 146 61229
rect -84 60569 84 60603
rect -84 60461 84 60495
rect -146 59835 -112 60411
rect 112 59835 146 60411
rect -84 59751 84 59785
rect -84 59643 84 59677
rect -146 59017 -112 59593
rect 112 59017 146 59593
rect -84 58933 84 58967
rect -84 58825 84 58859
rect -146 58199 -112 58775
rect 112 58199 146 58775
rect -84 58115 84 58149
rect -84 58007 84 58041
rect -146 57381 -112 57957
rect 112 57381 146 57957
rect -84 57297 84 57331
rect -84 57189 84 57223
rect -146 56563 -112 57139
rect 112 56563 146 57139
rect -84 56479 84 56513
rect -84 56371 84 56405
rect -146 55745 -112 56321
rect 112 55745 146 56321
rect -84 55661 84 55695
rect -84 55553 84 55587
rect -146 54927 -112 55503
rect 112 54927 146 55503
rect -84 54843 84 54877
rect -84 54735 84 54769
rect -146 54109 -112 54685
rect 112 54109 146 54685
rect -84 54025 84 54059
rect -84 53917 84 53951
rect -146 53291 -112 53867
rect 112 53291 146 53867
rect -84 53207 84 53241
rect -84 53099 84 53133
rect -146 52473 -112 53049
rect 112 52473 146 53049
rect -84 52389 84 52423
rect -84 52281 84 52315
rect -146 51655 -112 52231
rect 112 51655 146 52231
rect -84 51571 84 51605
rect -84 51463 84 51497
rect -146 50837 -112 51413
rect 112 50837 146 51413
rect -84 50753 84 50787
rect -84 50645 84 50679
rect -146 50019 -112 50595
rect 112 50019 146 50595
rect -84 49935 84 49969
rect -84 49827 84 49861
rect -146 49201 -112 49777
rect 112 49201 146 49777
rect -84 49117 84 49151
rect -84 49009 84 49043
rect -146 48383 -112 48959
rect 112 48383 146 48959
rect -84 48299 84 48333
rect -84 48191 84 48225
rect -146 47565 -112 48141
rect 112 47565 146 48141
rect -84 47481 84 47515
rect -84 47373 84 47407
rect -146 46747 -112 47323
rect 112 46747 146 47323
rect -84 46663 84 46697
rect -84 46555 84 46589
rect -146 45929 -112 46505
rect 112 45929 146 46505
rect -84 45845 84 45879
rect -84 45737 84 45771
rect -146 45111 -112 45687
rect 112 45111 146 45687
rect -84 45027 84 45061
rect -84 44919 84 44953
rect -146 44293 -112 44869
rect 112 44293 146 44869
rect -84 44209 84 44243
rect -84 44101 84 44135
rect -146 43475 -112 44051
rect 112 43475 146 44051
rect -84 43391 84 43425
rect -84 43283 84 43317
rect -146 42657 -112 43233
rect 112 42657 146 43233
rect -84 42573 84 42607
rect -84 42465 84 42499
rect -146 41839 -112 42415
rect 112 41839 146 42415
rect -84 41755 84 41789
rect -84 41647 84 41681
rect -146 41021 -112 41597
rect 112 41021 146 41597
rect -84 40937 84 40971
rect -84 40829 84 40863
rect -146 40203 -112 40779
rect 112 40203 146 40779
rect -84 40119 84 40153
rect -84 40011 84 40045
rect -146 39385 -112 39961
rect 112 39385 146 39961
rect -84 39301 84 39335
rect -84 39193 84 39227
rect -146 38567 -112 39143
rect 112 38567 146 39143
rect -84 38483 84 38517
rect -84 38375 84 38409
rect -146 37749 -112 38325
rect 112 37749 146 38325
rect -84 37665 84 37699
rect -84 37557 84 37591
rect -146 36931 -112 37507
rect 112 36931 146 37507
rect -84 36847 84 36881
rect -84 36739 84 36773
rect -146 36113 -112 36689
rect 112 36113 146 36689
rect -84 36029 84 36063
rect -84 35921 84 35955
rect -146 35295 -112 35871
rect 112 35295 146 35871
rect -84 35211 84 35245
rect -84 35103 84 35137
rect -146 34477 -112 35053
rect 112 34477 146 35053
rect -84 34393 84 34427
rect -84 34285 84 34319
rect -146 33659 -112 34235
rect 112 33659 146 34235
rect -84 33575 84 33609
rect -84 33467 84 33501
rect -146 32841 -112 33417
rect 112 32841 146 33417
rect -84 32757 84 32791
rect -84 32649 84 32683
rect -146 32023 -112 32599
rect 112 32023 146 32599
rect -84 31939 84 31973
rect -84 31831 84 31865
rect -146 31205 -112 31781
rect 112 31205 146 31781
rect -84 31121 84 31155
rect -84 31013 84 31047
rect -146 30387 -112 30963
rect 112 30387 146 30963
rect -84 30303 84 30337
rect -84 30195 84 30229
rect -146 29569 -112 30145
rect 112 29569 146 30145
rect -84 29485 84 29519
rect -84 29377 84 29411
rect -146 28751 -112 29327
rect 112 28751 146 29327
rect -84 28667 84 28701
rect -84 28559 84 28593
rect -146 27933 -112 28509
rect 112 27933 146 28509
rect -84 27849 84 27883
rect -84 27741 84 27775
rect -146 27115 -112 27691
rect 112 27115 146 27691
rect -84 27031 84 27065
rect -84 26923 84 26957
rect -146 26297 -112 26873
rect 112 26297 146 26873
rect -84 26213 84 26247
rect -84 26105 84 26139
rect -146 25479 -112 26055
rect 112 25479 146 26055
rect -84 25395 84 25429
rect -84 25287 84 25321
rect -146 24661 -112 25237
rect 112 24661 146 25237
rect -84 24577 84 24611
rect -84 24469 84 24503
rect -146 23843 -112 24419
rect 112 23843 146 24419
rect -84 23759 84 23793
rect -84 23651 84 23685
rect -146 23025 -112 23601
rect 112 23025 146 23601
rect -84 22941 84 22975
rect -84 22833 84 22867
rect -146 22207 -112 22783
rect 112 22207 146 22783
rect -84 22123 84 22157
rect -84 22015 84 22049
rect -146 21389 -112 21965
rect 112 21389 146 21965
rect -84 21305 84 21339
rect -84 21197 84 21231
rect -146 20571 -112 21147
rect 112 20571 146 21147
rect -84 20487 84 20521
rect -84 20379 84 20413
rect -146 19753 -112 20329
rect 112 19753 146 20329
rect -84 19669 84 19703
rect -84 19561 84 19595
rect -146 18935 -112 19511
rect 112 18935 146 19511
rect -84 18851 84 18885
rect -84 18743 84 18777
rect -146 18117 -112 18693
rect 112 18117 146 18693
rect -84 18033 84 18067
rect -84 17925 84 17959
rect -146 17299 -112 17875
rect 112 17299 146 17875
rect -84 17215 84 17249
rect -84 17107 84 17141
rect -146 16481 -112 17057
rect 112 16481 146 17057
rect -84 16397 84 16431
rect -84 16289 84 16323
rect -146 15663 -112 16239
rect 112 15663 146 16239
rect -84 15579 84 15613
rect -84 15471 84 15505
rect -146 14845 -112 15421
rect 112 14845 146 15421
rect -84 14761 84 14795
rect -84 14653 84 14687
rect -146 14027 -112 14603
rect 112 14027 146 14603
rect -84 13943 84 13977
rect -84 13835 84 13869
rect -146 13209 -112 13785
rect 112 13209 146 13785
rect -84 13125 84 13159
rect -84 13017 84 13051
rect -146 12391 -112 12967
rect 112 12391 146 12967
rect -84 12307 84 12341
rect -84 12199 84 12233
rect -146 11573 -112 12149
rect 112 11573 146 12149
rect -84 11489 84 11523
rect -84 11381 84 11415
rect -146 10755 -112 11331
rect 112 10755 146 11331
rect -84 10671 84 10705
rect -84 10563 84 10597
rect -146 9937 -112 10513
rect 112 9937 146 10513
rect -84 9853 84 9887
rect -84 9745 84 9779
rect -146 9119 -112 9695
rect 112 9119 146 9695
rect -84 9035 84 9069
rect -84 8927 84 8961
rect -146 8301 -112 8877
rect 112 8301 146 8877
rect -84 8217 84 8251
rect -84 8109 84 8143
rect -146 7483 -112 8059
rect 112 7483 146 8059
rect -84 7399 84 7433
rect -84 7291 84 7325
rect -146 6665 -112 7241
rect 112 6665 146 7241
rect -84 6581 84 6615
rect -84 6473 84 6507
rect -146 5847 -112 6423
rect 112 5847 146 6423
rect -84 5763 84 5797
rect -84 5655 84 5689
rect -146 5029 -112 5605
rect 112 5029 146 5605
rect -84 4945 84 4979
rect -84 4837 84 4871
rect -146 4211 -112 4787
rect 112 4211 146 4787
rect -84 4127 84 4161
rect -84 4019 84 4053
rect -146 3393 -112 3969
rect 112 3393 146 3969
rect -84 3309 84 3343
rect -84 3201 84 3235
rect -146 2575 -112 3151
rect 112 2575 146 3151
rect -84 2491 84 2525
rect -84 2383 84 2417
rect -146 1757 -112 2333
rect 112 1757 146 2333
rect -84 1673 84 1707
rect -84 1565 84 1599
rect -146 939 -112 1515
rect 112 939 146 1515
rect -84 855 84 889
rect -84 747 84 781
rect -146 121 -112 697
rect 112 121 146 697
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -697 -112 -121
rect 112 -697 146 -121
rect -84 -781 84 -747
rect -84 -889 84 -855
rect -146 -1515 -112 -939
rect 112 -1515 146 -939
rect -84 -1599 84 -1565
rect -84 -1707 84 -1673
rect -146 -2333 -112 -1757
rect 112 -2333 146 -1757
rect -84 -2417 84 -2383
rect -84 -2525 84 -2491
rect -146 -3151 -112 -2575
rect 112 -3151 146 -2575
rect -84 -3235 84 -3201
rect -84 -3343 84 -3309
rect -146 -3969 -112 -3393
rect 112 -3969 146 -3393
rect -84 -4053 84 -4019
rect -84 -4161 84 -4127
rect -146 -4787 -112 -4211
rect 112 -4787 146 -4211
rect -84 -4871 84 -4837
rect -84 -4979 84 -4945
rect -146 -5605 -112 -5029
rect 112 -5605 146 -5029
rect -84 -5689 84 -5655
rect -84 -5797 84 -5763
rect -146 -6423 -112 -5847
rect 112 -6423 146 -5847
rect -84 -6507 84 -6473
rect -84 -6615 84 -6581
rect -146 -7241 -112 -6665
rect 112 -7241 146 -6665
rect -84 -7325 84 -7291
rect -84 -7433 84 -7399
rect -146 -8059 -112 -7483
rect 112 -8059 146 -7483
rect -84 -8143 84 -8109
rect -84 -8251 84 -8217
rect -146 -8877 -112 -8301
rect 112 -8877 146 -8301
rect -84 -8961 84 -8927
rect -84 -9069 84 -9035
rect -146 -9695 -112 -9119
rect 112 -9695 146 -9119
rect -84 -9779 84 -9745
rect -84 -9887 84 -9853
rect -146 -10513 -112 -9937
rect 112 -10513 146 -9937
rect -84 -10597 84 -10563
rect -84 -10705 84 -10671
rect -146 -11331 -112 -10755
rect 112 -11331 146 -10755
rect -84 -11415 84 -11381
rect -84 -11523 84 -11489
rect -146 -12149 -112 -11573
rect 112 -12149 146 -11573
rect -84 -12233 84 -12199
rect -84 -12341 84 -12307
rect -146 -12967 -112 -12391
rect 112 -12967 146 -12391
rect -84 -13051 84 -13017
rect -84 -13159 84 -13125
rect -146 -13785 -112 -13209
rect 112 -13785 146 -13209
rect -84 -13869 84 -13835
rect -84 -13977 84 -13943
rect -146 -14603 -112 -14027
rect 112 -14603 146 -14027
rect -84 -14687 84 -14653
rect -84 -14795 84 -14761
rect -146 -15421 -112 -14845
rect 112 -15421 146 -14845
rect -84 -15505 84 -15471
rect -84 -15613 84 -15579
rect -146 -16239 -112 -15663
rect 112 -16239 146 -15663
rect -84 -16323 84 -16289
rect -84 -16431 84 -16397
rect -146 -17057 -112 -16481
rect 112 -17057 146 -16481
rect -84 -17141 84 -17107
rect -84 -17249 84 -17215
rect -146 -17875 -112 -17299
rect 112 -17875 146 -17299
rect -84 -17959 84 -17925
rect -84 -18067 84 -18033
rect -146 -18693 -112 -18117
rect 112 -18693 146 -18117
rect -84 -18777 84 -18743
rect -84 -18885 84 -18851
rect -146 -19511 -112 -18935
rect 112 -19511 146 -18935
rect -84 -19595 84 -19561
rect -84 -19703 84 -19669
rect -146 -20329 -112 -19753
rect 112 -20329 146 -19753
rect -84 -20413 84 -20379
rect -84 -20521 84 -20487
rect -146 -21147 -112 -20571
rect 112 -21147 146 -20571
rect -84 -21231 84 -21197
rect -84 -21339 84 -21305
rect -146 -21965 -112 -21389
rect 112 -21965 146 -21389
rect -84 -22049 84 -22015
rect -84 -22157 84 -22123
rect -146 -22783 -112 -22207
rect 112 -22783 146 -22207
rect -84 -22867 84 -22833
rect -84 -22975 84 -22941
rect -146 -23601 -112 -23025
rect 112 -23601 146 -23025
rect -84 -23685 84 -23651
rect -84 -23793 84 -23759
rect -146 -24419 -112 -23843
rect 112 -24419 146 -23843
rect -84 -24503 84 -24469
rect -84 -24611 84 -24577
rect -146 -25237 -112 -24661
rect 112 -25237 146 -24661
rect -84 -25321 84 -25287
rect -84 -25429 84 -25395
rect -146 -26055 -112 -25479
rect 112 -26055 146 -25479
rect -84 -26139 84 -26105
rect -84 -26247 84 -26213
rect -146 -26873 -112 -26297
rect 112 -26873 146 -26297
rect -84 -26957 84 -26923
rect -84 -27065 84 -27031
rect -146 -27691 -112 -27115
rect 112 -27691 146 -27115
rect -84 -27775 84 -27741
rect -84 -27883 84 -27849
rect -146 -28509 -112 -27933
rect 112 -28509 146 -27933
rect -84 -28593 84 -28559
rect -84 -28701 84 -28667
rect -146 -29327 -112 -28751
rect 112 -29327 146 -28751
rect -84 -29411 84 -29377
rect -84 -29519 84 -29485
rect -146 -30145 -112 -29569
rect 112 -30145 146 -29569
rect -84 -30229 84 -30195
rect -84 -30337 84 -30303
rect -146 -30963 -112 -30387
rect 112 -30963 146 -30387
rect -84 -31047 84 -31013
rect -84 -31155 84 -31121
rect -146 -31781 -112 -31205
rect 112 -31781 146 -31205
rect -84 -31865 84 -31831
rect -84 -31973 84 -31939
rect -146 -32599 -112 -32023
rect 112 -32599 146 -32023
rect -84 -32683 84 -32649
rect -84 -32791 84 -32757
rect -146 -33417 -112 -32841
rect 112 -33417 146 -32841
rect -84 -33501 84 -33467
rect -84 -33609 84 -33575
rect -146 -34235 -112 -33659
rect 112 -34235 146 -33659
rect -84 -34319 84 -34285
rect -84 -34427 84 -34393
rect -146 -35053 -112 -34477
rect 112 -35053 146 -34477
rect -84 -35137 84 -35103
rect -84 -35245 84 -35211
rect -146 -35871 -112 -35295
rect 112 -35871 146 -35295
rect -84 -35955 84 -35921
rect -84 -36063 84 -36029
rect -146 -36689 -112 -36113
rect 112 -36689 146 -36113
rect -84 -36773 84 -36739
rect -84 -36881 84 -36847
rect -146 -37507 -112 -36931
rect 112 -37507 146 -36931
rect -84 -37591 84 -37557
rect -84 -37699 84 -37665
rect -146 -38325 -112 -37749
rect 112 -38325 146 -37749
rect -84 -38409 84 -38375
rect -84 -38517 84 -38483
rect -146 -39143 -112 -38567
rect 112 -39143 146 -38567
rect -84 -39227 84 -39193
rect -84 -39335 84 -39301
rect -146 -39961 -112 -39385
rect 112 -39961 146 -39385
rect -84 -40045 84 -40011
rect -84 -40153 84 -40119
rect -146 -40779 -112 -40203
rect 112 -40779 146 -40203
rect -84 -40863 84 -40829
rect -84 -40971 84 -40937
rect -146 -41597 -112 -41021
rect 112 -41597 146 -41021
rect -84 -41681 84 -41647
rect -84 -41789 84 -41755
rect -146 -42415 -112 -41839
rect 112 -42415 146 -41839
rect -84 -42499 84 -42465
rect -84 -42607 84 -42573
rect -146 -43233 -112 -42657
rect 112 -43233 146 -42657
rect -84 -43317 84 -43283
rect -84 -43425 84 -43391
rect -146 -44051 -112 -43475
rect 112 -44051 146 -43475
rect -84 -44135 84 -44101
rect -84 -44243 84 -44209
rect -146 -44869 -112 -44293
rect 112 -44869 146 -44293
rect -84 -44953 84 -44919
rect -84 -45061 84 -45027
rect -146 -45687 -112 -45111
rect 112 -45687 146 -45111
rect -84 -45771 84 -45737
rect -84 -45879 84 -45845
rect -146 -46505 -112 -45929
rect 112 -46505 146 -45929
rect -84 -46589 84 -46555
rect -84 -46697 84 -46663
rect -146 -47323 -112 -46747
rect 112 -47323 146 -46747
rect -84 -47407 84 -47373
rect -84 -47515 84 -47481
rect -146 -48141 -112 -47565
rect 112 -48141 146 -47565
rect -84 -48225 84 -48191
rect -84 -48333 84 -48299
rect -146 -48959 -112 -48383
rect 112 -48959 146 -48383
rect -84 -49043 84 -49009
rect -84 -49151 84 -49117
rect -146 -49777 -112 -49201
rect 112 -49777 146 -49201
rect -84 -49861 84 -49827
rect -84 -49969 84 -49935
rect -146 -50595 -112 -50019
rect 112 -50595 146 -50019
rect -84 -50679 84 -50645
rect -84 -50787 84 -50753
rect -146 -51413 -112 -50837
rect 112 -51413 146 -50837
rect -84 -51497 84 -51463
rect -84 -51605 84 -51571
rect -146 -52231 -112 -51655
rect 112 -52231 146 -51655
rect -84 -52315 84 -52281
rect -84 -52423 84 -52389
rect -146 -53049 -112 -52473
rect 112 -53049 146 -52473
rect -84 -53133 84 -53099
rect -84 -53241 84 -53207
rect -146 -53867 -112 -53291
rect 112 -53867 146 -53291
rect -84 -53951 84 -53917
rect -84 -54059 84 -54025
rect -146 -54685 -112 -54109
rect 112 -54685 146 -54109
rect -84 -54769 84 -54735
rect -84 -54877 84 -54843
rect -146 -55503 -112 -54927
rect 112 -55503 146 -54927
rect -84 -55587 84 -55553
rect -84 -55695 84 -55661
rect -146 -56321 -112 -55745
rect 112 -56321 146 -55745
rect -84 -56405 84 -56371
rect -84 -56513 84 -56479
rect -146 -57139 -112 -56563
rect 112 -57139 146 -56563
rect -84 -57223 84 -57189
rect -84 -57331 84 -57297
rect -146 -57957 -112 -57381
rect 112 -57957 146 -57381
rect -84 -58041 84 -58007
rect -84 -58149 84 -58115
rect -146 -58775 -112 -58199
rect 112 -58775 146 -58199
rect -84 -58859 84 -58825
rect -84 -58967 84 -58933
rect -146 -59593 -112 -59017
rect 112 -59593 146 -59017
rect -84 -59677 84 -59643
rect -84 -59785 84 -59751
rect -146 -60411 -112 -59835
rect 112 -60411 146 -59835
rect -84 -60495 84 -60461
rect -84 -60603 84 -60569
rect -146 -61229 -112 -60653
rect 112 -61229 146 -60653
rect -84 -61313 84 -61279
rect -84 -61421 84 -61387
rect -146 -62047 -112 -61471
rect 112 -62047 146 -61471
rect -84 -62131 84 -62097
rect -84 -62239 84 -62205
rect -146 -62865 -112 -62289
rect 112 -62865 146 -62289
rect -84 -62949 84 -62915
rect -84 -63057 84 -63023
rect -146 -63683 -112 -63107
rect 112 -63683 146 -63107
rect -84 -63767 84 -63733
rect -84 -63875 84 -63841
rect -146 -64501 -112 -63925
rect 112 -64501 146 -63925
rect -84 -64585 84 -64551
rect -84 -64693 84 -64659
rect -146 -65319 -112 -64743
rect 112 -65319 146 -64743
rect -84 -65403 84 -65369
rect -84 -65511 84 -65477
rect -146 -66137 -112 -65561
rect 112 -66137 146 -65561
rect -84 -66221 84 -66187
rect -84 -66329 84 -66295
rect -146 -66955 -112 -66379
rect 112 -66955 146 -66379
rect -84 -67039 84 -67005
rect -84 -67147 84 -67113
rect -146 -67773 -112 -67197
rect 112 -67773 146 -67197
rect -84 -67857 84 -67823
rect -84 -67965 84 -67931
rect -146 -68591 -112 -68015
rect 112 -68591 146 -68015
rect -84 -68675 84 -68641
rect -84 -68783 84 -68749
rect -146 -69409 -112 -68833
rect 112 -69409 146 -68833
rect -84 -69493 84 -69459
rect -84 -69601 84 -69567
rect -146 -70227 -112 -69651
rect 112 -70227 146 -69651
rect -84 -70311 84 -70277
rect -84 -70419 84 -70385
rect -146 -71045 -112 -70469
rect 112 -71045 146 -70469
rect -84 -71129 84 -71095
rect -84 -71237 84 -71203
rect -146 -71863 -112 -71287
rect 112 -71863 146 -71287
rect -84 -71947 84 -71913
rect -84 -72055 84 -72021
rect -146 -72681 -112 -72105
rect 112 -72681 146 -72105
rect -84 -72765 84 -72731
rect -84 -72873 84 -72839
rect -146 -73499 -112 -72923
rect 112 -73499 146 -72923
rect -84 -73583 84 -73549
rect -84 -73691 84 -73657
rect -146 -74317 -112 -73741
rect 112 -74317 146 -73741
rect -84 -74401 84 -74367
rect -84 -74509 84 -74475
rect -146 -75135 -112 -74559
rect 112 -75135 146 -74559
rect -84 -75219 84 -75185
rect -84 -75327 84 -75293
rect -146 -75953 -112 -75377
rect 112 -75953 146 -75377
rect -84 -76037 84 -76003
rect -84 -76145 84 -76111
rect -146 -76771 -112 -76195
rect 112 -76771 146 -76195
rect -84 -76855 84 -76821
rect -84 -76963 84 -76929
rect -146 -77589 -112 -77013
rect 112 -77589 146 -77013
rect -84 -77673 84 -77639
rect -84 -77781 84 -77747
rect -146 -78407 -112 -77831
rect 112 -78407 146 -77831
rect -84 -78491 84 -78457
rect -84 -78599 84 -78565
rect -146 -79225 -112 -78649
rect 112 -79225 146 -78649
rect -84 -79309 84 -79275
rect -84 -79417 84 -79383
rect -146 -80043 -112 -79467
rect 112 -80043 146 -79467
rect -84 -80127 84 -80093
rect -84 -80235 84 -80201
rect -146 -80861 -112 -80285
rect 112 -80861 146 -80285
rect -84 -80945 84 -80911
rect -84 -81053 84 -81019
rect -146 -81679 -112 -81103
rect 112 -81679 146 -81103
rect -84 -81763 84 -81729
rect -84 -81871 84 -81837
rect -146 -82497 -112 -81921
rect 112 -82497 146 -81921
rect -84 -82581 84 -82547
rect -84 -82689 84 -82655
rect -146 -83315 -112 -82739
rect 112 -83315 146 -82739
rect -84 -83399 84 -83365
rect -84 -83507 84 -83473
rect -146 -84133 -112 -83557
rect 112 -84133 146 -83557
rect -84 -84217 84 -84183
rect -84 -84325 84 -84291
rect -146 -84951 -112 -84375
rect 112 -84951 146 -84375
rect -84 -85035 84 -85001
rect -84 -85143 84 -85109
rect -146 -85769 -112 -85193
rect 112 -85769 146 -85193
rect -84 -85853 84 -85819
rect -84 -85961 84 -85927
rect -146 -86587 -112 -86011
rect 112 -86587 146 -86011
rect -84 -86671 84 -86637
rect -84 -86779 84 -86745
rect -146 -87405 -112 -86829
rect 112 -87405 146 -86829
rect -84 -87489 84 -87455
rect -84 -87597 84 -87563
rect -146 -88223 -112 -87647
rect 112 -88223 146 -87647
rect -84 -88307 84 -88273
rect -84 -88415 84 -88381
rect -146 -89041 -112 -88465
rect 112 -89041 146 -88465
rect -84 -89125 84 -89091
rect -84 -89233 84 -89199
rect -146 -89859 -112 -89283
rect 112 -89859 146 -89283
rect -84 -89943 84 -89909
rect -84 -90051 84 -90017
rect -146 -90677 -112 -90101
rect 112 -90677 146 -90101
rect -84 -90761 84 -90727
rect -84 -90869 84 -90835
rect -146 -91495 -112 -90919
rect 112 -91495 146 -90919
rect -84 -91579 84 -91545
rect -84 -91687 84 -91653
rect -146 -92313 -112 -91737
rect 112 -92313 146 -91737
rect -84 -92397 84 -92363
rect -84 -92505 84 -92471
rect -146 -93131 -112 -92555
rect 112 -93131 146 -92555
rect -84 -93215 84 -93181
rect -84 -93323 84 -93289
rect -146 -93949 -112 -93373
rect 112 -93949 146 -93373
rect -84 -94033 84 -93999
rect -84 -94141 84 -94107
rect -146 -94767 -112 -94191
rect 112 -94767 146 -94191
rect -84 -94851 84 -94817
rect -84 -94959 84 -94925
rect -146 -95585 -112 -95009
rect 112 -95585 146 -95009
rect -84 -95669 84 -95635
rect -84 -95777 84 -95743
rect -146 -96403 -112 -95827
rect 112 -96403 146 -95827
rect -84 -96487 84 -96453
rect -84 -96595 84 -96561
rect -146 -97221 -112 -96645
rect 112 -97221 146 -96645
rect -84 -97305 84 -97271
rect -84 -97413 84 -97379
rect -146 -98039 -112 -97463
rect 112 -98039 146 -97463
rect -84 -98123 84 -98089
rect -84 -98231 84 -98197
rect -146 -98857 -112 -98281
rect 112 -98857 146 -98281
rect -84 -98941 84 -98907
rect -84 -99049 84 -99015
rect -146 -99675 -112 -99099
rect 112 -99675 146 -99099
rect -84 -99759 84 -99725
rect -84 -99867 84 -99833
rect -146 -100493 -112 -99917
rect 112 -100493 146 -99917
rect -84 -100577 84 -100543
rect -84 -100685 84 -100651
rect -146 -101311 -112 -100735
rect 112 -101311 146 -100735
rect -84 -101395 84 -101361
rect -84 -101503 84 -101469
rect -146 -102129 -112 -101553
rect 112 -102129 146 -101553
rect -84 -102213 84 -102179
rect -84 -102321 84 -102287
rect -146 -102947 -112 -102371
rect 112 -102947 146 -102371
rect -84 -103031 84 -102997
rect -84 -103139 84 -103105
rect -146 -103765 -112 -103189
rect 112 -103765 146 -103189
rect -84 -103849 84 -103815
rect -84 -103957 84 -103923
rect -146 -104583 -112 -104007
rect 112 -104583 146 -104007
rect -84 -104667 84 -104633
<< metal1 >>
rect -96 104667 96 104673
rect -96 104633 -84 104667
rect 84 104633 96 104667
rect -96 104627 96 104633
rect -152 104583 -106 104595
rect -152 104007 -146 104583
rect -112 104007 -106 104583
rect -152 103995 -106 104007
rect 106 104583 152 104595
rect 106 104007 112 104583
rect 146 104007 152 104583
rect 106 103995 152 104007
rect -96 103957 96 103963
rect -96 103923 -84 103957
rect 84 103923 96 103957
rect -96 103917 96 103923
rect -96 103849 96 103855
rect -96 103815 -84 103849
rect 84 103815 96 103849
rect -96 103809 96 103815
rect -152 103765 -106 103777
rect -152 103189 -146 103765
rect -112 103189 -106 103765
rect -152 103177 -106 103189
rect 106 103765 152 103777
rect 106 103189 112 103765
rect 146 103189 152 103765
rect 106 103177 152 103189
rect -96 103139 96 103145
rect -96 103105 -84 103139
rect 84 103105 96 103139
rect -96 103099 96 103105
rect -96 103031 96 103037
rect -96 102997 -84 103031
rect 84 102997 96 103031
rect -96 102991 96 102997
rect -152 102947 -106 102959
rect -152 102371 -146 102947
rect -112 102371 -106 102947
rect -152 102359 -106 102371
rect 106 102947 152 102959
rect 106 102371 112 102947
rect 146 102371 152 102947
rect 106 102359 152 102371
rect -96 102321 96 102327
rect -96 102287 -84 102321
rect 84 102287 96 102321
rect -96 102281 96 102287
rect -96 102213 96 102219
rect -96 102179 -84 102213
rect 84 102179 96 102213
rect -96 102173 96 102179
rect -152 102129 -106 102141
rect -152 101553 -146 102129
rect -112 101553 -106 102129
rect -152 101541 -106 101553
rect 106 102129 152 102141
rect 106 101553 112 102129
rect 146 101553 152 102129
rect 106 101541 152 101553
rect -96 101503 96 101509
rect -96 101469 -84 101503
rect 84 101469 96 101503
rect -96 101463 96 101469
rect -96 101395 96 101401
rect -96 101361 -84 101395
rect 84 101361 96 101395
rect -96 101355 96 101361
rect -152 101311 -106 101323
rect -152 100735 -146 101311
rect -112 100735 -106 101311
rect -152 100723 -106 100735
rect 106 101311 152 101323
rect 106 100735 112 101311
rect 146 100735 152 101311
rect 106 100723 152 100735
rect -96 100685 96 100691
rect -96 100651 -84 100685
rect 84 100651 96 100685
rect -96 100645 96 100651
rect -96 100577 96 100583
rect -96 100543 -84 100577
rect 84 100543 96 100577
rect -96 100537 96 100543
rect -152 100493 -106 100505
rect -152 99917 -146 100493
rect -112 99917 -106 100493
rect -152 99905 -106 99917
rect 106 100493 152 100505
rect 106 99917 112 100493
rect 146 99917 152 100493
rect 106 99905 152 99917
rect -96 99867 96 99873
rect -96 99833 -84 99867
rect 84 99833 96 99867
rect -96 99827 96 99833
rect -96 99759 96 99765
rect -96 99725 -84 99759
rect 84 99725 96 99759
rect -96 99719 96 99725
rect -152 99675 -106 99687
rect -152 99099 -146 99675
rect -112 99099 -106 99675
rect -152 99087 -106 99099
rect 106 99675 152 99687
rect 106 99099 112 99675
rect 146 99099 152 99675
rect 106 99087 152 99099
rect -96 99049 96 99055
rect -96 99015 -84 99049
rect 84 99015 96 99049
rect -96 99009 96 99015
rect -96 98941 96 98947
rect -96 98907 -84 98941
rect 84 98907 96 98941
rect -96 98901 96 98907
rect -152 98857 -106 98869
rect -152 98281 -146 98857
rect -112 98281 -106 98857
rect -152 98269 -106 98281
rect 106 98857 152 98869
rect 106 98281 112 98857
rect 146 98281 152 98857
rect 106 98269 152 98281
rect -96 98231 96 98237
rect -96 98197 -84 98231
rect 84 98197 96 98231
rect -96 98191 96 98197
rect -96 98123 96 98129
rect -96 98089 -84 98123
rect 84 98089 96 98123
rect -96 98083 96 98089
rect -152 98039 -106 98051
rect -152 97463 -146 98039
rect -112 97463 -106 98039
rect -152 97451 -106 97463
rect 106 98039 152 98051
rect 106 97463 112 98039
rect 146 97463 152 98039
rect 106 97451 152 97463
rect -96 97413 96 97419
rect -96 97379 -84 97413
rect 84 97379 96 97413
rect -96 97373 96 97379
rect -96 97305 96 97311
rect -96 97271 -84 97305
rect 84 97271 96 97305
rect -96 97265 96 97271
rect -152 97221 -106 97233
rect -152 96645 -146 97221
rect -112 96645 -106 97221
rect -152 96633 -106 96645
rect 106 97221 152 97233
rect 106 96645 112 97221
rect 146 96645 152 97221
rect 106 96633 152 96645
rect -96 96595 96 96601
rect -96 96561 -84 96595
rect 84 96561 96 96595
rect -96 96555 96 96561
rect -96 96487 96 96493
rect -96 96453 -84 96487
rect 84 96453 96 96487
rect -96 96447 96 96453
rect -152 96403 -106 96415
rect -152 95827 -146 96403
rect -112 95827 -106 96403
rect -152 95815 -106 95827
rect 106 96403 152 96415
rect 106 95827 112 96403
rect 146 95827 152 96403
rect 106 95815 152 95827
rect -96 95777 96 95783
rect -96 95743 -84 95777
rect 84 95743 96 95777
rect -96 95737 96 95743
rect -96 95669 96 95675
rect -96 95635 -84 95669
rect 84 95635 96 95669
rect -96 95629 96 95635
rect -152 95585 -106 95597
rect -152 95009 -146 95585
rect -112 95009 -106 95585
rect -152 94997 -106 95009
rect 106 95585 152 95597
rect 106 95009 112 95585
rect 146 95009 152 95585
rect 106 94997 152 95009
rect -96 94959 96 94965
rect -96 94925 -84 94959
rect 84 94925 96 94959
rect -96 94919 96 94925
rect -96 94851 96 94857
rect -96 94817 -84 94851
rect 84 94817 96 94851
rect -96 94811 96 94817
rect -152 94767 -106 94779
rect -152 94191 -146 94767
rect -112 94191 -106 94767
rect -152 94179 -106 94191
rect 106 94767 152 94779
rect 106 94191 112 94767
rect 146 94191 152 94767
rect 106 94179 152 94191
rect -96 94141 96 94147
rect -96 94107 -84 94141
rect 84 94107 96 94141
rect -96 94101 96 94107
rect -96 94033 96 94039
rect -96 93999 -84 94033
rect 84 93999 96 94033
rect -96 93993 96 93999
rect -152 93949 -106 93961
rect -152 93373 -146 93949
rect -112 93373 -106 93949
rect -152 93361 -106 93373
rect 106 93949 152 93961
rect 106 93373 112 93949
rect 146 93373 152 93949
rect 106 93361 152 93373
rect -96 93323 96 93329
rect -96 93289 -84 93323
rect 84 93289 96 93323
rect -96 93283 96 93289
rect -96 93215 96 93221
rect -96 93181 -84 93215
rect 84 93181 96 93215
rect -96 93175 96 93181
rect -152 93131 -106 93143
rect -152 92555 -146 93131
rect -112 92555 -106 93131
rect -152 92543 -106 92555
rect 106 93131 152 93143
rect 106 92555 112 93131
rect 146 92555 152 93131
rect 106 92543 152 92555
rect -96 92505 96 92511
rect -96 92471 -84 92505
rect 84 92471 96 92505
rect -96 92465 96 92471
rect -96 92397 96 92403
rect -96 92363 -84 92397
rect 84 92363 96 92397
rect -96 92357 96 92363
rect -152 92313 -106 92325
rect -152 91737 -146 92313
rect -112 91737 -106 92313
rect -152 91725 -106 91737
rect 106 92313 152 92325
rect 106 91737 112 92313
rect 146 91737 152 92313
rect 106 91725 152 91737
rect -96 91687 96 91693
rect -96 91653 -84 91687
rect 84 91653 96 91687
rect -96 91647 96 91653
rect -96 91579 96 91585
rect -96 91545 -84 91579
rect 84 91545 96 91579
rect -96 91539 96 91545
rect -152 91495 -106 91507
rect -152 90919 -146 91495
rect -112 90919 -106 91495
rect -152 90907 -106 90919
rect 106 91495 152 91507
rect 106 90919 112 91495
rect 146 90919 152 91495
rect 106 90907 152 90919
rect -96 90869 96 90875
rect -96 90835 -84 90869
rect 84 90835 96 90869
rect -96 90829 96 90835
rect -96 90761 96 90767
rect -96 90727 -84 90761
rect 84 90727 96 90761
rect -96 90721 96 90727
rect -152 90677 -106 90689
rect -152 90101 -146 90677
rect -112 90101 -106 90677
rect -152 90089 -106 90101
rect 106 90677 152 90689
rect 106 90101 112 90677
rect 146 90101 152 90677
rect 106 90089 152 90101
rect -96 90051 96 90057
rect -96 90017 -84 90051
rect 84 90017 96 90051
rect -96 90011 96 90017
rect -96 89943 96 89949
rect -96 89909 -84 89943
rect 84 89909 96 89943
rect -96 89903 96 89909
rect -152 89859 -106 89871
rect -152 89283 -146 89859
rect -112 89283 -106 89859
rect -152 89271 -106 89283
rect 106 89859 152 89871
rect 106 89283 112 89859
rect 146 89283 152 89859
rect 106 89271 152 89283
rect -96 89233 96 89239
rect -96 89199 -84 89233
rect 84 89199 96 89233
rect -96 89193 96 89199
rect -96 89125 96 89131
rect -96 89091 -84 89125
rect 84 89091 96 89125
rect -96 89085 96 89091
rect -152 89041 -106 89053
rect -152 88465 -146 89041
rect -112 88465 -106 89041
rect -152 88453 -106 88465
rect 106 89041 152 89053
rect 106 88465 112 89041
rect 146 88465 152 89041
rect 106 88453 152 88465
rect -96 88415 96 88421
rect -96 88381 -84 88415
rect 84 88381 96 88415
rect -96 88375 96 88381
rect -96 88307 96 88313
rect -96 88273 -84 88307
rect 84 88273 96 88307
rect -96 88267 96 88273
rect -152 88223 -106 88235
rect -152 87647 -146 88223
rect -112 87647 -106 88223
rect -152 87635 -106 87647
rect 106 88223 152 88235
rect 106 87647 112 88223
rect 146 87647 152 88223
rect 106 87635 152 87647
rect -96 87597 96 87603
rect -96 87563 -84 87597
rect 84 87563 96 87597
rect -96 87557 96 87563
rect -96 87489 96 87495
rect -96 87455 -84 87489
rect 84 87455 96 87489
rect -96 87449 96 87455
rect -152 87405 -106 87417
rect -152 86829 -146 87405
rect -112 86829 -106 87405
rect -152 86817 -106 86829
rect 106 87405 152 87417
rect 106 86829 112 87405
rect 146 86829 152 87405
rect 106 86817 152 86829
rect -96 86779 96 86785
rect -96 86745 -84 86779
rect 84 86745 96 86779
rect -96 86739 96 86745
rect -96 86671 96 86677
rect -96 86637 -84 86671
rect 84 86637 96 86671
rect -96 86631 96 86637
rect -152 86587 -106 86599
rect -152 86011 -146 86587
rect -112 86011 -106 86587
rect -152 85999 -106 86011
rect 106 86587 152 86599
rect 106 86011 112 86587
rect 146 86011 152 86587
rect 106 85999 152 86011
rect -96 85961 96 85967
rect -96 85927 -84 85961
rect 84 85927 96 85961
rect -96 85921 96 85927
rect -96 85853 96 85859
rect -96 85819 -84 85853
rect 84 85819 96 85853
rect -96 85813 96 85819
rect -152 85769 -106 85781
rect -152 85193 -146 85769
rect -112 85193 -106 85769
rect -152 85181 -106 85193
rect 106 85769 152 85781
rect 106 85193 112 85769
rect 146 85193 152 85769
rect 106 85181 152 85193
rect -96 85143 96 85149
rect -96 85109 -84 85143
rect 84 85109 96 85143
rect -96 85103 96 85109
rect -96 85035 96 85041
rect -96 85001 -84 85035
rect 84 85001 96 85035
rect -96 84995 96 85001
rect -152 84951 -106 84963
rect -152 84375 -146 84951
rect -112 84375 -106 84951
rect -152 84363 -106 84375
rect 106 84951 152 84963
rect 106 84375 112 84951
rect 146 84375 152 84951
rect 106 84363 152 84375
rect -96 84325 96 84331
rect -96 84291 -84 84325
rect 84 84291 96 84325
rect -96 84285 96 84291
rect -96 84217 96 84223
rect -96 84183 -84 84217
rect 84 84183 96 84217
rect -96 84177 96 84183
rect -152 84133 -106 84145
rect -152 83557 -146 84133
rect -112 83557 -106 84133
rect -152 83545 -106 83557
rect 106 84133 152 84145
rect 106 83557 112 84133
rect 146 83557 152 84133
rect 106 83545 152 83557
rect -96 83507 96 83513
rect -96 83473 -84 83507
rect 84 83473 96 83507
rect -96 83467 96 83473
rect -96 83399 96 83405
rect -96 83365 -84 83399
rect 84 83365 96 83399
rect -96 83359 96 83365
rect -152 83315 -106 83327
rect -152 82739 -146 83315
rect -112 82739 -106 83315
rect -152 82727 -106 82739
rect 106 83315 152 83327
rect 106 82739 112 83315
rect 146 82739 152 83315
rect 106 82727 152 82739
rect -96 82689 96 82695
rect -96 82655 -84 82689
rect 84 82655 96 82689
rect -96 82649 96 82655
rect -96 82581 96 82587
rect -96 82547 -84 82581
rect 84 82547 96 82581
rect -96 82541 96 82547
rect -152 82497 -106 82509
rect -152 81921 -146 82497
rect -112 81921 -106 82497
rect -152 81909 -106 81921
rect 106 82497 152 82509
rect 106 81921 112 82497
rect 146 81921 152 82497
rect 106 81909 152 81921
rect -96 81871 96 81877
rect -96 81837 -84 81871
rect 84 81837 96 81871
rect -96 81831 96 81837
rect -96 81763 96 81769
rect -96 81729 -84 81763
rect 84 81729 96 81763
rect -96 81723 96 81729
rect -152 81679 -106 81691
rect -152 81103 -146 81679
rect -112 81103 -106 81679
rect -152 81091 -106 81103
rect 106 81679 152 81691
rect 106 81103 112 81679
rect 146 81103 152 81679
rect 106 81091 152 81103
rect -96 81053 96 81059
rect -96 81019 -84 81053
rect 84 81019 96 81053
rect -96 81013 96 81019
rect -96 80945 96 80951
rect -96 80911 -84 80945
rect 84 80911 96 80945
rect -96 80905 96 80911
rect -152 80861 -106 80873
rect -152 80285 -146 80861
rect -112 80285 -106 80861
rect -152 80273 -106 80285
rect 106 80861 152 80873
rect 106 80285 112 80861
rect 146 80285 152 80861
rect 106 80273 152 80285
rect -96 80235 96 80241
rect -96 80201 -84 80235
rect 84 80201 96 80235
rect -96 80195 96 80201
rect -96 80127 96 80133
rect -96 80093 -84 80127
rect 84 80093 96 80127
rect -96 80087 96 80093
rect -152 80043 -106 80055
rect -152 79467 -146 80043
rect -112 79467 -106 80043
rect -152 79455 -106 79467
rect 106 80043 152 80055
rect 106 79467 112 80043
rect 146 79467 152 80043
rect 106 79455 152 79467
rect -96 79417 96 79423
rect -96 79383 -84 79417
rect 84 79383 96 79417
rect -96 79377 96 79383
rect -96 79309 96 79315
rect -96 79275 -84 79309
rect 84 79275 96 79309
rect -96 79269 96 79275
rect -152 79225 -106 79237
rect -152 78649 -146 79225
rect -112 78649 -106 79225
rect -152 78637 -106 78649
rect 106 79225 152 79237
rect 106 78649 112 79225
rect 146 78649 152 79225
rect 106 78637 152 78649
rect -96 78599 96 78605
rect -96 78565 -84 78599
rect 84 78565 96 78599
rect -96 78559 96 78565
rect -96 78491 96 78497
rect -96 78457 -84 78491
rect 84 78457 96 78491
rect -96 78451 96 78457
rect -152 78407 -106 78419
rect -152 77831 -146 78407
rect -112 77831 -106 78407
rect -152 77819 -106 77831
rect 106 78407 152 78419
rect 106 77831 112 78407
rect 146 77831 152 78407
rect 106 77819 152 77831
rect -96 77781 96 77787
rect -96 77747 -84 77781
rect 84 77747 96 77781
rect -96 77741 96 77747
rect -96 77673 96 77679
rect -96 77639 -84 77673
rect 84 77639 96 77673
rect -96 77633 96 77639
rect -152 77589 -106 77601
rect -152 77013 -146 77589
rect -112 77013 -106 77589
rect -152 77001 -106 77013
rect 106 77589 152 77601
rect 106 77013 112 77589
rect 146 77013 152 77589
rect 106 77001 152 77013
rect -96 76963 96 76969
rect -96 76929 -84 76963
rect 84 76929 96 76963
rect -96 76923 96 76929
rect -96 76855 96 76861
rect -96 76821 -84 76855
rect 84 76821 96 76855
rect -96 76815 96 76821
rect -152 76771 -106 76783
rect -152 76195 -146 76771
rect -112 76195 -106 76771
rect -152 76183 -106 76195
rect 106 76771 152 76783
rect 106 76195 112 76771
rect 146 76195 152 76771
rect 106 76183 152 76195
rect -96 76145 96 76151
rect -96 76111 -84 76145
rect 84 76111 96 76145
rect -96 76105 96 76111
rect -96 76037 96 76043
rect -96 76003 -84 76037
rect 84 76003 96 76037
rect -96 75997 96 76003
rect -152 75953 -106 75965
rect -152 75377 -146 75953
rect -112 75377 -106 75953
rect -152 75365 -106 75377
rect 106 75953 152 75965
rect 106 75377 112 75953
rect 146 75377 152 75953
rect 106 75365 152 75377
rect -96 75327 96 75333
rect -96 75293 -84 75327
rect 84 75293 96 75327
rect -96 75287 96 75293
rect -96 75219 96 75225
rect -96 75185 -84 75219
rect 84 75185 96 75219
rect -96 75179 96 75185
rect -152 75135 -106 75147
rect -152 74559 -146 75135
rect -112 74559 -106 75135
rect -152 74547 -106 74559
rect 106 75135 152 75147
rect 106 74559 112 75135
rect 146 74559 152 75135
rect 106 74547 152 74559
rect -96 74509 96 74515
rect -96 74475 -84 74509
rect 84 74475 96 74509
rect -96 74469 96 74475
rect -96 74401 96 74407
rect -96 74367 -84 74401
rect 84 74367 96 74401
rect -96 74361 96 74367
rect -152 74317 -106 74329
rect -152 73741 -146 74317
rect -112 73741 -106 74317
rect -152 73729 -106 73741
rect 106 74317 152 74329
rect 106 73741 112 74317
rect 146 73741 152 74317
rect 106 73729 152 73741
rect -96 73691 96 73697
rect -96 73657 -84 73691
rect 84 73657 96 73691
rect -96 73651 96 73657
rect -96 73583 96 73589
rect -96 73549 -84 73583
rect 84 73549 96 73583
rect -96 73543 96 73549
rect -152 73499 -106 73511
rect -152 72923 -146 73499
rect -112 72923 -106 73499
rect -152 72911 -106 72923
rect 106 73499 152 73511
rect 106 72923 112 73499
rect 146 72923 152 73499
rect 106 72911 152 72923
rect -96 72873 96 72879
rect -96 72839 -84 72873
rect 84 72839 96 72873
rect -96 72833 96 72839
rect -96 72765 96 72771
rect -96 72731 -84 72765
rect 84 72731 96 72765
rect -96 72725 96 72731
rect -152 72681 -106 72693
rect -152 72105 -146 72681
rect -112 72105 -106 72681
rect -152 72093 -106 72105
rect 106 72681 152 72693
rect 106 72105 112 72681
rect 146 72105 152 72681
rect 106 72093 152 72105
rect -96 72055 96 72061
rect -96 72021 -84 72055
rect 84 72021 96 72055
rect -96 72015 96 72021
rect -96 71947 96 71953
rect -96 71913 -84 71947
rect 84 71913 96 71947
rect -96 71907 96 71913
rect -152 71863 -106 71875
rect -152 71287 -146 71863
rect -112 71287 -106 71863
rect -152 71275 -106 71287
rect 106 71863 152 71875
rect 106 71287 112 71863
rect 146 71287 152 71863
rect 106 71275 152 71287
rect -96 71237 96 71243
rect -96 71203 -84 71237
rect 84 71203 96 71237
rect -96 71197 96 71203
rect -96 71129 96 71135
rect -96 71095 -84 71129
rect 84 71095 96 71129
rect -96 71089 96 71095
rect -152 71045 -106 71057
rect -152 70469 -146 71045
rect -112 70469 -106 71045
rect -152 70457 -106 70469
rect 106 71045 152 71057
rect 106 70469 112 71045
rect 146 70469 152 71045
rect 106 70457 152 70469
rect -96 70419 96 70425
rect -96 70385 -84 70419
rect 84 70385 96 70419
rect -96 70379 96 70385
rect -96 70311 96 70317
rect -96 70277 -84 70311
rect 84 70277 96 70311
rect -96 70271 96 70277
rect -152 70227 -106 70239
rect -152 69651 -146 70227
rect -112 69651 -106 70227
rect -152 69639 -106 69651
rect 106 70227 152 70239
rect 106 69651 112 70227
rect 146 69651 152 70227
rect 106 69639 152 69651
rect -96 69601 96 69607
rect -96 69567 -84 69601
rect 84 69567 96 69601
rect -96 69561 96 69567
rect -96 69493 96 69499
rect -96 69459 -84 69493
rect 84 69459 96 69493
rect -96 69453 96 69459
rect -152 69409 -106 69421
rect -152 68833 -146 69409
rect -112 68833 -106 69409
rect -152 68821 -106 68833
rect 106 69409 152 69421
rect 106 68833 112 69409
rect 146 68833 152 69409
rect 106 68821 152 68833
rect -96 68783 96 68789
rect -96 68749 -84 68783
rect 84 68749 96 68783
rect -96 68743 96 68749
rect -96 68675 96 68681
rect -96 68641 -84 68675
rect 84 68641 96 68675
rect -96 68635 96 68641
rect -152 68591 -106 68603
rect -152 68015 -146 68591
rect -112 68015 -106 68591
rect -152 68003 -106 68015
rect 106 68591 152 68603
rect 106 68015 112 68591
rect 146 68015 152 68591
rect 106 68003 152 68015
rect -96 67965 96 67971
rect -96 67931 -84 67965
rect 84 67931 96 67965
rect -96 67925 96 67931
rect -96 67857 96 67863
rect -96 67823 -84 67857
rect 84 67823 96 67857
rect -96 67817 96 67823
rect -152 67773 -106 67785
rect -152 67197 -146 67773
rect -112 67197 -106 67773
rect -152 67185 -106 67197
rect 106 67773 152 67785
rect 106 67197 112 67773
rect 146 67197 152 67773
rect 106 67185 152 67197
rect -96 67147 96 67153
rect -96 67113 -84 67147
rect 84 67113 96 67147
rect -96 67107 96 67113
rect -96 67039 96 67045
rect -96 67005 -84 67039
rect 84 67005 96 67039
rect -96 66999 96 67005
rect -152 66955 -106 66967
rect -152 66379 -146 66955
rect -112 66379 -106 66955
rect -152 66367 -106 66379
rect 106 66955 152 66967
rect 106 66379 112 66955
rect 146 66379 152 66955
rect 106 66367 152 66379
rect -96 66329 96 66335
rect -96 66295 -84 66329
rect 84 66295 96 66329
rect -96 66289 96 66295
rect -96 66221 96 66227
rect -96 66187 -84 66221
rect 84 66187 96 66221
rect -96 66181 96 66187
rect -152 66137 -106 66149
rect -152 65561 -146 66137
rect -112 65561 -106 66137
rect -152 65549 -106 65561
rect 106 66137 152 66149
rect 106 65561 112 66137
rect 146 65561 152 66137
rect 106 65549 152 65561
rect -96 65511 96 65517
rect -96 65477 -84 65511
rect 84 65477 96 65511
rect -96 65471 96 65477
rect -96 65403 96 65409
rect -96 65369 -84 65403
rect 84 65369 96 65403
rect -96 65363 96 65369
rect -152 65319 -106 65331
rect -152 64743 -146 65319
rect -112 64743 -106 65319
rect -152 64731 -106 64743
rect 106 65319 152 65331
rect 106 64743 112 65319
rect 146 64743 152 65319
rect 106 64731 152 64743
rect -96 64693 96 64699
rect -96 64659 -84 64693
rect 84 64659 96 64693
rect -96 64653 96 64659
rect -96 64585 96 64591
rect -96 64551 -84 64585
rect 84 64551 96 64585
rect -96 64545 96 64551
rect -152 64501 -106 64513
rect -152 63925 -146 64501
rect -112 63925 -106 64501
rect -152 63913 -106 63925
rect 106 64501 152 64513
rect 106 63925 112 64501
rect 146 63925 152 64501
rect 106 63913 152 63925
rect -96 63875 96 63881
rect -96 63841 -84 63875
rect 84 63841 96 63875
rect -96 63835 96 63841
rect -96 63767 96 63773
rect -96 63733 -84 63767
rect 84 63733 96 63767
rect -96 63727 96 63733
rect -152 63683 -106 63695
rect -152 63107 -146 63683
rect -112 63107 -106 63683
rect -152 63095 -106 63107
rect 106 63683 152 63695
rect 106 63107 112 63683
rect 146 63107 152 63683
rect 106 63095 152 63107
rect -96 63057 96 63063
rect -96 63023 -84 63057
rect 84 63023 96 63057
rect -96 63017 96 63023
rect -96 62949 96 62955
rect -96 62915 -84 62949
rect 84 62915 96 62949
rect -96 62909 96 62915
rect -152 62865 -106 62877
rect -152 62289 -146 62865
rect -112 62289 -106 62865
rect -152 62277 -106 62289
rect 106 62865 152 62877
rect 106 62289 112 62865
rect 146 62289 152 62865
rect 106 62277 152 62289
rect -96 62239 96 62245
rect -96 62205 -84 62239
rect 84 62205 96 62239
rect -96 62199 96 62205
rect -96 62131 96 62137
rect -96 62097 -84 62131
rect 84 62097 96 62131
rect -96 62091 96 62097
rect -152 62047 -106 62059
rect -152 61471 -146 62047
rect -112 61471 -106 62047
rect -152 61459 -106 61471
rect 106 62047 152 62059
rect 106 61471 112 62047
rect 146 61471 152 62047
rect 106 61459 152 61471
rect -96 61421 96 61427
rect -96 61387 -84 61421
rect 84 61387 96 61421
rect -96 61381 96 61387
rect -96 61313 96 61319
rect -96 61279 -84 61313
rect 84 61279 96 61313
rect -96 61273 96 61279
rect -152 61229 -106 61241
rect -152 60653 -146 61229
rect -112 60653 -106 61229
rect -152 60641 -106 60653
rect 106 61229 152 61241
rect 106 60653 112 61229
rect 146 60653 152 61229
rect 106 60641 152 60653
rect -96 60603 96 60609
rect -96 60569 -84 60603
rect 84 60569 96 60603
rect -96 60563 96 60569
rect -96 60495 96 60501
rect -96 60461 -84 60495
rect 84 60461 96 60495
rect -96 60455 96 60461
rect -152 60411 -106 60423
rect -152 59835 -146 60411
rect -112 59835 -106 60411
rect -152 59823 -106 59835
rect 106 60411 152 60423
rect 106 59835 112 60411
rect 146 59835 152 60411
rect 106 59823 152 59835
rect -96 59785 96 59791
rect -96 59751 -84 59785
rect 84 59751 96 59785
rect -96 59745 96 59751
rect -96 59677 96 59683
rect -96 59643 -84 59677
rect 84 59643 96 59677
rect -96 59637 96 59643
rect -152 59593 -106 59605
rect -152 59017 -146 59593
rect -112 59017 -106 59593
rect -152 59005 -106 59017
rect 106 59593 152 59605
rect 106 59017 112 59593
rect 146 59017 152 59593
rect 106 59005 152 59017
rect -96 58967 96 58973
rect -96 58933 -84 58967
rect 84 58933 96 58967
rect -96 58927 96 58933
rect -96 58859 96 58865
rect -96 58825 -84 58859
rect 84 58825 96 58859
rect -96 58819 96 58825
rect -152 58775 -106 58787
rect -152 58199 -146 58775
rect -112 58199 -106 58775
rect -152 58187 -106 58199
rect 106 58775 152 58787
rect 106 58199 112 58775
rect 146 58199 152 58775
rect 106 58187 152 58199
rect -96 58149 96 58155
rect -96 58115 -84 58149
rect 84 58115 96 58149
rect -96 58109 96 58115
rect -96 58041 96 58047
rect -96 58007 -84 58041
rect 84 58007 96 58041
rect -96 58001 96 58007
rect -152 57957 -106 57969
rect -152 57381 -146 57957
rect -112 57381 -106 57957
rect -152 57369 -106 57381
rect 106 57957 152 57969
rect 106 57381 112 57957
rect 146 57381 152 57957
rect 106 57369 152 57381
rect -96 57331 96 57337
rect -96 57297 -84 57331
rect 84 57297 96 57331
rect -96 57291 96 57297
rect -96 57223 96 57229
rect -96 57189 -84 57223
rect 84 57189 96 57223
rect -96 57183 96 57189
rect -152 57139 -106 57151
rect -152 56563 -146 57139
rect -112 56563 -106 57139
rect -152 56551 -106 56563
rect 106 57139 152 57151
rect 106 56563 112 57139
rect 146 56563 152 57139
rect 106 56551 152 56563
rect -96 56513 96 56519
rect -96 56479 -84 56513
rect 84 56479 96 56513
rect -96 56473 96 56479
rect -96 56405 96 56411
rect -96 56371 -84 56405
rect 84 56371 96 56405
rect -96 56365 96 56371
rect -152 56321 -106 56333
rect -152 55745 -146 56321
rect -112 55745 -106 56321
rect -152 55733 -106 55745
rect 106 56321 152 56333
rect 106 55745 112 56321
rect 146 55745 152 56321
rect 106 55733 152 55745
rect -96 55695 96 55701
rect -96 55661 -84 55695
rect 84 55661 96 55695
rect -96 55655 96 55661
rect -96 55587 96 55593
rect -96 55553 -84 55587
rect 84 55553 96 55587
rect -96 55547 96 55553
rect -152 55503 -106 55515
rect -152 54927 -146 55503
rect -112 54927 -106 55503
rect -152 54915 -106 54927
rect 106 55503 152 55515
rect 106 54927 112 55503
rect 146 54927 152 55503
rect 106 54915 152 54927
rect -96 54877 96 54883
rect -96 54843 -84 54877
rect 84 54843 96 54877
rect -96 54837 96 54843
rect -96 54769 96 54775
rect -96 54735 -84 54769
rect 84 54735 96 54769
rect -96 54729 96 54735
rect -152 54685 -106 54697
rect -152 54109 -146 54685
rect -112 54109 -106 54685
rect -152 54097 -106 54109
rect 106 54685 152 54697
rect 106 54109 112 54685
rect 146 54109 152 54685
rect 106 54097 152 54109
rect -96 54059 96 54065
rect -96 54025 -84 54059
rect 84 54025 96 54059
rect -96 54019 96 54025
rect -96 53951 96 53957
rect -96 53917 -84 53951
rect 84 53917 96 53951
rect -96 53911 96 53917
rect -152 53867 -106 53879
rect -152 53291 -146 53867
rect -112 53291 -106 53867
rect -152 53279 -106 53291
rect 106 53867 152 53879
rect 106 53291 112 53867
rect 146 53291 152 53867
rect 106 53279 152 53291
rect -96 53241 96 53247
rect -96 53207 -84 53241
rect 84 53207 96 53241
rect -96 53201 96 53207
rect -96 53133 96 53139
rect -96 53099 -84 53133
rect 84 53099 96 53133
rect -96 53093 96 53099
rect -152 53049 -106 53061
rect -152 52473 -146 53049
rect -112 52473 -106 53049
rect -152 52461 -106 52473
rect 106 53049 152 53061
rect 106 52473 112 53049
rect 146 52473 152 53049
rect 106 52461 152 52473
rect -96 52423 96 52429
rect -96 52389 -84 52423
rect 84 52389 96 52423
rect -96 52383 96 52389
rect -96 52315 96 52321
rect -96 52281 -84 52315
rect 84 52281 96 52315
rect -96 52275 96 52281
rect -152 52231 -106 52243
rect -152 51655 -146 52231
rect -112 51655 -106 52231
rect -152 51643 -106 51655
rect 106 52231 152 52243
rect 106 51655 112 52231
rect 146 51655 152 52231
rect 106 51643 152 51655
rect -96 51605 96 51611
rect -96 51571 -84 51605
rect 84 51571 96 51605
rect -96 51565 96 51571
rect -96 51497 96 51503
rect -96 51463 -84 51497
rect 84 51463 96 51497
rect -96 51457 96 51463
rect -152 51413 -106 51425
rect -152 50837 -146 51413
rect -112 50837 -106 51413
rect -152 50825 -106 50837
rect 106 51413 152 51425
rect 106 50837 112 51413
rect 146 50837 152 51413
rect 106 50825 152 50837
rect -96 50787 96 50793
rect -96 50753 -84 50787
rect 84 50753 96 50787
rect -96 50747 96 50753
rect -96 50679 96 50685
rect -96 50645 -84 50679
rect 84 50645 96 50679
rect -96 50639 96 50645
rect -152 50595 -106 50607
rect -152 50019 -146 50595
rect -112 50019 -106 50595
rect -152 50007 -106 50019
rect 106 50595 152 50607
rect 106 50019 112 50595
rect 146 50019 152 50595
rect 106 50007 152 50019
rect -96 49969 96 49975
rect -96 49935 -84 49969
rect 84 49935 96 49969
rect -96 49929 96 49935
rect -96 49861 96 49867
rect -96 49827 -84 49861
rect 84 49827 96 49861
rect -96 49821 96 49827
rect -152 49777 -106 49789
rect -152 49201 -146 49777
rect -112 49201 -106 49777
rect -152 49189 -106 49201
rect 106 49777 152 49789
rect 106 49201 112 49777
rect 146 49201 152 49777
rect 106 49189 152 49201
rect -96 49151 96 49157
rect -96 49117 -84 49151
rect 84 49117 96 49151
rect -96 49111 96 49117
rect -96 49043 96 49049
rect -96 49009 -84 49043
rect 84 49009 96 49043
rect -96 49003 96 49009
rect -152 48959 -106 48971
rect -152 48383 -146 48959
rect -112 48383 -106 48959
rect -152 48371 -106 48383
rect 106 48959 152 48971
rect 106 48383 112 48959
rect 146 48383 152 48959
rect 106 48371 152 48383
rect -96 48333 96 48339
rect -96 48299 -84 48333
rect 84 48299 96 48333
rect -96 48293 96 48299
rect -96 48225 96 48231
rect -96 48191 -84 48225
rect 84 48191 96 48225
rect -96 48185 96 48191
rect -152 48141 -106 48153
rect -152 47565 -146 48141
rect -112 47565 -106 48141
rect -152 47553 -106 47565
rect 106 48141 152 48153
rect 106 47565 112 48141
rect 146 47565 152 48141
rect 106 47553 152 47565
rect -96 47515 96 47521
rect -96 47481 -84 47515
rect 84 47481 96 47515
rect -96 47475 96 47481
rect -96 47407 96 47413
rect -96 47373 -84 47407
rect 84 47373 96 47407
rect -96 47367 96 47373
rect -152 47323 -106 47335
rect -152 46747 -146 47323
rect -112 46747 -106 47323
rect -152 46735 -106 46747
rect 106 47323 152 47335
rect 106 46747 112 47323
rect 146 46747 152 47323
rect 106 46735 152 46747
rect -96 46697 96 46703
rect -96 46663 -84 46697
rect 84 46663 96 46697
rect -96 46657 96 46663
rect -96 46589 96 46595
rect -96 46555 -84 46589
rect 84 46555 96 46589
rect -96 46549 96 46555
rect -152 46505 -106 46517
rect -152 45929 -146 46505
rect -112 45929 -106 46505
rect -152 45917 -106 45929
rect 106 46505 152 46517
rect 106 45929 112 46505
rect 146 45929 152 46505
rect 106 45917 152 45929
rect -96 45879 96 45885
rect -96 45845 -84 45879
rect 84 45845 96 45879
rect -96 45839 96 45845
rect -96 45771 96 45777
rect -96 45737 -84 45771
rect 84 45737 96 45771
rect -96 45731 96 45737
rect -152 45687 -106 45699
rect -152 45111 -146 45687
rect -112 45111 -106 45687
rect -152 45099 -106 45111
rect 106 45687 152 45699
rect 106 45111 112 45687
rect 146 45111 152 45687
rect 106 45099 152 45111
rect -96 45061 96 45067
rect -96 45027 -84 45061
rect 84 45027 96 45061
rect -96 45021 96 45027
rect -96 44953 96 44959
rect -96 44919 -84 44953
rect 84 44919 96 44953
rect -96 44913 96 44919
rect -152 44869 -106 44881
rect -152 44293 -146 44869
rect -112 44293 -106 44869
rect -152 44281 -106 44293
rect 106 44869 152 44881
rect 106 44293 112 44869
rect 146 44293 152 44869
rect 106 44281 152 44293
rect -96 44243 96 44249
rect -96 44209 -84 44243
rect 84 44209 96 44243
rect -96 44203 96 44209
rect -96 44135 96 44141
rect -96 44101 -84 44135
rect 84 44101 96 44135
rect -96 44095 96 44101
rect -152 44051 -106 44063
rect -152 43475 -146 44051
rect -112 43475 -106 44051
rect -152 43463 -106 43475
rect 106 44051 152 44063
rect 106 43475 112 44051
rect 146 43475 152 44051
rect 106 43463 152 43475
rect -96 43425 96 43431
rect -96 43391 -84 43425
rect 84 43391 96 43425
rect -96 43385 96 43391
rect -96 43317 96 43323
rect -96 43283 -84 43317
rect 84 43283 96 43317
rect -96 43277 96 43283
rect -152 43233 -106 43245
rect -152 42657 -146 43233
rect -112 42657 -106 43233
rect -152 42645 -106 42657
rect 106 43233 152 43245
rect 106 42657 112 43233
rect 146 42657 152 43233
rect 106 42645 152 42657
rect -96 42607 96 42613
rect -96 42573 -84 42607
rect 84 42573 96 42607
rect -96 42567 96 42573
rect -96 42499 96 42505
rect -96 42465 -84 42499
rect 84 42465 96 42499
rect -96 42459 96 42465
rect -152 42415 -106 42427
rect -152 41839 -146 42415
rect -112 41839 -106 42415
rect -152 41827 -106 41839
rect 106 42415 152 42427
rect 106 41839 112 42415
rect 146 41839 152 42415
rect 106 41827 152 41839
rect -96 41789 96 41795
rect -96 41755 -84 41789
rect 84 41755 96 41789
rect -96 41749 96 41755
rect -96 41681 96 41687
rect -96 41647 -84 41681
rect 84 41647 96 41681
rect -96 41641 96 41647
rect -152 41597 -106 41609
rect -152 41021 -146 41597
rect -112 41021 -106 41597
rect -152 41009 -106 41021
rect 106 41597 152 41609
rect 106 41021 112 41597
rect 146 41021 152 41597
rect 106 41009 152 41021
rect -96 40971 96 40977
rect -96 40937 -84 40971
rect 84 40937 96 40971
rect -96 40931 96 40937
rect -96 40863 96 40869
rect -96 40829 -84 40863
rect 84 40829 96 40863
rect -96 40823 96 40829
rect -152 40779 -106 40791
rect -152 40203 -146 40779
rect -112 40203 -106 40779
rect -152 40191 -106 40203
rect 106 40779 152 40791
rect 106 40203 112 40779
rect 146 40203 152 40779
rect 106 40191 152 40203
rect -96 40153 96 40159
rect -96 40119 -84 40153
rect 84 40119 96 40153
rect -96 40113 96 40119
rect -96 40045 96 40051
rect -96 40011 -84 40045
rect 84 40011 96 40045
rect -96 40005 96 40011
rect -152 39961 -106 39973
rect -152 39385 -146 39961
rect -112 39385 -106 39961
rect -152 39373 -106 39385
rect 106 39961 152 39973
rect 106 39385 112 39961
rect 146 39385 152 39961
rect 106 39373 152 39385
rect -96 39335 96 39341
rect -96 39301 -84 39335
rect 84 39301 96 39335
rect -96 39295 96 39301
rect -96 39227 96 39233
rect -96 39193 -84 39227
rect 84 39193 96 39227
rect -96 39187 96 39193
rect -152 39143 -106 39155
rect -152 38567 -146 39143
rect -112 38567 -106 39143
rect -152 38555 -106 38567
rect 106 39143 152 39155
rect 106 38567 112 39143
rect 146 38567 152 39143
rect 106 38555 152 38567
rect -96 38517 96 38523
rect -96 38483 -84 38517
rect 84 38483 96 38517
rect -96 38477 96 38483
rect -96 38409 96 38415
rect -96 38375 -84 38409
rect 84 38375 96 38409
rect -96 38369 96 38375
rect -152 38325 -106 38337
rect -152 37749 -146 38325
rect -112 37749 -106 38325
rect -152 37737 -106 37749
rect 106 38325 152 38337
rect 106 37749 112 38325
rect 146 37749 152 38325
rect 106 37737 152 37749
rect -96 37699 96 37705
rect -96 37665 -84 37699
rect 84 37665 96 37699
rect -96 37659 96 37665
rect -96 37591 96 37597
rect -96 37557 -84 37591
rect 84 37557 96 37591
rect -96 37551 96 37557
rect -152 37507 -106 37519
rect -152 36931 -146 37507
rect -112 36931 -106 37507
rect -152 36919 -106 36931
rect 106 37507 152 37519
rect 106 36931 112 37507
rect 146 36931 152 37507
rect 106 36919 152 36931
rect -96 36881 96 36887
rect -96 36847 -84 36881
rect 84 36847 96 36881
rect -96 36841 96 36847
rect -96 36773 96 36779
rect -96 36739 -84 36773
rect 84 36739 96 36773
rect -96 36733 96 36739
rect -152 36689 -106 36701
rect -152 36113 -146 36689
rect -112 36113 -106 36689
rect -152 36101 -106 36113
rect 106 36689 152 36701
rect 106 36113 112 36689
rect 146 36113 152 36689
rect 106 36101 152 36113
rect -96 36063 96 36069
rect -96 36029 -84 36063
rect 84 36029 96 36063
rect -96 36023 96 36029
rect -96 35955 96 35961
rect -96 35921 -84 35955
rect 84 35921 96 35955
rect -96 35915 96 35921
rect -152 35871 -106 35883
rect -152 35295 -146 35871
rect -112 35295 -106 35871
rect -152 35283 -106 35295
rect 106 35871 152 35883
rect 106 35295 112 35871
rect 146 35295 152 35871
rect 106 35283 152 35295
rect -96 35245 96 35251
rect -96 35211 -84 35245
rect 84 35211 96 35245
rect -96 35205 96 35211
rect -96 35137 96 35143
rect -96 35103 -84 35137
rect 84 35103 96 35137
rect -96 35097 96 35103
rect -152 35053 -106 35065
rect -152 34477 -146 35053
rect -112 34477 -106 35053
rect -152 34465 -106 34477
rect 106 35053 152 35065
rect 106 34477 112 35053
rect 146 34477 152 35053
rect 106 34465 152 34477
rect -96 34427 96 34433
rect -96 34393 -84 34427
rect 84 34393 96 34427
rect -96 34387 96 34393
rect -96 34319 96 34325
rect -96 34285 -84 34319
rect 84 34285 96 34319
rect -96 34279 96 34285
rect -152 34235 -106 34247
rect -152 33659 -146 34235
rect -112 33659 -106 34235
rect -152 33647 -106 33659
rect 106 34235 152 34247
rect 106 33659 112 34235
rect 146 33659 152 34235
rect 106 33647 152 33659
rect -96 33609 96 33615
rect -96 33575 -84 33609
rect 84 33575 96 33609
rect -96 33569 96 33575
rect -96 33501 96 33507
rect -96 33467 -84 33501
rect 84 33467 96 33501
rect -96 33461 96 33467
rect -152 33417 -106 33429
rect -152 32841 -146 33417
rect -112 32841 -106 33417
rect -152 32829 -106 32841
rect 106 33417 152 33429
rect 106 32841 112 33417
rect 146 32841 152 33417
rect 106 32829 152 32841
rect -96 32791 96 32797
rect -96 32757 -84 32791
rect 84 32757 96 32791
rect -96 32751 96 32757
rect -96 32683 96 32689
rect -96 32649 -84 32683
rect 84 32649 96 32683
rect -96 32643 96 32649
rect -152 32599 -106 32611
rect -152 32023 -146 32599
rect -112 32023 -106 32599
rect -152 32011 -106 32023
rect 106 32599 152 32611
rect 106 32023 112 32599
rect 146 32023 152 32599
rect 106 32011 152 32023
rect -96 31973 96 31979
rect -96 31939 -84 31973
rect 84 31939 96 31973
rect -96 31933 96 31939
rect -96 31865 96 31871
rect -96 31831 -84 31865
rect 84 31831 96 31865
rect -96 31825 96 31831
rect -152 31781 -106 31793
rect -152 31205 -146 31781
rect -112 31205 -106 31781
rect -152 31193 -106 31205
rect 106 31781 152 31793
rect 106 31205 112 31781
rect 146 31205 152 31781
rect 106 31193 152 31205
rect -96 31155 96 31161
rect -96 31121 -84 31155
rect 84 31121 96 31155
rect -96 31115 96 31121
rect -96 31047 96 31053
rect -96 31013 -84 31047
rect 84 31013 96 31047
rect -96 31007 96 31013
rect -152 30963 -106 30975
rect -152 30387 -146 30963
rect -112 30387 -106 30963
rect -152 30375 -106 30387
rect 106 30963 152 30975
rect 106 30387 112 30963
rect 146 30387 152 30963
rect 106 30375 152 30387
rect -96 30337 96 30343
rect -96 30303 -84 30337
rect 84 30303 96 30337
rect -96 30297 96 30303
rect -96 30229 96 30235
rect -96 30195 -84 30229
rect 84 30195 96 30229
rect -96 30189 96 30195
rect -152 30145 -106 30157
rect -152 29569 -146 30145
rect -112 29569 -106 30145
rect -152 29557 -106 29569
rect 106 30145 152 30157
rect 106 29569 112 30145
rect 146 29569 152 30145
rect 106 29557 152 29569
rect -96 29519 96 29525
rect -96 29485 -84 29519
rect 84 29485 96 29519
rect -96 29479 96 29485
rect -96 29411 96 29417
rect -96 29377 -84 29411
rect 84 29377 96 29411
rect -96 29371 96 29377
rect -152 29327 -106 29339
rect -152 28751 -146 29327
rect -112 28751 -106 29327
rect -152 28739 -106 28751
rect 106 29327 152 29339
rect 106 28751 112 29327
rect 146 28751 152 29327
rect 106 28739 152 28751
rect -96 28701 96 28707
rect -96 28667 -84 28701
rect 84 28667 96 28701
rect -96 28661 96 28667
rect -96 28593 96 28599
rect -96 28559 -84 28593
rect 84 28559 96 28593
rect -96 28553 96 28559
rect -152 28509 -106 28521
rect -152 27933 -146 28509
rect -112 27933 -106 28509
rect -152 27921 -106 27933
rect 106 28509 152 28521
rect 106 27933 112 28509
rect 146 27933 152 28509
rect 106 27921 152 27933
rect -96 27883 96 27889
rect -96 27849 -84 27883
rect 84 27849 96 27883
rect -96 27843 96 27849
rect -96 27775 96 27781
rect -96 27741 -84 27775
rect 84 27741 96 27775
rect -96 27735 96 27741
rect -152 27691 -106 27703
rect -152 27115 -146 27691
rect -112 27115 -106 27691
rect -152 27103 -106 27115
rect 106 27691 152 27703
rect 106 27115 112 27691
rect 146 27115 152 27691
rect 106 27103 152 27115
rect -96 27065 96 27071
rect -96 27031 -84 27065
rect 84 27031 96 27065
rect -96 27025 96 27031
rect -96 26957 96 26963
rect -96 26923 -84 26957
rect 84 26923 96 26957
rect -96 26917 96 26923
rect -152 26873 -106 26885
rect -152 26297 -146 26873
rect -112 26297 -106 26873
rect -152 26285 -106 26297
rect 106 26873 152 26885
rect 106 26297 112 26873
rect 146 26297 152 26873
rect 106 26285 152 26297
rect -96 26247 96 26253
rect -96 26213 -84 26247
rect 84 26213 96 26247
rect -96 26207 96 26213
rect -96 26139 96 26145
rect -96 26105 -84 26139
rect 84 26105 96 26139
rect -96 26099 96 26105
rect -152 26055 -106 26067
rect -152 25479 -146 26055
rect -112 25479 -106 26055
rect -152 25467 -106 25479
rect 106 26055 152 26067
rect 106 25479 112 26055
rect 146 25479 152 26055
rect 106 25467 152 25479
rect -96 25429 96 25435
rect -96 25395 -84 25429
rect 84 25395 96 25429
rect -96 25389 96 25395
rect -96 25321 96 25327
rect -96 25287 -84 25321
rect 84 25287 96 25321
rect -96 25281 96 25287
rect -152 25237 -106 25249
rect -152 24661 -146 25237
rect -112 24661 -106 25237
rect -152 24649 -106 24661
rect 106 25237 152 25249
rect 106 24661 112 25237
rect 146 24661 152 25237
rect 106 24649 152 24661
rect -96 24611 96 24617
rect -96 24577 -84 24611
rect 84 24577 96 24611
rect -96 24571 96 24577
rect -96 24503 96 24509
rect -96 24469 -84 24503
rect 84 24469 96 24503
rect -96 24463 96 24469
rect -152 24419 -106 24431
rect -152 23843 -146 24419
rect -112 23843 -106 24419
rect -152 23831 -106 23843
rect 106 24419 152 24431
rect 106 23843 112 24419
rect 146 23843 152 24419
rect 106 23831 152 23843
rect -96 23793 96 23799
rect -96 23759 -84 23793
rect 84 23759 96 23793
rect -96 23753 96 23759
rect -96 23685 96 23691
rect -96 23651 -84 23685
rect 84 23651 96 23685
rect -96 23645 96 23651
rect -152 23601 -106 23613
rect -152 23025 -146 23601
rect -112 23025 -106 23601
rect -152 23013 -106 23025
rect 106 23601 152 23613
rect 106 23025 112 23601
rect 146 23025 152 23601
rect 106 23013 152 23025
rect -96 22975 96 22981
rect -96 22941 -84 22975
rect 84 22941 96 22975
rect -96 22935 96 22941
rect -96 22867 96 22873
rect -96 22833 -84 22867
rect 84 22833 96 22867
rect -96 22827 96 22833
rect -152 22783 -106 22795
rect -152 22207 -146 22783
rect -112 22207 -106 22783
rect -152 22195 -106 22207
rect 106 22783 152 22795
rect 106 22207 112 22783
rect 146 22207 152 22783
rect 106 22195 152 22207
rect -96 22157 96 22163
rect -96 22123 -84 22157
rect 84 22123 96 22157
rect -96 22117 96 22123
rect -96 22049 96 22055
rect -96 22015 -84 22049
rect 84 22015 96 22049
rect -96 22009 96 22015
rect -152 21965 -106 21977
rect -152 21389 -146 21965
rect -112 21389 -106 21965
rect -152 21377 -106 21389
rect 106 21965 152 21977
rect 106 21389 112 21965
rect 146 21389 152 21965
rect 106 21377 152 21389
rect -96 21339 96 21345
rect -96 21305 -84 21339
rect 84 21305 96 21339
rect -96 21299 96 21305
rect -96 21231 96 21237
rect -96 21197 -84 21231
rect 84 21197 96 21231
rect -96 21191 96 21197
rect -152 21147 -106 21159
rect -152 20571 -146 21147
rect -112 20571 -106 21147
rect -152 20559 -106 20571
rect 106 21147 152 21159
rect 106 20571 112 21147
rect 146 20571 152 21147
rect 106 20559 152 20571
rect -96 20521 96 20527
rect -96 20487 -84 20521
rect 84 20487 96 20521
rect -96 20481 96 20487
rect -96 20413 96 20419
rect -96 20379 -84 20413
rect 84 20379 96 20413
rect -96 20373 96 20379
rect -152 20329 -106 20341
rect -152 19753 -146 20329
rect -112 19753 -106 20329
rect -152 19741 -106 19753
rect 106 20329 152 20341
rect 106 19753 112 20329
rect 146 19753 152 20329
rect 106 19741 152 19753
rect -96 19703 96 19709
rect -96 19669 -84 19703
rect 84 19669 96 19703
rect -96 19663 96 19669
rect -96 19595 96 19601
rect -96 19561 -84 19595
rect 84 19561 96 19595
rect -96 19555 96 19561
rect -152 19511 -106 19523
rect -152 18935 -146 19511
rect -112 18935 -106 19511
rect -152 18923 -106 18935
rect 106 19511 152 19523
rect 106 18935 112 19511
rect 146 18935 152 19511
rect 106 18923 152 18935
rect -96 18885 96 18891
rect -96 18851 -84 18885
rect 84 18851 96 18885
rect -96 18845 96 18851
rect -96 18777 96 18783
rect -96 18743 -84 18777
rect 84 18743 96 18777
rect -96 18737 96 18743
rect -152 18693 -106 18705
rect -152 18117 -146 18693
rect -112 18117 -106 18693
rect -152 18105 -106 18117
rect 106 18693 152 18705
rect 106 18117 112 18693
rect 146 18117 152 18693
rect 106 18105 152 18117
rect -96 18067 96 18073
rect -96 18033 -84 18067
rect 84 18033 96 18067
rect -96 18027 96 18033
rect -96 17959 96 17965
rect -96 17925 -84 17959
rect 84 17925 96 17959
rect -96 17919 96 17925
rect -152 17875 -106 17887
rect -152 17299 -146 17875
rect -112 17299 -106 17875
rect -152 17287 -106 17299
rect 106 17875 152 17887
rect 106 17299 112 17875
rect 146 17299 152 17875
rect 106 17287 152 17299
rect -96 17249 96 17255
rect -96 17215 -84 17249
rect 84 17215 96 17249
rect -96 17209 96 17215
rect -96 17141 96 17147
rect -96 17107 -84 17141
rect 84 17107 96 17141
rect -96 17101 96 17107
rect -152 17057 -106 17069
rect -152 16481 -146 17057
rect -112 16481 -106 17057
rect -152 16469 -106 16481
rect 106 17057 152 17069
rect 106 16481 112 17057
rect 146 16481 152 17057
rect 106 16469 152 16481
rect -96 16431 96 16437
rect -96 16397 -84 16431
rect 84 16397 96 16431
rect -96 16391 96 16397
rect -96 16323 96 16329
rect -96 16289 -84 16323
rect 84 16289 96 16323
rect -96 16283 96 16289
rect -152 16239 -106 16251
rect -152 15663 -146 16239
rect -112 15663 -106 16239
rect -152 15651 -106 15663
rect 106 16239 152 16251
rect 106 15663 112 16239
rect 146 15663 152 16239
rect 106 15651 152 15663
rect -96 15613 96 15619
rect -96 15579 -84 15613
rect 84 15579 96 15613
rect -96 15573 96 15579
rect -96 15505 96 15511
rect -96 15471 -84 15505
rect 84 15471 96 15505
rect -96 15465 96 15471
rect -152 15421 -106 15433
rect -152 14845 -146 15421
rect -112 14845 -106 15421
rect -152 14833 -106 14845
rect 106 15421 152 15433
rect 106 14845 112 15421
rect 146 14845 152 15421
rect 106 14833 152 14845
rect -96 14795 96 14801
rect -96 14761 -84 14795
rect 84 14761 96 14795
rect -96 14755 96 14761
rect -96 14687 96 14693
rect -96 14653 -84 14687
rect 84 14653 96 14687
rect -96 14647 96 14653
rect -152 14603 -106 14615
rect -152 14027 -146 14603
rect -112 14027 -106 14603
rect -152 14015 -106 14027
rect 106 14603 152 14615
rect 106 14027 112 14603
rect 146 14027 152 14603
rect 106 14015 152 14027
rect -96 13977 96 13983
rect -96 13943 -84 13977
rect 84 13943 96 13977
rect -96 13937 96 13943
rect -96 13869 96 13875
rect -96 13835 -84 13869
rect 84 13835 96 13869
rect -96 13829 96 13835
rect -152 13785 -106 13797
rect -152 13209 -146 13785
rect -112 13209 -106 13785
rect -152 13197 -106 13209
rect 106 13785 152 13797
rect 106 13209 112 13785
rect 146 13209 152 13785
rect 106 13197 152 13209
rect -96 13159 96 13165
rect -96 13125 -84 13159
rect 84 13125 96 13159
rect -96 13119 96 13125
rect -96 13051 96 13057
rect -96 13017 -84 13051
rect 84 13017 96 13051
rect -96 13011 96 13017
rect -152 12967 -106 12979
rect -152 12391 -146 12967
rect -112 12391 -106 12967
rect -152 12379 -106 12391
rect 106 12967 152 12979
rect 106 12391 112 12967
rect 146 12391 152 12967
rect 106 12379 152 12391
rect -96 12341 96 12347
rect -96 12307 -84 12341
rect 84 12307 96 12341
rect -96 12301 96 12307
rect -96 12233 96 12239
rect -96 12199 -84 12233
rect 84 12199 96 12233
rect -96 12193 96 12199
rect -152 12149 -106 12161
rect -152 11573 -146 12149
rect -112 11573 -106 12149
rect -152 11561 -106 11573
rect 106 12149 152 12161
rect 106 11573 112 12149
rect 146 11573 152 12149
rect 106 11561 152 11573
rect -96 11523 96 11529
rect -96 11489 -84 11523
rect 84 11489 96 11523
rect -96 11483 96 11489
rect -96 11415 96 11421
rect -96 11381 -84 11415
rect 84 11381 96 11415
rect -96 11375 96 11381
rect -152 11331 -106 11343
rect -152 10755 -146 11331
rect -112 10755 -106 11331
rect -152 10743 -106 10755
rect 106 11331 152 11343
rect 106 10755 112 11331
rect 146 10755 152 11331
rect 106 10743 152 10755
rect -96 10705 96 10711
rect -96 10671 -84 10705
rect 84 10671 96 10705
rect -96 10665 96 10671
rect -96 10597 96 10603
rect -96 10563 -84 10597
rect 84 10563 96 10597
rect -96 10557 96 10563
rect -152 10513 -106 10525
rect -152 9937 -146 10513
rect -112 9937 -106 10513
rect -152 9925 -106 9937
rect 106 10513 152 10525
rect 106 9937 112 10513
rect 146 9937 152 10513
rect 106 9925 152 9937
rect -96 9887 96 9893
rect -96 9853 -84 9887
rect 84 9853 96 9887
rect -96 9847 96 9853
rect -96 9779 96 9785
rect -96 9745 -84 9779
rect 84 9745 96 9779
rect -96 9739 96 9745
rect -152 9695 -106 9707
rect -152 9119 -146 9695
rect -112 9119 -106 9695
rect -152 9107 -106 9119
rect 106 9695 152 9707
rect 106 9119 112 9695
rect 146 9119 152 9695
rect 106 9107 152 9119
rect -96 9069 96 9075
rect -96 9035 -84 9069
rect 84 9035 96 9069
rect -96 9029 96 9035
rect -96 8961 96 8967
rect -96 8927 -84 8961
rect 84 8927 96 8961
rect -96 8921 96 8927
rect -152 8877 -106 8889
rect -152 8301 -146 8877
rect -112 8301 -106 8877
rect -152 8289 -106 8301
rect 106 8877 152 8889
rect 106 8301 112 8877
rect 146 8301 152 8877
rect 106 8289 152 8301
rect -96 8251 96 8257
rect -96 8217 -84 8251
rect 84 8217 96 8251
rect -96 8211 96 8217
rect -96 8143 96 8149
rect -96 8109 -84 8143
rect 84 8109 96 8143
rect -96 8103 96 8109
rect -152 8059 -106 8071
rect -152 7483 -146 8059
rect -112 7483 -106 8059
rect -152 7471 -106 7483
rect 106 8059 152 8071
rect 106 7483 112 8059
rect 146 7483 152 8059
rect 106 7471 152 7483
rect -96 7433 96 7439
rect -96 7399 -84 7433
rect 84 7399 96 7433
rect -96 7393 96 7399
rect -96 7325 96 7331
rect -96 7291 -84 7325
rect 84 7291 96 7325
rect -96 7285 96 7291
rect -152 7241 -106 7253
rect -152 6665 -146 7241
rect -112 6665 -106 7241
rect -152 6653 -106 6665
rect 106 7241 152 7253
rect 106 6665 112 7241
rect 146 6665 152 7241
rect 106 6653 152 6665
rect -96 6615 96 6621
rect -96 6581 -84 6615
rect 84 6581 96 6615
rect -96 6575 96 6581
rect -96 6507 96 6513
rect -96 6473 -84 6507
rect 84 6473 96 6507
rect -96 6467 96 6473
rect -152 6423 -106 6435
rect -152 5847 -146 6423
rect -112 5847 -106 6423
rect -152 5835 -106 5847
rect 106 6423 152 6435
rect 106 5847 112 6423
rect 146 5847 152 6423
rect 106 5835 152 5847
rect -96 5797 96 5803
rect -96 5763 -84 5797
rect 84 5763 96 5797
rect -96 5757 96 5763
rect -96 5689 96 5695
rect -96 5655 -84 5689
rect 84 5655 96 5689
rect -96 5649 96 5655
rect -152 5605 -106 5617
rect -152 5029 -146 5605
rect -112 5029 -106 5605
rect -152 5017 -106 5029
rect 106 5605 152 5617
rect 106 5029 112 5605
rect 146 5029 152 5605
rect 106 5017 152 5029
rect -96 4979 96 4985
rect -96 4945 -84 4979
rect 84 4945 96 4979
rect -96 4939 96 4945
rect -96 4871 96 4877
rect -96 4837 -84 4871
rect 84 4837 96 4871
rect -96 4831 96 4837
rect -152 4787 -106 4799
rect -152 4211 -146 4787
rect -112 4211 -106 4787
rect -152 4199 -106 4211
rect 106 4787 152 4799
rect 106 4211 112 4787
rect 146 4211 152 4787
rect 106 4199 152 4211
rect -96 4161 96 4167
rect -96 4127 -84 4161
rect 84 4127 96 4161
rect -96 4121 96 4127
rect -96 4053 96 4059
rect -96 4019 -84 4053
rect 84 4019 96 4053
rect -96 4013 96 4019
rect -152 3969 -106 3981
rect -152 3393 -146 3969
rect -112 3393 -106 3969
rect -152 3381 -106 3393
rect 106 3969 152 3981
rect 106 3393 112 3969
rect 146 3393 152 3969
rect 106 3381 152 3393
rect -96 3343 96 3349
rect -96 3309 -84 3343
rect 84 3309 96 3343
rect -96 3303 96 3309
rect -96 3235 96 3241
rect -96 3201 -84 3235
rect 84 3201 96 3235
rect -96 3195 96 3201
rect -152 3151 -106 3163
rect -152 2575 -146 3151
rect -112 2575 -106 3151
rect -152 2563 -106 2575
rect 106 3151 152 3163
rect 106 2575 112 3151
rect 146 2575 152 3151
rect 106 2563 152 2575
rect -96 2525 96 2531
rect -96 2491 -84 2525
rect 84 2491 96 2525
rect -96 2485 96 2491
rect -96 2417 96 2423
rect -96 2383 -84 2417
rect 84 2383 96 2417
rect -96 2377 96 2383
rect -152 2333 -106 2345
rect -152 1757 -146 2333
rect -112 1757 -106 2333
rect -152 1745 -106 1757
rect 106 2333 152 2345
rect 106 1757 112 2333
rect 146 1757 152 2333
rect 106 1745 152 1757
rect -96 1707 96 1713
rect -96 1673 -84 1707
rect 84 1673 96 1707
rect -96 1667 96 1673
rect -96 1599 96 1605
rect -96 1565 -84 1599
rect 84 1565 96 1599
rect -96 1559 96 1565
rect -152 1515 -106 1527
rect -152 939 -146 1515
rect -112 939 -106 1515
rect -152 927 -106 939
rect 106 1515 152 1527
rect 106 939 112 1515
rect 146 939 152 1515
rect 106 927 152 939
rect -96 889 96 895
rect -96 855 -84 889
rect 84 855 96 889
rect -96 849 96 855
rect -96 781 96 787
rect -96 747 -84 781
rect 84 747 96 781
rect -96 741 96 747
rect -152 697 -106 709
rect -152 121 -146 697
rect -112 121 -106 697
rect -152 109 -106 121
rect 106 697 152 709
rect 106 121 112 697
rect 146 121 152 697
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -697 -146 -121
rect -112 -697 -106 -121
rect -152 -709 -106 -697
rect 106 -121 152 -109
rect 106 -697 112 -121
rect 146 -697 152 -121
rect 106 -709 152 -697
rect -96 -747 96 -741
rect -96 -781 -84 -747
rect 84 -781 96 -747
rect -96 -787 96 -781
rect -96 -855 96 -849
rect -96 -889 -84 -855
rect 84 -889 96 -855
rect -96 -895 96 -889
rect -152 -939 -106 -927
rect -152 -1515 -146 -939
rect -112 -1515 -106 -939
rect -152 -1527 -106 -1515
rect 106 -939 152 -927
rect 106 -1515 112 -939
rect 146 -1515 152 -939
rect 106 -1527 152 -1515
rect -96 -1565 96 -1559
rect -96 -1599 -84 -1565
rect 84 -1599 96 -1565
rect -96 -1605 96 -1599
rect -96 -1673 96 -1667
rect -96 -1707 -84 -1673
rect 84 -1707 96 -1673
rect -96 -1713 96 -1707
rect -152 -1757 -106 -1745
rect -152 -2333 -146 -1757
rect -112 -2333 -106 -1757
rect -152 -2345 -106 -2333
rect 106 -1757 152 -1745
rect 106 -2333 112 -1757
rect 146 -2333 152 -1757
rect 106 -2345 152 -2333
rect -96 -2383 96 -2377
rect -96 -2417 -84 -2383
rect 84 -2417 96 -2383
rect -96 -2423 96 -2417
rect -96 -2491 96 -2485
rect -96 -2525 -84 -2491
rect 84 -2525 96 -2491
rect -96 -2531 96 -2525
rect -152 -2575 -106 -2563
rect -152 -3151 -146 -2575
rect -112 -3151 -106 -2575
rect -152 -3163 -106 -3151
rect 106 -2575 152 -2563
rect 106 -3151 112 -2575
rect 146 -3151 152 -2575
rect 106 -3163 152 -3151
rect -96 -3201 96 -3195
rect -96 -3235 -84 -3201
rect 84 -3235 96 -3201
rect -96 -3241 96 -3235
rect -96 -3309 96 -3303
rect -96 -3343 -84 -3309
rect 84 -3343 96 -3309
rect -96 -3349 96 -3343
rect -152 -3393 -106 -3381
rect -152 -3969 -146 -3393
rect -112 -3969 -106 -3393
rect -152 -3981 -106 -3969
rect 106 -3393 152 -3381
rect 106 -3969 112 -3393
rect 146 -3969 152 -3393
rect 106 -3981 152 -3969
rect -96 -4019 96 -4013
rect -96 -4053 -84 -4019
rect 84 -4053 96 -4019
rect -96 -4059 96 -4053
rect -96 -4127 96 -4121
rect -96 -4161 -84 -4127
rect 84 -4161 96 -4127
rect -96 -4167 96 -4161
rect -152 -4211 -106 -4199
rect -152 -4787 -146 -4211
rect -112 -4787 -106 -4211
rect -152 -4799 -106 -4787
rect 106 -4211 152 -4199
rect 106 -4787 112 -4211
rect 146 -4787 152 -4211
rect 106 -4799 152 -4787
rect -96 -4837 96 -4831
rect -96 -4871 -84 -4837
rect 84 -4871 96 -4837
rect -96 -4877 96 -4871
rect -96 -4945 96 -4939
rect -96 -4979 -84 -4945
rect 84 -4979 96 -4945
rect -96 -4985 96 -4979
rect -152 -5029 -106 -5017
rect -152 -5605 -146 -5029
rect -112 -5605 -106 -5029
rect -152 -5617 -106 -5605
rect 106 -5029 152 -5017
rect 106 -5605 112 -5029
rect 146 -5605 152 -5029
rect 106 -5617 152 -5605
rect -96 -5655 96 -5649
rect -96 -5689 -84 -5655
rect 84 -5689 96 -5655
rect -96 -5695 96 -5689
rect -96 -5763 96 -5757
rect -96 -5797 -84 -5763
rect 84 -5797 96 -5763
rect -96 -5803 96 -5797
rect -152 -5847 -106 -5835
rect -152 -6423 -146 -5847
rect -112 -6423 -106 -5847
rect -152 -6435 -106 -6423
rect 106 -5847 152 -5835
rect 106 -6423 112 -5847
rect 146 -6423 152 -5847
rect 106 -6435 152 -6423
rect -96 -6473 96 -6467
rect -96 -6507 -84 -6473
rect 84 -6507 96 -6473
rect -96 -6513 96 -6507
rect -96 -6581 96 -6575
rect -96 -6615 -84 -6581
rect 84 -6615 96 -6581
rect -96 -6621 96 -6615
rect -152 -6665 -106 -6653
rect -152 -7241 -146 -6665
rect -112 -7241 -106 -6665
rect -152 -7253 -106 -7241
rect 106 -6665 152 -6653
rect 106 -7241 112 -6665
rect 146 -7241 152 -6665
rect 106 -7253 152 -7241
rect -96 -7291 96 -7285
rect -96 -7325 -84 -7291
rect 84 -7325 96 -7291
rect -96 -7331 96 -7325
rect -96 -7399 96 -7393
rect -96 -7433 -84 -7399
rect 84 -7433 96 -7399
rect -96 -7439 96 -7433
rect -152 -7483 -106 -7471
rect -152 -8059 -146 -7483
rect -112 -8059 -106 -7483
rect -152 -8071 -106 -8059
rect 106 -7483 152 -7471
rect 106 -8059 112 -7483
rect 146 -8059 152 -7483
rect 106 -8071 152 -8059
rect -96 -8109 96 -8103
rect -96 -8143 -84 -8109
rect 84 -8143 96 -8109
rect -96 -8149 96 -8143
rect -96 -8217 96 -8211
rect -96 -8251 -84 -8217
rect 84 -8251 96 -8217
rect -96 -8257 96 -8251
rect -152 -8301 -106 -8289
rect -152 -8877 -146 -8301
rect -112 -8877 -106 -8301
rect -152 -8889 -106 -8877
rect 106 -8301 152 -8289
rect 106 -8877 112 -8301
rect 146 -8877 152 -8301
rect 106 -8889 152 -8877
rect -96 -8927 96 -8921
rect -96 -8961 -84 -8927
rect 84 -8961 96 -8927
rect -96 -8967 96 -8961
rect -96 -9035 96 -9029
rect -96 -9069 -84 -9035
rect 84 -9069 96 -9035
rect -96 -9075 96 -9069
rect -152 -9119 -106 -9107
rect -152 -9695 -146 -9119
rect -112 -9695 -106 -9119
rect -152 -9707 -106 -9695
rect 106 -9119 152 -9107
rect 106 -9695 112 -9119
rect 146 -9695 152 -9119
rect 106 -9707 152 -9695
rect -96 -9745 96 -9739
rect -96 -9779 -84 -9745
rect 84 -9779 96 -9745
rect -96 -9785 96 -9779
rect -96 -9853 96 -9847
rect -96 -9887 -84 -9853
rect 84 -9887 96 -9853
rect -96 -9893 96 -9887
rect -152 -9937 -106 -9925
rect -152 -10513 -146 -9937
rect -112 -10513 -106 -9937
rect -152 -10525 -106 -10513
rect 106 -9937 152 -9925
rect 106 -10513 112 -9937
rect 146 -10513 152 -9937
rect 106 -10525 152 -10513
rect -96 -10563 96 -10557
rect -96 -10597 -84 -10563
rect 84 -10597 96 -10563
rect -96 -10603 96 -10597
rect -96 -10671 96 -10665
rect -96 -10705 -84 -10671
rect 84 -10705 96 -10671
rect -96 -10711 96 -10705
rect -152 -10755 -106 -10743
rect -152 -11331 -146 -10755
rect -112 -11331 -106 -10755
rect -152 -11343 -106 -11331
rect 106 -10755 152 -10743
rect 106 -11331 112 -10755
rect 146 -11331 152 -10755
rect 106 -11343 152 -11331
rect -96 -11381 96 -11375
rect -96 -11415 -84 -11381
rect 84 -11415 96 -11381
rect -96 -11421 96 -11415
rect -96 -11489 96 -11483
rect -96 -11523 -84 -11489
rect 84 -11523 96 -11489
rect -96 -11529 96 -11523
rect -152 -11573 -106 -11561
rect -152 -12149 -146 -11573
rect -112 -12149 -106 -11573
rect -152 -12161 -106 -12149
rect 106 -11573 152 -11561
rect 106 -12149 112 -11573
rect 146 -12149 152 -11573
rect 106 -12161 152 -12149
rect -96 -12199 96 -12193
rect -96 -12233 -84 -12199
rect 84 -12233 96 -12199
rect -96 -12239 96 -12233
rect -96 -12307 96 -12301
rect -96 -12341 -84 -12307
rect 84 -12341 96 -12307
rect -96 -12347 96 -12341
rect -152 -12391 -106 -12379
rect -152 -12967 -146 -12391
rect -112 -12967 -106 -12391
rect -152 -12979 -106 -12967
rect 106 -12391 152 -12379
rect 106 -12967 112 -12391
rect 146 -12967 152 -12391
rect 106 -12979 152 -12967
rect -96 -13017 96 -13011
rect -96 -13051 -84 -13017
rect 84 -13051 96 -13017
rect -96 -13057 96 -13051
rect -96 -13125 96 -13119
rect -96 -13159 -84 -13125
rect 84 -13159 96 -13125
rect -96 -13165 96 -13159
rect -152 -13209 -106 -13197
rect -152 -13785 -146 -13209
rect -112 -13785 -106 -13209
rect -152 -13797 -106 -13785
rect 106 -13209 152 -13197
rect 106 -13785 112 -13209
rect 146 -13785 152 -13209
rect 106 -13797 152 -13785
rect -96 -13835 96 -13829
rect -96 -13869 -84 -13835
rect 84 -13869 96 -13835
rect -96 -13875 96 -13869
rect -96 -13943 96 -13937
rect -96 -13977 -84 -13943
rect 84 -13977 96 -13943
rect -96 -13983 96 -13977
rect -152 -14027 -106 -14015
rect -152 -14603 -146 -14027
rect -112 -14603 -106 -14027
rect -152 -14615 -106 -14603
rect 106 -14027 152 -14015
rect 106 -14603 112 -14027
rect 146 -14603 152 -14027
rect 106 -14615 152 -14603
rect -96 -14653 96 -14647
rect -96 -14687 -84 -14653
rect 84 -14687 96 -14653
rect -96 -14693 96 -14687
rect -96 -14761 96 -14755
rect -96 -14795 -84 -14761
rect 84 -14795 96 -14761
rect -96 -14801 96 -14795
rect -152 -14845 -106 -14833
rect -152 -15421 -146 -14845
rect -112 -15421 -106 -14845
rect -152 -15433 -106 -15421
rect 106 -14845 152 -14833
rect 106 -15421 112 -14845
rect 146 -15421 152 -14845
rect 106 -15433 152 -15421
rect -96 -15471 96 -15465
rect -96 -15505 -84 -15471
rect 84 -15505 96 -15471
rect -96 -15511 96 -15505
rect -96 -15579 96 -15573
rect -96 -15613 -84 -15579
rect 84 -15613 96 -15579
rect -96 -15619 96 -15613
rect -152 -15663 -106 -15651
rect -152 -16239 -146 -15663
rect -112 -16239 -106 -15663
rect -152 -16251 -106 -16239
rect 106 -15663 152 -15651
rect 106 -16239 112 -15663
rect 146 -16239 152 -15663
rect 106 -16251 152 -16239
rect -96 -16289 96 -16283
rect -96 -16323 -84 -16289
rect 84 -16323 96 -16289
rect -96 -16329 96 -16323
rect -96 -16397 96 -16391
rect -96 -16431 -84 -16397
rect 84 -16431 96 -16397
rect -96 -16437 96 -16431
rect -152 -16481 -106 -16469
rect -152 -17057 -146 -16481
rect -112 -17057 -106 -16481
rect -152 -17069 -106 -17057
rect 106 -16481 152 -16469
rect 106 -17057 112 -16481
rect 146 -17057 152 -16481
rect 106 -17069 152 -17057
rect -96 -17107 96 -17101
rect -96 -17141 -84 -17107
rect 84 -17141 96 -17107
rect -96 -17147 96 -17141
rect -96 -17215 96 -17209
rect -96 -17249 -84 -17215
rect 84 -17249 96 -17215
rect -96 -17255 96 -17249
rect -152 -17299 -106 -17287
rect -152 -17875 -146 -17299
rect -112 -17875 -106 -17299
rect -152 -17887 -106 -17875
rect 106 -17299 152 -17287
rect 106 -17875 112 -17299
rect 146 -17875 152 -17299
rect 106 -17887 152 -17875
rect -96 -17925 96 -17919
rect -96 -17959 -84 -17925
rect 84 -17959 96 -17925
rect -96 -17965 96 -17959
rect -96 -18033 96 -18027
rect -96 -18067 -84 -18033
rect 84 -18067 96 -18033
rect -96 -18073 96 -18067
rect -152 -18117 -106 -18105
rect -152 -18693 -146 -18117
rect -112 -18693 -106 -18117
rect -152 -18705 -106 -18693
rect 106 -18117 152 -18105
rect 106 -18693 112 -18117
rect 146 -18693 152 -18117
rect 106 -18705 152 -18693
rect -96 -18743 96 -18737
rect -96 -18777 -84 -18743
rect 84 -18777 96 -18743
rect -96 -18783 96 -18777
rect -96 -18851 96 -18845
rect -96 -18885 -84 -18851
rect 84 -18885 96 -18851
rect -96 -18891 96 -18885
rect -152 -18935 -106 -18923
rect -152 -19511 -146 -18935
rect -112 -19511 -106 -18935
rect -152 -19523 -106 -19511
rect 106 -18935 152 -18923
rect 106 -19511 112 -18935
rect 146 -19511 152 -18935
rect 106 -19523 152 -19511
rect -96 -19561 96 -19555
rect -96 -19595 -84 -19561
rect 84 -19595 96 -19561
rect -96 -19601 96 -19595
rect -96 -19669 96 -19663
rect -96 -19703 -84 -19669
rect 84 -19703 96 -19669
rect -96 -19709 96 -19703
rect -152 -19753 -106 -19741
rect -152 -20329 -146 -19753
rect -112 -20329 -106 -19753
rect -152 -20341 -106 -20329
rect 106 -19753 152 -19741
rect 106 -20329 112 -19753
rect 146 -20329 152 -19753
rect 106 -20341 152 -20329
rect -96 -20379 96 -20373
rect -96 -20413 -84 -20379
rect 84 -20413 96 -20379
rect -96 -20419 96 -20413
rect -96 -20487 96 -20481
rect -96 -20521 -84 -20487
rect 84 -20521 96 -20487
rect -96 -20527 96 -20521
rect -152 -20571 -106 -20559
rect -152 -21147 -146 -20571
rect -112 -21147 -106 -20571
rect -152 -21159 -106 -21147
rect 106 -20571 152 -20559
rect 106 -21147 112 -20571
rect 146 -21147 152 -20571
rect 106 -21159 152 -21147
rect -96 -21197 96 -21191
rect -96 -21231 -84 -21197
rect 84 -21231 96 -21197
rect -96 -21237 96 -21231
rect -96 -21305 96 -21299
rect -96 -21339 -84 -21305
rect 84 -21339 96 -21305
rect -96 -21345 96 -21339
rect -152 -21389 -106 -21377
rect -152 -21965 -146 -21389
rect -112 -21965 -106 -21389
rect -152 -21977 -106 -21965
rect 106 -21389 152 -21377
rect 106 -21965 112 -21389
rect 146 -21965 152 -21389
rect 106 -21977 152 -21965
rect -96 -22015 96 -22009
rect -96 -22049 -84 -22015
rect 84 -22049 96 -22015
rect -96 -22055 96 -22049
rect -96 -22123 96 -22117
rect -96 -22157 -84 -22123
rect 84 -22157 96 -22123
rect -96 -22163 96 -22157
rect -152 -22207 -106 -22195
rect -152 -22783 -146 -22207
rect -112 -22783 -106 -22207
rect -152 -22795 -106 -22783
rect 106 -22207 152 -22195
rect 106 -22783 112 -22207
rect 146 -22783 152 -22207
rect 106 -22795 152 -22783
rect -96 -22833 96 -22827
rect -96 -22867 -84 -22833
rect 84 -22867 96 -22833
rect -96 -22873 96 -22867
rect -96 -22941 96 -22935
rect -96 -22975 -84 -22941
rect 84 -22975 96 -22941
rect -96 -22981 96 -22975
rect -152 -23025 -106 -23013
rect -152 -23601 -146 -23025
rect -112 -23601 -106 -23025
rect -152 -23613 -106 -23601
rect 106 -23025 152 -23013
rect 106 -23601 112 -23025
rect 146 -23601 152 -23025
rect 106 -23613 152 -23601
rect -96 -23651 96 -23645
rect -96 -23685 -84 -23651
rect 84 -23685 96 -23651
rect -96 -23691 96 -23685
rect -96 -23759 96 -23753
rect -96 -23793 -84 -23759
rect 84 -23793 96 -23759
rect -96 -23799 96 -23793
rect -152 -23843 -106 -23831
rect -152 -24419 -146 -23843
rect -112 -24419 -106 -23843
rect -152 -24431 -106 -24419
rect 106 -23843 152 -23831
rect 106 -24419 112 -23843
rect 146 -24419 152 -23843
rect 106 -24431 152 -24419
rect -96 -24469 96 -24463
rect -96 -24503 -84 -24469
rect 84 -24503 96 -24469
rect -96 -24509 96 -24503
rect -96 -24577 96 -24571
rect -96 -24611 -84 -24577
rect 84 -24611 96 -24577
rect -96 -24617 96 -24611
rect -152 -24661 -106 -24649
rect -152 -25237 -146 -24661
rect -112 -25237 -106 -24661
rect -152 -25249 -106 -25237
rect 106 -24661 152 -24649
rect 106 -25237 112 -24661
rect 146 -25237 152 -24661
rect 106 -25249 152 -25237
rect -96 -25287 96 -25281
rect -96 -25321 -84 -25287
rect 84 -25321 96 -25287
rect -96 -25327 96 -25321
rect -96 -25395 96 -25389
rect -96 -25429 -84 -25395
rect 84 -25429 96 -25395
rect -96 -25435 96 -25429
rect -152 -25479 -106 -25467
rect -152 -26055 -146 -25479
rect -112 -26055 -106 -25479
rect -152 -26067 -106 -26055
rect 106 -25479 152 -25467
rect 106 -26055 112 -25479
rect 146 -26055 152 -25479
rect 106 -26067 152 -26055
rect -96 -26105 96 -26099
rect -96 -26139 -84 -26105
rect 84 -26139 96 -26105
rect -96 -26145 96 -26139
rect -96 -26213 96 -26207
rect -96 -26247 -84 -26213
rect 84 -26247 96 -26213
rect -96 -26253 96 -26247
rect -152 -26297 -106 -26285
rect -152 -26873 -146 -26297
rect -112 -26873 -106 -26297
rect -152 -26885 -106 -26873
rect 106 -26297 152 -26285
rect 106 -26873 112 -26297
rect 146 -26873 152 -26297
rect 106 -26885 152 -26873
rect -96 -26923 96 -26917
rect -96 -26957 -84 -26923
rect 84 -26957 96 -26923
rect -96 -26963 96 -26957
rect -96 -27031 96 -27025
rect -96 -27065 -84 -27031
rect 84 -27065 96 -27031
rect -96 -27071 96 -27065
rect -152 -27115 -106 -27103
rect -152 -27691 -146 -27115
rect -112 -27691 -106 -27115
rect -152 -27703 -106 -27691
rect 106 -27115 152 -27103
rect 106 -27691 112 -27115
rect 146 -27691 152 -27115
rect 106 -27703 152 -27691
rect -96 -27741 96 -27735
rect -96 -27775 -84 -27741
rect 84 -27775 96 -27741
rect -96 -27781 96 -27775
rect -96 -27849 96 -27843
rect -96 -27883 -84 -27849
rect 84 -27883 96 -27849
rect -96 -27889 96 -27883
rect -152 -27933 -106 -27921
rect -152 -28509 -146 -27933
rect -112 -28509 -106 -27933
rect -152 -28521 -106 -28509
rect 106 -27933 152 -27921
rect 106 -28509 112 -27933
rect 146 -28509 152 -27933
rect 106 -28521 152 -28509
rect -96 -28559 96 -28553
rect -96 -28593 -84 -28559
rect 84 -28593 96 -28559
rect -96 -28599 96 -28593
rect -96 -28667 96 -28661
rect -96 -28701 -84 -28667
rect 84 -28701 96 -28667
rect -96 -28707 96 -28701
rect -152 -28751 -106 -28739
rect -152 -29327 -146 -28751
rect -112 -29327 -106 -28751
rect -152 -29339 -106 -29327
rect 106 -28751 152 -28739
rect 106 -29327 112 -28751
rect 146 -29327 152 -28751
rect 106 -29339 152 -29327
rect -96 -29377 96 -29371
rect -96 -29411 -84 -29377
rect 84 -29411 96 -29377
rect -96 -29417 96 -29411
rect -96 -29485 96 -29479
rect -96 -29519 -84 -29485
rect 84 -29519 96 -29485
rect -96 -29525 96 -29519
rect -152 -29569 -106 -29557
rect -152 -30145 -146 -29569
rect -112 -30145 -106 -29569
rect -152 -30157 -106 -30145
rect 106 -29569 152 -29557
rect 106 -30145 112 -29569
rect 146 -30145 152 -29569
rect 106 -30157 152 -30145
rect -96 -30195 96 -30189
rect -96 -30229 -84 -30195
rect 84 -30229 96 -30195
rect -96 -30235 96 -30229
rect -96 -30303 96 -30297
rect -96 -30337 -84 -30303
rect 84 -30337 96 -30303
rect -96 -30343 96 -30337
rect -152 -30387 -106 -30375
rect -152 -30963 -146 -30387
rect -112 -30963 -106 -30387
rect -152 -30975 -106 -30963
rect 106 -30387 152 -30375
rect 106 -30963 112 -30387
rect 146 -30963 152 -30387
rect 106 -30975 152 -30963
rect -96 -31013 96 -31007
rect -96 -31047 -84 -31013
rect 84 -31047 96 -31013
rect -96 -31053 96 -31047
rect -96 -31121 96 -31115
rect -96 -31155 -84 -31121
rect 84 -31155 96 -31121
rect -96 -31161 96 -31155
rect -152 -31205 -106 -31193
rect -152 -31781 -146 -31205
rect -112 -31781 -106 -31205
rect -152 -31793 -106 -31781
rect 106 -31205 152 -31193
rect 106 -31781 112 -31205
rect 146 -31781 152 -31205
rect 106 -31793 152 -31781
rect -96 -31831 96 -31825
rect -96 -31865 -84 -31831
rect 84 -31865 96 -31831
rect -96 -31871 96 -31865
rect -96 -31939 96 -31933
rect -96 -31973 -84 -31939
rect 84 -31973 96 -31939
rect -96 -31979 96 -31973
rect -152 -32023 -106 -32011
rect -152 -32599 -146 -32023
rect -112 -32599 -106 -32023
rect -152 -32611 -106 -32599
rect 106 -32023 152 -32011
rect 106 -32599 112 -32023
rect 146 -32599 152 -32023
rect 106 -32611 152 -32599
rect -96 -32649 96 -32643
rect -96 -32683 -84 -32649
rect 84 -32683 96 -32649
rect -96 -32689 96 -32683
rect -96 -32757 96 -32751
rect -96 -32791 -84 -32757
rect 84 -32791 96 -32757
rect -96 -32797 96 -32791
rect -152 -32841 -106 -32829
rect -152 -33417 -146 -32841
rect -112 -33417 -106 -32841
rect -152 -33429 -106 -33417
rect 106 -32841 152 -32829
rect 106 -33417 112 -32841
rect 146 -33417 152 -32841
rect 106 -33429 152 -33417
rect -96 -33467 96 -33461
rect -96 -33501 -84 -33467
rect 84 -33501 96 -33467
rect -96 -33507 96 -33501
rect -96 -33575 96 -33569
rect -96 -33609 -84 -33575
rect 84 -33609 96 -33575
rect -96 -33615 96 -33609
rect -152 -33659 -106 -33647
rect -152 -34235 -146 -33659
rect -112 -34235 -106 -33659
rect -152 -34247 -106 -34235
rect 106 -33659 152 -33647
rect 106 -34235 112 -33659
rect 146 -34235 152 -33659
rect 106 -34247 152 -34235
rect -96 -34285 96 -34279
rect -96 -34319 -84 -34285
rect 84 -34319 96 -34285
rect -96 -34325 96 -34319
rect -96 -34393 96 -34387
rect -96 -34427 -84 -34393
rect 84 -34427 96 -34393
rect -96 -34433 96 -34427
rect -152 -34477 -106 -34465
rect -152 -35053 -146 -34477
rect -112 -35053 -106 -34477
rect -152 -35065 -106 -35053
rect 106 -34477 152 -34465
rect 106 -35053 112 -34477
rect 146 -35053 152 -34477
rect 106 -35065 152 -35053
rect -96 -35103 96 -35097
rect -96 -35137 -84 -35103
rect 84 -35137 96 -35103
rect -96 -35143 96 -35137
rect -96 -35211 96 -35205
rect -96 -35245 -84 -35211
rect 84 -35245 96 -35211
rect -96 -35251 96 -35245
rect -152 -35295 -106 -35283
rect -152 -35871 -146 -35295
rect -112 -35871 -106 -35295
rect -152 -35883 -106 -35871
rect 106 -35295 152 -35283
rect 106 -35871 112 -35295
rect 146 -35871 152 -35295
rect 106 -35883 152 -35871
rect -96 -35921 96 -35915
rect -96 -35955 -84 -35921
rect 84 -35955 96 -35921
rect -96 -35961 96 -35955
rect -96 -36029 96 -36023
rect -96 -36063 -84 -36029
rect 84 -36063 96 -36029
rect -96 -36069 96 -36063
rect -152 -36113 -106 -36101
rect -152 -36689 -146 -36113
rect -112 -36689 -106 -36113
rect -152 -36701 -106 -36689
rect 106 -36113 152 -36101
rect 106 -36689 112 -36113
rect 146 -36689 152 -36113
rect 106 -36701 152 -36689
rect -96 -36739 96 -36733
rect -96 -36773 -84 -36739
rect 84 -36773 96 -36739
rect -96 -36779 96 -36773
rect -96 -36847 96 -36841
rect -96 -36881 -84 -36847
rect 84 -36881 96 -36847
rect -96 -36887 96 -36881
rect -152 -36931 -106 -36919
rect -152 -37507 -146 -36931
rect -112 -37507 -106 -36931
rect -152 -37519 -106 -37507
rect 106 -36931 152 -36919
rect 106 -37507 112 -36931
rect 146 -37507 152 -36931
rect 106 -37519 152 -37507
rect -96 -37557 96 -37551
rect -96 -37591 -84 -37557
rect 84 -37591 96 -37557
rect -96 -37597 96 -37591
rect -96 -37665 96 -37659
rect -96 -37699 -84 -37665
rect 84 -37699 96 -37665
rect -96 -37705 96 -37699
rect -152 -37749 -106 -37737
rect -152 -38325 -146 -37749
rect -112 -38325 -106 -37749
rect -152 -38337 -106 -38325
rect 106 -37749 152 -37737
rect 106 -38325 112 -37749
rect 146 -38325 152 -37749
rect 106 -38337 152 -38325
rect -96 -38375 96 -38369
rect -96 -38409 -84 -38375
rect 84 -38409 96 -38375
rect -96 -38415 96 -38409
rect -96 -38483 96 -38477
rect -96 -38517 -84 -38483
rect 84 -38517 96 -38483
rect -96 -38523 96 -38517
rect -152 -38567 -106 -38555
rect -152 -39143 -146 -38567
rect -112 -39143 -106 -38567
rect -152 -39155 -106 -39143
rect 106 -38567 152 -38555
rect 106 -39143 112 -38567
rect 146 -39143 152 -38567
rect 106 -39155 152 -39143
rect -96 -39193 96 -39187
rect -96 -39227 -84 -39193
rect 84 -39227 96 -39193
rect -96 -39233 96 -39227
rect -96 -39301 96 -39295
rect -96 -39335 -84 -39301
rect 84 -39335 96 -39301
rect -96 -39341 96 -39335
rect -152 -39385 -106 -39373
rect -152 -39961 -146 -39385
rect -112 -39961 -106 -39385
rect -152 -39973 -106 -39961
rect 106 -39385 152 -39373
rect 106 -39961 112 -39385
rect 146 -39961 152 -39385
rect 106 -39973 152 -39961
rect -96 -40011 96 -40005
rect -96 -40045 -84 -40011
rect 84 -40045 96 -40011
rect -96 -40051 96 -40045
rect -96 -40119 96 -40113
rect -96 -40153 -84 -40119
rect 84 -40153 96 -40119
rect -96 -40159 96 -40153
rect -152 -40203 -106 -40191
rect -152 -40779 -146 -40203
rect -112 -40779 -106 -40203
rect -152 -40791 -106 -40779
rect 106 -40203 152 -40191
rect 106 -40779 112 -40203
rect 146 -40779 152 -40203
rect 106 -40791 152 -40779
rect -96 -40829 96 -40823
rect -96 -40863 -84 -40829
rect 84 -40863 96 -40829
rect -96 -40869 96 -40863
rect -96 -40937 96 -40931
rect -96 -40971 -84 -40937
rect 84 -40971 96 -40937
rect -96 -40977 96 -40971
rect -152 -41021 -106 -41009
rect -152 -41597 -146 -41021
rect -112 -41597 -106 -41021
rect -152 -41609 -106 -41597
rect 106 -41021 152 -41009
rect 106 -41597 112 -41021
rect 146 -41597 152 -41021
rect 106 -41609 152 -41597
rect -96 -41647 96 -41641
rect -96 -41681 -84 -41647
rect 84 -41681 96 -41647
rect -96 -41687 96 -41681
rect -96 -41755 96 -41749
rect -96 -41789 -84 -41755
rect 84 -41789 96 -41755
rect -96 -41795 96 -41789
rect -152 -41839 -106 -41827
rect -152 -42415 -146 -41839
rect -112 -42415 -106 -41839
rect -152 -42427 -106 -42415
rect 106 -41839 152 -41827
rect 106 -42415 112 -41839
rect 146 -42415 152 -41839
rect 106 -42427 152 -42415
rect -96 -42465 96 -42459
rect -96 -42499 -84 -42465
rect 84 -42499 96 -42465
rect -96 -42505 96 -42499
rect -96 -42573 96 -42567
rect -96 -42607 -84 -42573
rect 84 -42607 96 -42573
rect -96 -42613 96 -42607
rect -152 -42657 -106 -42645
rect -152 -43233 -146 -42657
rect -112 -43233 -106 -42657
rect -152 -43245 -106 -43233
rect 106 -42657 152 -42645
rect 106 -43233 112 -42657
rect 146 -43233 152 -42657
rect 106 -43245 152 -43233
rect -96 -43283 96 -43277
rect -96 -43317 -84 -43283
rect 84 -43317 96 -43283
rect -96 -43323 96 -43317
rect -96 -43391 96 -43385
rect -96 -43425 -84 -43391
rect 84 -43425 96 -43391
rect -96 -43431 96 -43425
rect -152 -43475 -106 -43463
rect -152 -44051 -146 -43475
rect -112 -44051 -106 -43475
rect -152 -44063 -106 -44051
rect 106 -43475 152 -43463
rect 106 -44051 112 -43475
rect 146 -44051 152 -43475
rect 106 -44063 152 -44051
rect -96 -44101 96 -44095
rect -96 -44135 -84 -44101
rect 84 -44135 96 -44101
rect -96 -44141 96 -44135
rect -96 -44209 96 -44203
rect -96 -44243 -84 -44209
rect 84 -44243 96 -44209
rect -96 -44249 96 -44243
rect -152 -44293 -106 -44281
rect -152 -44869 -146 -44293
rect -112 -44869 -106 -44293
rect -152 -44881 -106 -44869
rect 106 -44293 152 -44281
rect 106 -44869 112 -44293
rect 146 -44869 152 -44293
rect 106 -44881 152 -44869
rect -96 -44919 96 -44913
rect -96 -44953 -84 -44919
rect 84 -44953 96 -44919
rect -96 -44959 96 -44953
rect -96 -45027 96 -45021
rect -96 -45061 -84 -45027
rect 84 -45061 96 -45027
rect -96 -45067 96 -45061
rect -152 -45111 -106 -45099
rect -152 -45687 -146 -45111
rect -112 -45687 -106 -45111
rect -152 -45699 -106 -45687
rect 106 -45111 152 -45099
rect 106 -45687 112 -45111
rect 146 -45687 152 -45111
rect 106 -45699 152 -45687
rect -96 -45737 96 -45731
rect -96 -45771 -84 -45737
rect 84 -45771 96 -45737
rect -96 -45777 96 -45771
rect -96 -45845 96 -45839
rect -96 -45879 -84 -45845
rect 84 -45879 96 -45845
rect -96 -45885 96 -45879
rect -152 -45929 -106 -45917
rect -152 -46505 -146 -45929
rect -112 -46505 -106 -45929
rect -152 -46517 -106 -46505
rect 106 -45929 152 -45917
rect 106 -46505 112 -45929
rect 146 -46505 152 -45929
rect 106 -46517 152 -46505
rect -96 -46555 96 -46549
rect -96 -46589 -84 -46555
rect 84 -46589 96 -46555
rect -96 -46595 96 -46589
rect -96 -46663 96 -46657
rect -96 -46697 -84 -46663
rect 84 -46697 96 -46663
rect -96 -46703 96 -46697
rect -152 -46747 -106 -46735
rect -152 -47323 -146 -46747
rect -112 -47323 -106 -46747
rect -152 -47335 -106 -47323
rect 106 -46747 152 -46735
rect 106 -47323 112 -46747
rect 146 -47323 152 -46747
rect 106 -47335 152 -47323
rect -96 -47373 96 -47367
rect -96 -47407 -84 -47373
rect 84 -47407 96 -47373
rect -96 -47413 96 -47407
rect -96 -47481 96 -47475
rect -96 -47515 -84 -47481
rect 84 -47515 96 -47481
rect -96 -47521 96 -47515
rect -152 -47565 -106 -47553
rect -152 -48141 -146 -47565
rect -112 -48141 -106 -47565
rect -152 -48153 -106 -48141
rect 106 -47565 152 -47553
rect 106 -48141 112 -47565
rect 146 -48141 152 -47565
rect 106 -48153 152 -48141
rect -96 -48191 96 -48185
rect -96 -48225 -84 -48191
rect 84 -48225 96 -48191
rect -96 -48231 96 -48225
rect -96 -48299 96 -48293
rect -96 -48333 -84 -48299
rect 84 -48333 96 -48299
rect -96 -48339 96 -48333
rect -152 -48383 -106 -48371
rect -152 -48959 -146 -48383
rect -112 -48959 -106 -48383
rect -152 -48971 -106 -48959
rect 106 -48383 152 -48371
rect 106 -48959 112 -48383
rect 146 -48959 152 -48383
rect 106 -48971 152 -48959
rect -96 -49009 96 -49003
rect -96 -49043 -84 -49009
rect 84 -49043 96 -49009
rect -96 -49049 96 -49043
rect -96 -49117 96 -49111
rect -96 -49151 -84 -49117
rect 84 -49151 96 -49117
rect -96 -49157 96 -49151
rect -152 -49201 -106 -49189
rect -152 -49777 -146 -49201
rect -112 -49777 -106 -49201
rect -152 -49789 -106 -49777
rect 106 -49201 152 -49189
rect 106 -49777 112 -49201
rect 146 -49777 152 -49201
rect 106 -49789 152 -49777
rect -96 -49827 96 -49821
rect -96 -49861 -84 -49827
rect 84 -49861 96 -49827
rect -96 -49867 96 -49861
rect -96 -49935 96 -49929
rect -96 -49969 -84 -49935
rect 84 -49969 96 -49935
rect -96 -49975 96 -49969
rect -152 -50019 -106 -50007
rect -152 -50595 -146 -50019
rect -112 -50595 -106 -50019
rect -152 -50607 -106 -50595
rect 106 -50019 152 -50007
rect 106 -50595 112 -50019
rect 146 -50595 152 -50019
rect 106 -50607 152 -50595
rect -96 -50645 96 -50639
rect -96 -50679 -84 -50645
rect 84 -50679 96 -50645
rect -96 -50685 96 -50679
rect -96 -50753 96 -50747
rect -96 -50787 -84 -50753
rect 84 -50787 96 -50753
rect -96 -50793 96 -50787
rect -152 -50837 -106 -50825
rect -152 -51413 -146 -50837
rect -112 -51413 -106 -50837
rect -152 -51425 -106 -51413
rect 106 -50837 152 -50825
rect 106 -51413 112 -50837
rect 146 -51413 152 -50837
rect 106 -51425 152 -51413
rect -96 -51463 96 -51457
rect -96 -51497 -84 -51463
rect 84 -51497 96 -51463
rect -96 -51503 96 -51497
rect -96 -51571 96 -51565
rect -96 -51605 -84 -51571
rect 84 -51605 96 -51571
rect -96 -51611 96 -51605
rect -152 -51655 -106 -51643
rect -152 -52231 -146 -51655
rect -112 -52231 -106 -51655
rect -152 -52243 -106 -52231
rect 106 -51655 152 -51643
rect 106 -52231 112 -51655
rect 146 -52231 152 -51655
rect 106 -52243 152 -52231
rect -96 -52281 96 -52275
rect -96 -52315 -84 -52281
rect 84 -52315 96 -52281
rect -96 -52321 96 -52315
rect -96 -52389 96 -52383
rect -96 -52423 -84 -52389
rect 84 -52423 96 -52389
rect -96 -52429 96 -52423
rect -152 -52473 -106 -52461
rect -152 -53049 -146 -52473
rect -112 -53049 -106 -52473
rect -152 -53061 -106 -53049
rect 106 -52473 152 -52461
rect 106 -53049 112 -52473
rect 146 -53049 152 -52473
rect 106 -53061 152 -53049
rect -96 -53099 96 -53093
rect -96 -53133 -84 -53099
rect 84 -53133 96 -53099
rect -96 -53139 96 -53133
rect -96 -53207 96 -53201
rect -96 -53241 -84 -53207
rect 84 -53241 96 -53207
rect -96 -53247 96 -53241
rect -152 -53291 -106 -53279
rect -152 -53867 -146 -53291
rect -112 -53867 -106 -53291
rect -152 -53879 -106 -53867
rect 106 -53291 152 -53279
rect 106 -53867 112 -53291
rect 146 -53867 152 -53291
rect 106 -53879 152 -53867
rect -96 -53917 96 -53911
rect -96 -53951 -84 -53917
rect 84 -53951 96 -53917
rect -96 -53957 96 -53951
rect -96 -54025 96 -54019
rect -96 -54059 -84 -54025
rect 84 -54059 96 -54025
rect -96 -54065 96 -54059
rect -152 -54109 -106 -54097
rect -152 -54685 -146 -54109
rect -112 -54685 -106 -54109
rect -152 -54697 -106 -54685
rect 106 -54109 152 -54097
rect 106 -54685 112 -54109
rect 146 -54685 152 -54109
rect 106 -54697 152 -54685
rect -96 -54735 96 -54729
rect -96 -54769 -84 -54735
rect 84 -54769 96 -54735
rect -96 -54775 96 -54769
rect -96 -54843 96 -54837
rect -96 -54877 -84 -54843
rect 84 -54877 96 -54843
rect -96 -54883 96 -54877
rect -152 -54927 -106 -54915
rect -152 -55503 -146 -54927
rect -112 -55503 -106 -54927
rect -152 -55515 -106 -55503
rect 106 -54927 152 -54915
rect 106 -55503 112 -54927
rect 146 -55503 152 -54927
rect 106 -55515 152 -55503
rect -96 -55553 96 -55547
rect -96 -55587 -84 -55553
rect 84 -55587 96 -55553
rect -96 -55593 96 -55587
rect -96 -55661 96 -55655
rect -96 -55695 -84 -55661
rect 84 -55695 96 -55661
rect -96 -55701 96 -55695
rect -152 -55745 -106 -55733
rect -152 -56321 -146 -55745
rect -112 -56321 -106 -55745
rect -152 -56333 -106 -56321
rect 106 -55745 152 -55733
rect 106 -56321 112 -55745
rect 146 -56321 152 -55745
rect 106 -56333 152 -56321
rect -96 -56371 96 -56365
rect -96 -56405 -84 -56371
rect 84 -56405 96 -56371
rect -96 -56411 96 -56405
rect -96 -56479 96 -56473
rect -96 -56513 -84 -56479
rect 84 -56513 96 -56479
rect -96 -56519 96 -56513
rect -152 -56563 -106 -56551
rect -152 -57139 -146 -56563
rect -112 -57139 -106 -56563
rect -152 -57151 -106 -57139
rect 106 -56563 152 -56551
rect 106 -57139 112 -56563
rect 146 -57139 152 -56563
rect 106 -57151 152 -57139
rect -96 -57189 96 -57183
rect -96 -57223 -84 -57189
rect 84 -57223 96 -57189
rect -96 -57229 96 -57223
rect -96 -57297 96 -57291
rect -96 -57331 -84 -57297
rect 84 -57331 96 -57297
rect -96 -57337 96 -57331
rect -152 -57381 -106 -57369
rect -152 -57957 -146 -57381
rect -112 -57957 -106 -57381
rect -152 -57969 -106 -57957
rect 106 -57381 152 -57369
rect 106 -57957 112 -57381
rect 146 -57957 152 -57381
rect 106 -57969 152 -57957
rect -96 -58007 96 -58001
rect -96 -58041 -84 -58007
rect 84 -58041 96 -58007
rect -96 -58047 96 -58041
rect -96 -58115 96 -58109
rect -96 -58149 -84 -58115
rect 84 -58149 96 -58115
rect -96 -58155 96 -58149
rect -152 -58199 -106 -58187
rect -152 -58775 -146 -58199
rect -112 -58775 -106 -58199
rect -152 -58787 -106 -58775
rect 106 -58199 152 -58187
rect 106 -58775 112 -58199
rect 146 -58775 152 -58199
rect 106 -58787 152 -58775
rect -96 -58825 96 -58819
rect -96 -58859 -84 -58825
rect 84 -58859 96 -58825
rect -96 -58865 96 -58859
rect -96 -58933 96 -58927
rect -96 -58967 -84 -58933
rect 84 -58967 96 -58933
rect -96 -58973 96 -58967
rect -152 -59017 -106 -59005
rect -152 -59593 -146 -59017
rect -112 -59593 -106 -59017
rect -152 -59605 -106 -59593
rect 106 -59017 152 -59005
rect 106 -59593 112 -59017
rect 146 -59593 152 -59017
rect 106 -59605 152 -59593
rect -96 -59643 96 -59637
rect -96 -59677 -84 -59643
rect 84 -59677 96 -59643
rect -96 -59683 96 -59677
rect -96 -59751 96 -59745
rect -96 -59785 -84 -59751
rect 84 -59785 96 -59751
rect -96 -59791 96 -59785
rect -152 -59835 -106 -59823
rect -152 -60411 -146 -59835
rect -112 -60411 -106 -59835
rect -152 -60423 -106 -60411
rect 106 -59835 152 -59823
rect 106 -60411 112 -59835
rect 146 -60411 152 -59835
rect 106 -60423 152 -60411
rect -96 -60461 96 -60455
rect -96 -60495 -84 -60461
rect 84 -60495 96 -60461
rect -96 -60501 96 -60495
rect -96 -60569 96 -60563
rect -96 -60603 -84 -60569
rect 84 -60603 96 -60569
rect -96 -60609 96 -60603
rect -152 -60653 -106 -60641
rect -152 -61229 -146 -60653
rect -112 -61229 -106 -60653
rect -152 -61241 -106 -61229
rect 106 -60653 152 -60641
rect 106 -61229 112 -60653
rect 146 -61229 152 -60653
rect 106 -61241 152 -61229
rect -96 -61279 96 -61273
rect -96 -61313 -84 -61279
rect 84 -61313 96 -61279
rect -96 -61319 96 -61313
rect -96 -61387 96 -61381
rect -96 -61421 -84 -61387
rect 84 -61421 96 -61387
rect -96 -61427 96 -61421
rect -152 -61471 -106 -61459
rect -152 -62047 -146 -61471
rect -112 -62047 -106 -61471
rect -152 -62059 -106 -62047
rect 106 -61471 152 -61459
rect 106 -62047 112 -61471
rect 146 -62047 152 -61471
rect 106 -62059 152 -62047
rect -96 -62097 96 -62091
rect -96 -62131 -84 -62097
rect 84 -62131 96 -62097
rect -96 -62137 96 -62131
rect -96 -62205 96 -62199
rect -96 -62239 -84 -62205
rect 84 -62239 96 -62205
rect -96 -62245 96 -62239
rect -152 -62289 -106 -62277
rect -152 -62865 -146 -62289
rect -112 -62865 -106 -62289
rect -152 -62877 -106 -62865
rect 106 -62289 152 -62277
rect 106 -62865 112 -62289
rect 146 -62865 152 -62289
rect 106 -62877 152 -62865
rect -96 -62915 96 -62909
rect -96 -62949 -84 -62915
rect 84 -62949 96 -62915
rect -96 -62955 96 -62949
rect -96 -63023 96 -63017
rect -96 -63057 -84 -63023
rect 84 -63057 96 -63023
rect -96 -63063 96 -63057
rect -152 -63107 -106 -63095
rect -152 -63683 -146 -63107
rect -112 -63683 -106 -63107
rect -152 -63695 -106 -63683
rect 106 -63107 152 -63095
rect 106 -63683 112 -63107
rect 146 -63683 152 -63107
rect 106 -63695 152 -63683
rect -96 -63733 96 -63727
rect -96 -63767 -84 -63733
rect 84 -63767 96 -63733
rect -96 -63773 96 -63767
rect -96 -63841 96 -63835
rect -96 -63875 -84 -63841
rect 84 -63875 96 -63841
rect -96 -63881 96 -63875
rect -152 -63925 -106 -63913
rect -152 -64501 -146 -63925
rect -112 -64501 -106 -63925
rect -152 -64513 -106 -64501
rect 106 -63925 152 -63913
rect 106 -64501 112 -63925
rect 146 -64501 152 -63925
rect 106 -64513 152 -64501
rect -96 -64551 96 -64545
rect -96 -64585 -84 -64551
rect 84 -64585 96 -64551
rect -96 -64591 96 -64585
rect -96 -64659 96 -64653
rect -96 -64693 -84 -64659
rect 84 -64693 96 -64659
rect -96 -64699 96 -64693
rect -152 -64743 -106 -64731
rect -152 -65319 -146 -64743
rect -112 -65319 -106 -64743
rect -152 -65331 -106 -65319
rect 106 -64743 152 -64731
rect 106 -65319 112 -64743
rect 146 -65319 152 -64743
rect 106 -65331 152 -65319
rect -96 -65369 96 -65363
rect -96 -65403 -84 -65369
rect 84 -65403 96 -65369
rect -96 -65409 96 -65403
rect -96 -65477 96 -65471
rect -96 -65511 -84 -65477
rect 84 -65511 96 -65477
rect -96 -65517 96 -65511
rect -152 -65561 -106 -65549
rect -152 -66137 -146 -65561
rect -112 -66137 -106 -65561
rect -152 -66149 -106 -66137
rect 106 -65561 152 -65549
rect 106 -66137 112 -65561
rect 146 -66137 152 -65561
rect 106 -66149 152 -66137
rect -96 -66187 96 -66181
rect -96 -66221 -84 -66187
rect 84 -66221 96 -66187
rect -96 -66227 96 -66221
rect -96 -66295 96 -66289
rect -96 -66329 -84 -66295
rect 84 -66329 96 -66295
rect -96 -66335 96 -66329
rect -152 -66379 -106 -66367
rect -152 -66955 -146 -66379
rect -112 -66955 -106 -66379
rect -152 -66967 -106 -66955
rect 106 -66379 152 -66367
rect 106 -66955 112 -66379
rect 146 -66955 152 -66379
rect 106 -66967 152 -66955
rect -96 -67005 96 -66999
rect -96 -67039 -84 -67005
rect 84 -67039 96 -67005
rect -96 -67045 96 -67039
rect -96 -67113 96 -67107
rect -96 -67147 -84 -67113
rect 84 -67147 96 -67113
rect -96 -67153 96 -67147
rect -152 -67197 -106 -67185
rect -152 -67773 -146 -67197
rect -112 -67773 -106 -67197
rect -152 -67785 -106 -67773
rect 106 -67197 152 -67185
rect 106 -67773 112 -67197
rect 146 -67773 152 -67197
rect 106 -67785 152 -67773
rect -96 -67823 96 -67817
rect -96 -67857 -84 -67823
rect 84 -67857 96 -67823
rect -96 -67863 96 -67857
rect -96 -67931 96 -67925
rect -96 -67965 -84 -67931
rect 84 -67965 96 -67931
rect -96 -67971 96 -67965
rect -152 -68015 -106 -68003
rect -152 -68591 -146 -68015
rect -112 -68591 -106 -68015
rect -152 -68603 -106 -68591
rect 106 -68015 152 -68003
rect 106 -68591 112 -68015
rect 146 -68591 152 -68015
rect 106 -68603 152 -68591
rect -96 -68641 96 -68635
rect -96 -68675 -84 -68641
rect 84 -68675 96 -68641
rect -96 -68681 96 -68675
rect -96 -68749 96 -68743
rect -96 -68783 -84 -68749
rect 84 -68783 96 -68749
rect -96 -68789 96 -68783
rect -152 -68833 -106 -68821
rect -152 -69409 -146 -68833
rect -112 -69409 -106 -68833
rect -152 -69421 -106 -69409
rect 106 -68833 152 -68821
rect 106 -69409 112 -68833
rect 146 -69409 152 -68833
rect 106 -69421 152 -69409
rect -96 -69459 96 -69453
rect -96 -69493 -84 -69459
rect 84 -69493 96 -69459
rect -96 -69499 96 -69493
rect -96 -69567 96 -69561
rect -96 -69601 -84 -69567
rect 84 -69601 96 -69567
rect -96 -69607 96 -69601
rect -152 -69651 -106 -69639
rect -152 -70227 -146 -69651
rect -112 -70227 -106 -69651
rect -152 -70239 -106 -70227
rect 106 -69651 152 -69639
rect 106 -70227 112 -69651
rect 146 -70227 152 -69651
rect 106 -70239 152 -70227
rect -96 -70277 96 -70271
rect -96 -70311 -84 -70277
rect 84 -70311 96 -70277
rect -96 -70317 96 -70311
rect -96 -70385 96 -70379
rect -96 -70419 -84 -70385
rect 84 -70419 96 -70385
rect -96 -70425 96 -70419
rect -152 -70469 -106 -70457
rect -152 -71045 -146 -70469
rect -112 -71045 -106 -70469
rect -152 -71057 -106 -71045
rect 106 -70469 152 -70457
rect 106 -71045 112 -70469
rect 146 -71045 152 -70469
rect 106 -71057 152 -71045
rect -96 -71095 96 -71089
rect -96 -71129 -84 -71095
rect 84 -71129 96 -71095
rect -96 -71135 96 -71129
rect -96 -71203 96 -71197
rect -96 -71237 -84 -71203
rect 84 -71237 96 -71203
rect -96 -71243 96 -71237
rect -152 -71287 -106 -71275
rect -152 -71863 -146 -71287
rect -112 -71863 -106 -71287
rect -152 -71875 -106 -71863
rect 106 -71287 152 -71275
rect 106 -71863 112 -71287
rect 146 -71863 152 -71287
rect 106 -71875 152 -71863
rect -96 -71913 96 -71907
rect -96 -71947 -84 -71913
rect 84 -71947 96 -71913
rect -96 -71953 96 -71947
rect -96 -72021 96 -72015
rect -96 -72055 -84 -72021
rect 84 -72055 96 -72021
rect -96 -72061 96 -72055
rect -152 -72105 -106 -72093
rect -152 -72681 -146 -72105
rect -112 -72681 -106 -72105
rect -152 -72693 -106 -72681
rect 106 -72105 152 -72093
rect 106 -72681 112 -72105
rect 146 -72681 152 -72105
rect 106 -72693 152 -72681
rect -96 -72731 96 -72725
rect -96 -72765 -84 -72731
rect 84 -72765 96 -72731
rect -96 -72771 96 -72765
rect -96 -72839 96 -72833
rect -96 -72873 -84 -72839
rect 84 -72873 96 -72839
rect -96 -72879 96 -72873
rect -152 -72923 -106 -72911
rect -152 -73499 -146 -72923
rect -112 -73499 -106 -72923
rect -152 -73511 -106 -73499
rect 106 -72923 152 -72911
rect 106 -73499 112 -72923
rect 146 -73499 152 -72923
rect 106 -73511 152 -73499
rect -96 -73549 96 -73543
rect -96 -73583 -84 -73549
rect 84 -73583 96 -73549
rect -96 -73589 96 -73583
rect -96 -73657 96 -73651
rect -96 -73691 -84 -73657
rect 84 -73691 96 -73657
rect -96 -73697 96 -73691
rect -152 -73741 -106 -73729
rect -152 -74317 -146 -73741
rect -112 -74317 -106 -73741
rect -152 -74329 -106 -74317
rect 106 -73741 152 -73729
rect 106 -74317 112 -73741
rect 146 -74317 152 -73741
rect 106 -74329 152 -74317
rect -96 -74367 96 -74361
rect -96 -74401 -84 -74367
rect 84 -74401 96 -74367
rect -96 -74407 96 -74401
rect -96 -74475 96 -74469
rect -96 -74509 -84 -74475
rect 84 -74509 96 -74475
rect -96 -74515 96 -74509
rect -152 -74559 -106 -74547
rect -152 -75135 -146 -74559
rect -112 -75135 -106 -74559
rect -152 -75147 -106 -75135
rect 106 -74559 152 -74547
rect 106 -75135 112 -74559
rect 146 -75135 152 -74559
rect 106 -75147 152 -75135
rect -96 -75185 96 -75179
rect -96 -75219 -84 -75185
rect 84 -75219 96 -75185
rect -96 -75225 96 -75219
rect -96 -75293 96 -75287
rect -96 -75327 -84 -75293
rect 84 -75327 96 -75293
rect -96 -75333 96 -75327
rect -152 -75377 -106 -75365
rect -152 -75953 -146 -75377
rect -112 -75953 -106 -75377
rect -152 -75965 -106 -75953
rect 106 -75377 152 -75365
rect 106 -75953 112 -75377
rect 146 -75953 152 -75377
rect 106 -75965 152 -75953
rect -96 -76003 96 -75997
rect -96 -76037 -84 -76003
rect 84 -76037 96 -76003
rect -96 -76043 96 -76037
rect -96 -76111 96 -76105
rect -96 -76145 -84 -76111
rect 84 -76145 96 -76111
rect -96 -76151 96 -76145
rect -152 -76195 -106 -76183
rect -152 -76771 -146 -76195
rect -112 -76771 -106 -76195
rect -152 -76783 -106 -76771
rect 106 -76195 152 -76183
rect 106 -76771 112 -76195
rect 146 -76771 152 -76195
rect 106 -76783 152 -76771
rect -96 -76821 96 -76815
rect -96 -76855 -84 -76821
rect 84 -76855 96 -76821
rect -96 -76861 96 -76855
rect -96 -76929 96 -76923
rect -96 -76963 -84 -76929
rect 84 -76963 96 -76929
rect -96 -76969 96 -76963
rect -152 -77013 -106 -77001
rect -152 -77589 -146 -77013
rect -112 -77589 -106 -77013
rect -152 -77601 -106 -77589
rect 106 -77013 152 -77001
rect 106 -77589 112 -77013
rect 146 -77589 152 -77013
rect 106 -77601 152 -77589
rect -96 -77639 96 -77633
rect -96 -77673 -84 -77639
rect 84 -77673 96 -77639
rect -96 -77679 96 -77673
rect -96 -77747 96 -77741
rect -96 -77781 -84 -77747
rect 84 -77781 96 -77747
rect -96 -77787 96 -77781
rect -152 -77831 -106 -77819
rect -152 -78407 -146 -77831
rect -112 -78407 -106 -77831
rect -152 -78419 -106 -78407
rect 106 -77831 152 -77819
rect 106 -78407 112 -77831
rect 146 -78407 152 -77831
rect 106 -78419 152 -78407
rect -96 -78457 96 -78451
rect -96 -78491 -84 -78457
rect 84 -78491 96 -78457
rect -96 -78497 96 -78491
rect -96 -78565 96 -78559
rect -96 -78599 -84 -78565
rect 84 -78599 96 -78565
rect -96 -78605 96 -78599
rect -152 -78649 -106 -78637
rect -152 -79225 -146 -78649
rect -112 -79225 -106 -78649
rect -152 -79237 -106 -79225
rect 106 -78649 152 -78637
rect 106 -79225 112 -78649
rect 146 -79225 152 -78649
rect 106 -79237 152 -79225
rect -96 -79275 96 -79269
rect -96 -79309 -84 -79275
rect 84 -79309 96 -79275
rect -96 -79315 96 -79309
rect -96 -79383 96 -79377
rect -96 -79417 -84 -79383
rect 84 -79417 96 -79383
rect -96 -79423 96 -79417
rect -152 -79467 -106 -79455
rect -152 -80043 -146 -79467
rect -112 -80043 -106 -79467
rect -152 -80055 -106 -80043
rect 106 -79467 152 -79455
rect 106 -80043 112 -79467
rect 146 -80043 152 -79467
rect 106 -80055 152 -80043
rect -96 -80093 96 -80087
rect -96 -80127 -84 -80093
rect 84 -80127 96 -80093
rect -96 -80133 96 -80127
rect -96 -80201 96 -80195
rect -96 -80235 -84 -80201
rect 84 -80235 96 -80201
rect -96 -80241 96 -80235
rect -152 -80285 -106 -80273
rect -152 -80861 -146 -80285
rect -112 -80861 -106 -80285
rect -152 -80873 -106 -80861
rect 106 -80285 152 -80273
rect 106 -80861 112 -80285
rect 146 -80861 152 -80285
rect 106 -80873 152 -80861
rect -96 -80911 96 -80905
rect -96 -80945 -84 -80911
rect 84 -80945 96 -80911
rect -96 -80951 96 -80945
rect -96 -81019 96 -81013
rect -96 -81053 -84 -81019
rect 84 -81053 96 -81019
rect -96 -81059 96 -81053
rect -152 -81103 -106 -81091
rect -152 -81679 -146 -81103
rect -112 -81679 -106 -81103
rect -152 -81691 -106 -81679
rect 106 -81103 152 -81091
rect 106 -81679 112 -81103
rect 146 -81679 152 -81103
rect 106 -81691 152 -81679
rect -96 -81729 96 -81723
rect -96 -81763 -84 -81729
rect 84 -81763 96 -81729
rect -96 -81769 96 -81763
rect -96 -81837 96 -81831
rect -96 -81871 -84 -81837
rect 84 -81871 96 -81837
rect -96 -81877 96 -81871
rect -152 -81921 -106 -81909
rect -152 -82497 -146 -81921
rect -112 -82497 -106 -81921
rect -152 -82509 -106 -82497
rect 106 -81921 152 -81909
rect 106 -82497 112 -81921
rect 146 -82497 152 -81921
rect 106 -82509 152 -82497
rect -96 -82547 96 -82541
rect -96 -82581 -84 -82547
rect 84 -82581 96 -82547
rect -96 -82587 96 -82581
rect -96 -82655 96 -82649
rect -96 -82689 -84 -82655
rect 84 -82689 96 -82655
rect -96 -82695 96 -82689
rect -152 -82739 -106 -82727
rect -152 -83315 -146 -82739
rect -112 -83315 -106 -82739
rect -152 -83327 -106 -83315
rect 106 -82739 152 -82727
rect 106 -83315 112 -82739
rect 146 -83315 152 -82739
rect 106 -83327 152 -83315
rect -96 -83365 96 -83359
rect -96 -83399 -84 -83365
rect 84 -83399 96 -83365
rect -96 -83405 96 -83399
rect -96 -83473 96 -83467
rect -96 -83507 -84 -83473
rect 84 -83507 96 -83473
rect -96 -83513 96 -83507
rect -152 -83557 -106 -83545
rect -152 -84133 -146 -83557
rect -112 -84133 -106 -83557
rect -152 -84145 -106 -84133
rect 106 -83557 152 -83545
rect 106 -84133 112 -83557
rect 146 -84133 152 -83557
rect 106 -84145 152 -84133
rect -96 -84183 96 -84177
rect -96 -84217 -84 -84183
rect 84 -84217 96 -84183
rect -96 -84223 96 -84217
rect -96 -84291 96 -84285
rect -96 -84325 -84 -84291
rect 84 -84325 96 -84291
rect -96 -84331 96 -84325
rect -152 -84375 -106 -84363
rect -152 -84951 -146 -84375
rect -112 -84951 -106 -84375
rect -152 -84963 -106 -84951
rect 106 -84375 152 -84363
rect 106 -84951 112 -84375
rect 146 -84951 152 -84375
rect 106 -84963 152 -84951
rect -96 -85001 96 -84995
rect -96 -85035 -84 -85001
rect 84 -85035 96 -85001
rect -96 -85041 96 -85035
rect -96 -85109 96 -85103
rect -96 -85143 -84 -85109
rect 84 -85143 96 -85109
rect -96 -85149 96 -85143
rect -152 -85193 -106 -85181
rect -152 -85769 -146 -85193
rect -112 -85769 -106 -85193
rect -152 -85781 -106 -85769
rect 106 -85193 152 -85181
rect 106 -85769 112 -85193
rect 146 -85769 152 -85193
rect 106 -85781 152 -85769
rect -96 -85819 96 -85813
rect -96 -85853 -84 -85819
rect 84 -85853 96 -85819
rect -96 -85859 96 -85853
rect -96 -85927 96 -85921
rect -96 -85961 -84 -85927
rect 84 -85961 96 -85927
rect -96 -85967 96 -85961
rect -152 -86011 -106 -85999
rect -152 -86587 -146 -86011
rect -112 -86587 -106 -86011
rect -152 -86599 -106 -86587
rect 106 -86011 152 -85999
rect 106 -86587 112 -86011
rect 146 -86587 152 -86011
rect 106 -86599 152 -86587
rect -96 -86637 96 -86631
rect -96 -86671 -84 -86637
rect 84 -86671 96 -86637
rect -96 -86677 96 -86671
rect -96 -86745 96 -86739
rect -96 -86779 -84 -86745
rect 84 -86779 96 -86745
rect -96 -86785 96 -86779
rect -152 -86829 -106 -86817
rect -152 -87405 -146 -86829
rect -112 -87405 -106 -86829
rect -152 -87417 -106 -87405
rect 106 -86829 152 -86817
rect 106 -87405 112 -86829
rect 146 -87405 152 -86829
rect 106 -87417 152 -87405
rect -96 -87455 96 -87449
rect -96 -87489 -84 -87455
rect 84 -87489 96 -87455
rect -96 -87495 96 -87489
rect -96 -87563 96 -87557
rect -96 -87597 -84 -87563
rect 84 -87597 96 -87563
rect -96 -87603 96 -87597
rect -152 -87647 -106 -87635
rect -152 -88223 -146 -87647
rect -112 -88223 -106 -87647
rect -152 -88235 -106 -88223
rect 106 -87647 152 -87635
rect 106 -88223 112 -87647
rect 146 -88223 152 -87647
rect 106 -88235 152 -88223
rect -96 -88273 96 -88267
rect -96 -88307 -84 -88273
rect 84 -88307 96 -88273
rect -96 -88313 96 -88307
rect -96 -88381 96 -88375
rect -96 -88415 -84 -88381
rect 84 -88415 96 -88381
rect -96 -88421 96 -88415
rect -152 -88465 -106 -88453
rect -152 -89041 -146 -88465
rect -112 -89041 -106 -88465
rect -152 -89053 -106 -89041
rect 106 -88465 152 -88453
rect 106 -89041 112 -88465
rect 146 -89041 152 -88465
rect 106 -89053 152 -89041
rect -96 -89091 96 -89085
rect -96 -89125 -84 -89091
rect 84 -89125 96 -89091
rect -96 -89131 96 -89125
rect -96 -89199 96 -89193
rect -96 -89233 -84 -89199
rect 84 -89233 96 -89199
rect -96 -89239 96 -89233
rect -152 -89283 -106 -89271
rect -152 -89859 -146 -89283
rect -112 -89859 -106 -89283
rect -152 -89871 -106 -89859
rect 106 -89283 152 -89271
rect 106 -89859 112 -89283
rect 146 -89859 152 -89283
rect 106 -89871 152 -89859
rect -96 -89909 96 -89903
rect -96 -89943 -84 -89909
rect 84 -89943 96 -89909
rect -96 -89949 96 -89943
rect -96 -90017 96 -90011
rect -96 -90051 -84 -90017
rect 84 -90051 96 -90017
rect -96 -90057 96 -90051
rect -152 -90101 -106 -90089
rect -152 -90677 -146 -90101
rect -112 -90677 -106 -90101
rect -152 -90689 -106 -90677
rect 106 -90101 152 -90089
rect 106 -90677 112 -90101
rect 146 -90677 152 -90101
rect 106 -90689 152 -90677
rect -96 -90727 96 -90721
rect -96 -90761 -84 -90727
rect 84 -90761 96 -90727
rect -96 -90767 96 -90761
rect -96 -90835 96 -90829
rect -96 -90869 -84 -90835
rect 84 -90869 96 -90835
rect -96 -90875 96 -90869
rect -152 -90919 -106 -90907
rect -152 -91495 -146 -90919
rect -112 -91495 -106 -90919
rect -152 -91507 -106 -91495
rect 106 -90919 152 -90907
rect 106 -91495 112 -90919
rect 146 -91495 152 -90919
rect 106 -91507 152 -91495
rect -96 -91545 96 -91539
rect -96 -91579 -84 -91545
rect 84 -91579 96 -91545
rect -96 -91585 96 -91579
rect -96 -91653 96 -91647
rect -96 -91687 -84 -91653
rect 84 -91687 96 -91653
rect -96 -91693 96 -91687
rect -152 -91737 -106 -91725
rect -152 -92313 -146 -91737
rect -112 -92313 -106 -91737
rect -152 -92325 -106 -92313
rect 106 -91737 152 -91725
rect 106 -92313 112 -91737
rect 146 -92313 152 -91737
rect 106 -92325 152 -92313
rect -96 -92363 96 -92357
rect -96 -92397 -84 -92363
rect 84 -92397 96 -92363
rect -96 -92403 96 -92397
rect -96 -92471 96 -92465
rect -96 -92505 -84 -92471
rect 84 -92505 96 -92471
rect -96 -92511 96 -92505
rect -152 -92555 -106 -92543
rect -152 -93131 -146 -92555
rect -112 -93131 -106 -92555
rect -152 -93143 -106 -93131
rect 106 -92555 152 -92543
rect 106 -93131 112 -92555
rect 146 -93131 152 -92555
rect 106 -93143 152 -93131
rect -96 -93181 96 -93175
rect -96 -93215 -84 -93181
rect 84 -93215 96 -93181
rect -96 -93221 96 -93215
rect -96 -93289 96 -93283
rect -96 -93323 -84 -93289
rect 84 -93323 96 -93289
rect -96 -93329 96 -93323
rect -152 -93373 -106 -93361
rect -152 -93949 -146 -93373
rect -112 -93949 -106 -93373
rect -152 -93961 -106 -93949
rect 106 -93373 152 -93361
rect 106 -93949 112 -93373
rect 146 -93949 152 -93373
rect 106 -93961 152 -93949
rect -96 -93999 96 -93993
rect -96 -94033 -84 -93999
rect 84 -94033 96 -93999
rect -96 -94039 96 -94033
rect -96 -94107 96 -94101
rect -96 -94141 -84 -94107
rect 84 -94141 96 -94107
rect -96 -94147 96 -94141
rect -152 -94191 -106 -94179
rect -152 -94767 -146 -94191
rect -112 -94767 -106 -94191
rect -152 -94779 -106 -94767
rect 106 -94191 152 -94179
rect 106 -94767 112 -94191
rect 146 -94767 152 -94191
rect 106 -94779 152 -94767
rect -96 -94817 96 -94811
rect -96 -94851 -84 -94817
rect 84 -94851 96 -94817
rect -96 -94857 96 -94851
rect -96 -94925 96 -94919
rect -96 -94959 -84 -94925
rect 84 -94959 96 -94925
rect -96 -94965 96 -94959
rect -152 -95009 -106 -94997
rect -152 -95585 -146 -95009
rect -112 -95585 -106 -95009
rect -152 -95597 -106 -95585
rect 106 -95009 152 -94997
rect 106 -95585 112 -95009
rect 146 -95585 152 -95009
rect 106 -95597 152 -95585
rect -96 -95635 96 -95629
rect -96 -95669 -84 -95635
rect 84 -95669 96 -95635
rect -96 -95675 96 -95669
rect -96 -95743 96 -95737
rect -96 -95777 -84 -95743
rect 84 -95777 96 -95743
rect -96 -95783 96 -95777
rect -152 -95827 -106 -95815
rect -152 -96403 -146 -95827
rect -112 -96403 -106 -95827
rect -152 -96415 -106 -96403
rect 106 -95827 152 -95815
rect 106 -96403 112 -95827
rect 146 -96403 152 -95827
rect 106 -96415 152 -96403
rect -96 -96453 96 -96447
rect -96 -96487 -84 -96453
rect 84 -96487 96 -96453
rect -96 -96493 96 -96487
rect -96 -96561 96 -96555
rect -96 -96595 -84 -96561
rect 84 -96595 96 -96561
rect -96 -96601 96 -96595
rect -152 -96645 -106 -96633
rect -152 -97221 -146 -96645
rect -112 -97221 -106 -96645
rect -152 -97233 -106 -97221
rect 106 -96645 152 -96633
rect 106 -97221 112 -96645
rect 146 -97221 152 -96645
rect 106 -97233 152 -97221
rect -96 -97271 96 -97265
rect -96 -97305 -84 -97271
rect 84 -97305 96 -97271
rect -96 -97311 96 -97305
rect -96 -97379 96 -97373
rect -96 -97413 -84 -97379
rect 84 -97413 96 -97379
rect -96 -97419 96 -97413
rect -152 -97463 -106 -97451
rect -152 -98039 -146 -97463
rect -112 -98039 -106 -97463
rect -152 -98051 -106 -98039
rect 106 -97463 152 -97451
rect 106 -98039 112 -97463
rect 146 -98039 152 -97463
rect 106 -98051 152 -98039
rect -96 -98089 96 -98083
rect -96 -98123 -84 -98089
rect 84 -98123 96 -98089
rect -96 -98129 96 -98123
rect -96 -98197 96 -98191
rect -96 -98231 -84 -98197
rect 84 -98231 96 -98197
rect -96 -98237 96 -98231
rect -152 -98281 -106 -98269
rect -152 -98857 -146 -98281
rect -112 -98857 -106 -98281
rect -152 -98869 -106 -98857
rect 106 -98281 152 -98269
rect 106 -98857 112 -98281
rect 146 -98857 152 -98281
rect 106 -98869 152 -98857
rect -96 -98907 96 -98901
rect -96 -98941 -84 -98907
rect 84 -98941 96 -98907
rect -96 -98947 96 -98941
rect -96 -99015 96 -99009
rect -96 -99049 -84 -99015
rect 84 -99049 96 -99015
rect -96 -99055 96 -99049
rect -152 -99099 -106 -99087
rect -152 -99675 -146 -99099
rect -112 -99675 -106 -99099
rect -152 -99687 -106 -99675
rect 106 -99099 152 -99087
rect 106 -99675 112 -99099
rect 146 -99675 152 -99099
rect 106 -99687 152 -99675
rect -96 -99725 96 -99719
rect -96 -99759 -84 -99725
rect 84 -99759 96 -99725
rect -96 -99765 96 -99759
rect -96 -99833 96 -99827
rect -96 -99867 -84 -99833
rect 84 -99867 96 -99833
rect -96 -99873 96 -99867
rect -152 -99917 -106 -99905
rect -152 -100493 -146 -99917
rect -112 -100493 -106 -99917
rect -152 -100505 -106 -100493
rect 106 -99917 152 -99905
rect 106 -100493 112 -99917
rect 146 -100493 152 -99917
rect 106 -100505 152 -100493
rect -96 -100543 96 -100537
rect -96 -100577 -84 -100543
rect 84 -100577 96 -100543
rect -96 -100583 96 -100577
rect -96 -100651 96 -100645
rect -96 -100685 -84 -100651
rect 84 -100685 96 -100651
rect -96 -100691 96 -100685
rect -152 -100735 -106 -100723
rect -152 -101311 -146 -100735
rect -112 -101311 -106 -100735
rect -152 -101323 -106 -101311
rect 106 -100735 152 -100723
rect 106 -101311 112 -100735
rect 146 -101311 152 -100735
rect 106 -101323 152 -101311
rect -96 -101361 96 -101355
rect -96 -101395 -84 -101361
rect 84 -101395 96 -101361
rect -96 -101401 96 -101395
rect -96 -101469 96 -101463
rect -96 -101503 -84 -101469
rect 84 -101503 96 -101469
rect -96 -101509 96 -101503
rect -152 -101553 -106 -101541
rect -152 -102129 -146 -101553
rect -112 -102129 -106 -101553
rect -152 -102141 -106 -102129
rect 106 -101553 152 -101541
rect 106 -102129 112 -101553
rect 146 -102129 152 -101553
rect 106 -102141 152 -102129
rect -96 -102179 96 -102173
rect -96 -102213 -84 -102179
rect 84 -102213 96 -102179
rect -96 -102219 96 -102213
rect -96 -102287 96 -102281
rect -96 -102321 -84 -102287
rect 84 -102321 96 -102287
rect -96 -102327 96 -102321
rect -152 -102371 -106 -102359
rect -152 -102947 -146 -102371
rect -112 -102947 -106 -102371
rect -152 -102959 -106 -102947
rect 106 -102371 152 -102359
rect 106 -102947 112 -102371
rect 146 -102947 152 -102371
rect 106 -102959 152 -102947
rect -96 -102997 96 -102991
rect -96 -103031 -84 -102997
rect 84 -103031 96 -102997
rect -96 -103037 96 -103031
rect -96 -103105 96 -103099
rect -96 -103139 -84 -103105
rect 84 -103139 96 -103105
rect -96 -103145 96 -103139
rect -152 -103189 -106 -103177
rect -152 -103765 -146 -103189
rect -112 -103765 -106 -103189
rect -152 -103777 -106 -103765
rect 106 -103189 152 -103177
rect 106 -103765 112 -103189
rect 146 -103765 152 -103189
rect 106 -103777 152 -103765
rect -96 -103815 96 -103809
rect -96 -103849 -84 -103815
rect 84 -103849 96 -103815
rect -96 -103855 96 -103849
rect -96 -103923 96 -103917
rect -96 -103957 -84 -103923
rect 84 -103957 96 -103923
rect -96 -103963 96 -103957
rect -152 -104007 -106 -103995
rect -152 -104583 -146 -104007
rect -112 -104583 -106 -104007
rect -152 -104595 -106 -104583
rect 106 -104007 152 -103995
rect 106 -104583 112 -104007
rect 146 -104583 152 -104007
rect 106 -104595 152 -104583
rect -96 -104633 96 -104627
rect -96 -104667 -84 -104633
rect 84 -104667 96 -104633
rect -96 -104673 96 -104667
<< properties >>
string FIXED_BBOX -263 -104788 263 104788
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 1.0 m 256 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
