magic
tech sky130A
timestamp 1717401419
<< pwell >>
rect -164 -429 164 429
<< mvnmos >>
rect -50 -300 50 300
<< mvndiff >>
rect -79 294 -50 300
rect -79 -294 -73 294
rect -56 -294 -50 294
rect -79 -300 -50 -294
rect 50 294 79 300
rect 50 -294 56 294
rect 73 -294 79 294
rect 50 -300 79 -294
<< mvndiffc >>
rect -73 -294 -56 294
rect 56 -294 73 294
<< mvpsubdiff >>
rect -146 405 146 411
rect -146 388 -92 405
rect 92 388 146 405
rect -146 382 146 388
rect -146 357 -117 382
rect -146 -357 -140 357
rect -123 -357 -117 357
rect 117 357 146 382
rect -146 -382 -117 -357
rect 117 -357 123 357
rect 140 -357 146 357
rect 117 -382 146 -357
rect -146 -388 146 -382
rect -146 -405 -92 -388
rect 92 -405 146 -388
rect -146 -411 146 -405
<< mvpsubdiffcont >>
rect -92 388 92 405
rect -140 -357 -123 357
rect 123 -357 140 357
rect -92 -405 92 -388
<< poly >>
rect -50 336 50 344
rect -50 319 -42 336
rect 42 319 50 336
rect -50 300 50 319
rect -50 -319 50 -300
rect -50 -336 -42 -319
rect 42 -336 50 -319
rect -50 -344 50 -336
<< polycont >>
rect -42 319 42 336
rect -42 -336 42 -319
<< locali >>
rect -140 388 -92 405
rect 92 388 140 405
rect -140 357 -123 388
rect 123 357 140 388
rect -50 319 -42 336
rect 42 319 50 336
rect -73 294 -56 302
rect -73 -302 -56 -294
rect 56 294 73 302
rect 56 -302 73 -294
rect -50 -336 -42 -319
rect 42 -336 50 -319
rect -140 -388 -123 -357
rect 123 -388 140 -357
rect -140 -405 -92 -388
rect 92 -405 140 -388
<< viali >>
rect -42 319 42 336
rect -73 -294 -56 294
rect 56 -294 73 294
rect -42 -336 42 -319
<< metal1 >>
rect -48 336 48 339
rect -48 319 -42 336
rect 42 319 48 336
rect -48 316 48 319
rect -76 294 -53 300
rect -76 -294 -73 294
rect -56 -294 -53 294
rect -76 -300 -53 -294
rect 53 294 76 300
rect 53 -294 56 294
rect 73 -294 76 294
rect 53 -300 76 -294
rect -48 -319 48 -316
rect -48 -336 -42 -319
rect 42 -336 48 -319
rect -48 -339 48 -336
<< properties >>
string FIXED_BBOX -131 -396 131 396
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
