magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 10032 -2965 10148 -2899
rect 9884 -3232 9894 -3219
rect 9818 -3274 9894 -3232
rect 9946 -3274 10148 -3219
rect 9962 -3277 10148 -3274
rect 13228 -3232 13238 -3219
rect 13162 -3274 13238 -3232
rect 10076 -3393 10276 -3385
rect 10092 -3397 10260 -3393
rect 10018 -3574 10118 -3450
rect 13162 -3514 13306 -3274
rect 10018 -3628 10020 -3574
rect 13162 -3600 13336 -3514
rect 13362 -3574 13462 -3450
rect 13362 -3628 13364 -3574
rect 9703 -4371 9847 -4324
rect 9884 -4371 9901 -4270
rect 13047 -4371 13191 -4324
rect 13228 -4371 13245 -4270
rect 9703 -4382 9819 -4371
rect 9789 -4407 9819 -4382
rect 9801 -4906 9819 -4407
rect 13047 -4382 13819 -4371
rect 13133 -4407 13819 -4382
rect 13145 -4436 13819 -4407
rect 10983 -4848 11030 -4483
rect 11037 -4848 11084 -4537
rect 13145 -4848 13878 -4436
rect 14327 -4848 14374 -4483
rect 14381 -4848 14428 -4537
rect 10952 -4943 11155 -4848
rect 13145 -4906 14499 -4848
rect 12572 -4943 14499 -4906
rect 10952 -5067 11657 -4943
rect 12572 -5067 15001 -4943
rect 10952 -6152 11710 -5067
rect 12572 -6022 15054 -5067
rect 13163 -6087 15054 -6022
rect 13754 -6147 15054 -6087
rect 13783 -6152 15054 -6147
rect 10563 -6170 11710 -6152
rect 13907 -6170 15054 -6152
rect 11001 -6181 11710 -6170
rect 14345 -6181 15054 -6170
rect 11001 -6217 11675 -6181
rect 14345 -6217 15019 -6181
rect 11184 -6235 11675 -6217
rect 14528 -6235 15019 -6217
<< error_s >>
rect 3344 -2965 3460 -2899
rect 6688 -2965 6804 -2899
rect 3460 -3219 3846 -3153
rect 6804 -3219 7190 -3153
rect 3196 -3232 3206 -3219
rect 3130 -3274 3206 -3232
rect 3258 -3274 3846 -3219
rect 6540 -3232 6550 -3219
rect 3130 -3277 3846 -3274
rect 3130 -3514 3274 -3277
rect 3460 -3299 3846 -3277
rect 3384 -3385 3846 -3299
rect 6474 -3274 6550 -3232
rect 6602 -3274 7190 -3219
rect 6474 -3277 7190 -3274
rect 3388 -3393 3588 -3385
rect 3404 -3397 3572 -3393
rect 3130 -3600 3304 -3514
rect 3330 -3574 3430 -3450
rect 6474 -3514 6618 -3277
rect 6804 -3299 7190 -3277
rect 6728 -3385 7190 -3299
rect 6732 -3393 6932 -3385
rect 6748 -3397 6916 -3393
rect 3330 -3628 3332 -3574
rect 6474 -3600 6648 -3514
rect 6674 -3574 6774 -3450
rect 6674 -3628 6676 -3574
rect 3015 -4371 3159 -4324
rect 3196 -4371 3213 -4270
rect 6359 -4371 6503 -4324
rect 6540 -4371 6557 -4270
rect 3015 -4382 3787 -4371
rect 6359 -4382 7131 -4371
rect 3101 -4407 3787 -4382
rect 6445 -4407 7131 -4382
rect 3113 -4436 3787 -4407
rect 6457 -4436 7131 -4407
rect 3113 -4848 3846 -4436
rect 4295 -4848 4342 -4483
rect 4349 -4848 4396 -4537
rect 6457 -4848 7190 -4436
rect 7639 -4848 7686 -4483
rect 7693 -4848 7740 -4537
rect 3113 -4906 4467 -4848
rect 6457 -4906 7811 -4848
rect 2540 -4943 4467 -4906
rect 5884 -4943 7811 -4906
rect 2540 -5067 4969 -4943
rect 5884 -5067 8313 -4943
rect 2540 -6022 5022 -5067
rect 5884 -6022 8366 -5067
rect 9228 -6022 9692 -4906
rect 3131 -6087 5022 -6022
rect 6475 -6087 8366 -6022
rect 3722 -6147 5022 -6087
rect 7066 -6147 8366 -6087
rect 3751 -6152 5022 -6147
rect 7095 -6152 8366 -6147
rect 3875 -6170 5022 -6152
rect 7219 -6170 8366 -6152
rect 4313 -6181 5022 -6170
rect 7657 -6181 8366 -6170
rect 4313 -6217 4987 -6181
rect 7657 -6217 8331 -6181
rect 4496 -6235 4987 -6217
rect 7840 -6235 8331 -6217
<< error_ps >>
rect 9818 -3514 9962 -3274
rect 10148 -3299 10534 -3153
rect 10072 -3385 10534 -3299
rect 9818 -3600 9992 -3514
rect 9819 -4436 10475 -4371
rect 9819 -4848 10534 -4436
rect 9819 -4906 10952 -4848
rect 9692 -6022 10952 -4906
rect 9819 -6087 10952 -6022
rect 10410 -6147 10952 -6087
rect 10439 -6152 10952 -6147
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use icell2scs  x1
timestamp 1717439242
transform 1 0 0 0 1 0
box 0 -6337 8432 458
use icell2scs  x2
timestamp 1717439242
transform 1 0 6688 0 1 0
box 0 -6337 8432 458
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
