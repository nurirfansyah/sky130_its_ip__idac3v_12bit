magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 3344 -2965 3460 -2899
rect 6688 -2965 6804 -2899
rect 10032 -2965 10148 -2899
rect 13376 -2965 13492 -2899
rect 16720 -2965 16836 -2899
rect 20064 -2965 20180 -2899
rect 23408 -2965 23524 -2899
rect 30096 -2965 30212 -2899
rect 33440 -2965 33556 -2899
rect 36784 -2965 36900 -2899
rect 40128 -2965 40244 -2899
rect 43472 -2965 43588 -2899
rect 46816 -2965 46932 -2899
rect 50160 -2965 50276 -2899
rect 3460 -3219 3846 -3153
rect 6804 -3219 7190 -3153
rect 10148 -3219 10534 -3153
rect 13492 -3219 13878 -3153
rect 16836 -3219 17222 -3153
rect 20180 -3219 20566 -3153
rect 23524 -3219 23910 -3153
rect 3196 -3232 3206 -3219
rect 3130 -3274 3206 -3232
rect 3258 -3274 3846 -3219
rect 6540 -3232 6550 -3219
rect 3130 -3277 3846 -3274
rect 3130 -3514 3274 -3277
rect 3460 -3299 3846 -3277
rect 3384 -3385 3846 -3299
rect 6474 -3274 6550 -3232
rect 6602 -3274 7190 -3219
rect 9884 -3232 9894 -3219
rect 6474 -3277 7190 -3274
rect 3388 -3393 3588 -3385
rect 3404 -3397 3572 -3393
rect 3130 -3600 3304 -3514
rect 3330 -3574 3430 -3450
rect 6474 -3514 6618 -3277
rect 6804 -3299 7190 -3277
rect 6728 -3385 7190 -3299
rect 9818 -3274 9894 -3232
rect 9946 -3274 10534 -3219
rect 13228 -3232 13238 -3219
rect 9818 -3277 10534 -3274
rect 6732 -3393 6932 -3385
rect 6748 -3397 6916 -3393
rect 3330 -3628 3332 -3574
rect 6474 -3600 6648 -3514
rect 6674 -3574 6774 -3450
rect 9818 -3514 9962 -3277
rect 10148 -3299 10534 -3277
rect 10072 -3385 10534 -3299
rect 13162 -3274 13238 -3232
rect 13290 -3274 13878 -3219
rect 16572 -3232 16582 -3219
rect 13162 -3277 13878 -3274
rect 10076 -3393 10276 -3385
rect 10092 -3397 10260 -3393
rect 6674 -3628 6676 -3574
rect 9818 -3600 9992 -3514
rect 10018 -3574 10118 -3450
rect 13162 -3514 13306 -3277
rect 13492 -3299 13878 -3277
rect 13416 -3385 13878 -3299
rect 16506 -3274 16582 -3232
rect 16634 -3274 17222 -3219
rect 19916 -3232 19926 -3219
rect 16506 -3277 17222 -3274
rect 13420 -3393 13620 -3385
rect 13436 -3397 13604 -3393
rect 10018 -3628 10020 -3574
rect 13162 -3600 13336 -3514
rect 13362 -3574 13462 -3450
rect 16506 -3514 16650 -3277
rect 16836 -3299 17222 -3277
rect 16760 -3385 17222 -3299
rect 19850 -3274 19926 -3232
rect 19978 -3274 20566 -3219
rect 23260 -3232 23270 -3219
rect 19850 -3277 20566 -3274
rect 16764 -3393 16964 -3385
rect 16780 -3397 16948 -3393
rect 13362 -3628 13364 -3574
rect 16506 -3600 16680 -3514
rect 16706 -3574 16806 -3450
rect 19850 -3514 19994 -3277
rect 20180 -3299 20566 -3277
rect 20104 -3385 20566 -3299
rect 23194 -3274 23270 -3232
rect 23322 -3274 23910 -3219
rect 23194 -3277 23910 -3274
rect 20108 -3393 20308 -3385
rect 20124 -3397 20292 -3393
rect 16706 -3628 16708 -3574
rect 19850 -3600 20024 -3514
rect 20050 -3574 20150 -3450
rect 23194 -3514 23338 -3277
rect 23524 -3299 23910 -3277
rect 23448 -3385 23910 -3299
rect 29948 -3232 29958 -3219
rect 23452 -3393 23652 -3385
rect 23468 -3397 23636 -3393
rect 20050 -3628 20052 -3574
rect 23194 -3600 23368 -3514
rect 23394 -3574 23494 -3450
rect 29882 -3274 29958 -3232
rect 30010 -3274 30212 -3219
rect 23394 -3628 23396 -3574
rect 30026 -3277 30212 -3274
rect 33556 -3219 33942 -3153
rect 36900 -3219 37286 -3153
rect 40244 -3219 40630 -3153
rect 43588 -3219 43974 -3153
rect 46932 -3219 47318 -3153
rect 50276 -3219 50662 -3153
rect 33292 -3232 33302 -3219
rect 33226 -3274 33302 -3232
rect 33354 -3274 33942 -3219
rect 36636 -3232 36646 -3219
rect 33226 -3277 33942 -3274
rect 30140 -3393 30340 -3385
rect 30156 -3397 30324 -3393
rect 30082 -3574 30182 -3450
rect 33226 -3514 33370 -3277
rect 33556 -3299 33942 -3277
rect 33480 -3385 33942 -3299
rect 36570 -3274 36646 -3232
rect 36698 -3274 37286 -3219
rect 39980 -3232 39990 -3219
rect 36570 -3277 37286 -3274
rect 33484 -3393 33684 -3385
rect 33500 -3397 33668 -3393
rect 30082 -3628 30084 -3574
rect 33226 -3600 33400 -3514
rect 33426 -3574 33526 -3450
rect 36570 -3514 36714 -3277
rect 36900 -3299 37286 -3277
rect 36824 -3385 37286 -3299
rect 39914 -3274 39990 -3232
rect 40042 -3274 40630 -3219
rect 43324 -3232 43334 -3219
rect 39914 -3277 40630 -3274
rect 36828 -3393 37028 -3385
rect 36844 -3397 37012 -3393
rect 33426 -3628 33428 -3574
rect 36570 -3600 36744 -3514
rect 36770 -3574 36870 -3450
rect 39914 -3514 40058 -3277
rect 40244 -3299 40630 -3277
rect 40168 -3385 40630 -3299
rect 43258 -3274 43334 -3232
rect 43386 -3274 43974 -3219
rect 46668 -3232 46678 -3219
rect 43258 -3277 43974 -3274
rect 40172 -3393 40372 -3385
rect 40188 -3397 40356 -3393
rect 36770 -3628 36772 -3574
rect 39914 -3600 40088 -3514
rect 40114 -3574 40214 -3450
rect 43258 -3514 43402 -3277
rect 43588 -3299 43974 -3277
rect 43512 -3385 43974 -3299
rect 46602 -3274 46678 -3232
rect 46730 -3274 47318 -3219
rect 50012 -3232 50022 -3219
rect 46602 -3277 47318 -3274
rect 43516 -3393 43716 -3385
rect 43532 -3397 43700 -3393
rect 40114 -3628 40116 -3574
rect 43258 -3600 43432 -3514
rect 43458 -3574 43558 -3450
rect 46602 -3514 46746 -3277
rect 46932 -3299 47318 -3277
rect 46856 -3385 47318 -3299
rect 49946 -3274 50022 -3232
rect 50074 -3274 50662 -3219
rect 53356 -3232 53366 -3219
rect 49946 -3277 50662 -3274
rect 46860 -3393 47060 -3385
rect 46876 -3397 47044 -3393
rect 43458 -3628 43460 -3574
rect 46602 -3600 46776 -3514
rect 46802 -3574 46902 -3450
rect 49946 -3514 50090 -3277
rect 50276 -3299 50662 -3277
rect 50200 -3385 50662 -3299
rect 53290 -3274 53366 -3232
rect 50204 -3393 50404 -3385
rect 50220 -3397 50388 -3393
rect 46802 -3628 46804 -3574
rect 49946 -3600 50120 -3514
rect 50146 -3574 50246 -3450
rect 53290 -3514 53434 -3274
rect 50146 -3628 50148 -3574
rect 53290 -3600 53464 -3514
rect 53490 -3574 53590 -3450
rect 53490 -3628 53492 -3574
rect 3015 -4371 3159 -4324
rect 3196 -4371 3213 -4270
rect 6359 -4371 6503 -4324
rect 6540 -4371 6557 -4270
rect 9703 -4371 9847 -4324
rect 9884 -4371 9901 -4270
rect 13047 -4371 13191 -4324
rect 13228 -4371 13245 -4270
rect 16391 -4371 16535 -4324
rect 16572 -4371 16589 -4270
rect 19735 -4371 19879 -4324
rect 19916 -4371 19933 -4270
rect 23079 -4371 23223 -4324
rect 23260 -4371 23277 -4270
rect 29767 -4371 29911 -4324
rect 29948 -4371 29965 -4270
rect 33111 -4371 33255 -4324
rect 33292 -4371 33309 -4270
rect 36455 -4371 36599 -4324
rect 36636 -4371 36653 -4270
rect 39799 -4371 39943 -4324
rect 39980 -4371 39997 -4270
rect 43143 -4371 43287 -4324
rect 43324 -4371 43341 -4270
rect 46487 -4371 46631 -4324
rect 46668 -4371 46685 -4270
rect 49831 -4371 49975 -4324
rect 50012 -4371 50029 -4270
rect 53175 -4371 53319 -4324
rect 53356 -4371 53373 -4270
rect 3015 -4382 3787 -4371
rect 6359 -4382 7131 -4371
rect 9703 -4382 10475 -4371
rect 13047 -4382 13819 -4371
rect 16391 -4382 17163 -4371
rect 19735 -4382 20507 -4371
rect 23079 -4382 23851 -4371
rect 29767 -4382 29883 -4371
rect 3101 -4407 3787 -4382
rect 6445 -4407 7131 -4382
rect 9789 -4407 10475 -4382
rect 13133 -4407 13819 -4382
rect 16477 -4407 17163 -4382
rect 19821 -4407 20507 -4382
rect 23165 -4407 23851 -4382
rect 29853 -4407 29883 -4382
rect 3113 -4436 3787 -4407
rect 6457 -4436 7131 -4407
rect 9801 -4436 10475 -4407
rect 13145 -4436 13819 -4407
rect 16489 -4436 17163 -4407
rect 19833 -4436 20507 -4407
rect 23177 -4436 23851 -4407
rect 3113 -4848 3846 -4436
rect 4295 -4848 4342 -4483
rect 4349 -4848 4396 -4537
rect 6457 -4848 7190 -4436
rect 7639 -4848 7686 -4483
rect 7693 -4848 7740 -4537
rect 9801 -4848 10534 -4436
rect 10983 -4848 11030 -4483
rect 11037 -4848 11084 -4537
rect 13145 -4848 13878 -4436
rect 14327 -4848 14374 -4483
rect 14381 -4848 14428 -4537
rect 16489 -4848 17222 -4436
rect 17671 -4848 17718 -4483
rect 17725 -4848 17772 -4537
rect 19833 -4848 20566 -4436
rect 21015 -4848 21062 -4483
rect 21069 -4848 21116 -4537
rect 23177 -4848 23910 -4436
rect 24359 -4848 24406 -4483
rect 24413 -4848 24460 -4537
rect 3113 -4906 4467 -4848
rect 6457 -4906 7811 -4848
rect 9801 -4906 11155 -4848
rect 13145 -4906 14499 -4848
rect 16489 -4906 17843 -4848
rect 19833 -4906 21187 -4848
rect 23177 -4906 24232 -4848
rect 2720 -4943 4467 -4906
rect 5884 -4943 7811 -4906
rect 9228 -4943 11155 -4906
rect 12572 -4943 14499 -4906
rect 15916 -4943 17843 -4906
rect 19260 -4943 21187 -4906
rect 2720 -5067 4969 -4943
rect 5884 -5067 8313 -4943
rect 9228 -5067 11657 -4943
rect 12572 -5067 15001 -4943
rect 15916 -5067 18345 -4943
rect 19260 -5067 21689 -4943
rect 2720 -6022 5022 -5067
rect 5884 -6022 8366 -5067
rect 9228 -6022 11710 -5067
rect 12572 -6022 15054 -5067
rect 15916 -6022 18398 -5067
rect 19260 -6022 21742 -5067
rect 22604 -6022 24232 -4906
rect 29865 -4906 29883 -4407
rect 33111 -4382 33883 -4371
rect 36455 -4382 37227 -4371
rect 39799 -4382 40571 -4371
rect 43143 -4382 43915 -4371
rect 46487 -4382 47259 -4371
rect 49831 -4382 50603 -4371
rect 53175 -4382 53947 -4371
rect 33197 -4407 33883 -4382
rect 36541 -4407 37227 -4382
rect 39885 -4407 40571 -4382
rect 43229 -4407 43915 -4382
rect 46573 -4407 47259 -4382
rect 49917 -4407 50603 -4382
rect 53261 -4407 53947 -4382
rect 33209 -4436 33883 -4407
rect 36553 -4436 37227 -4407
rect 39897 -4436 40571 -4407
rect 43241 -4436 43915 -4407
rect 46585 -4436 47259 -4407
rect 49929 -4436 50603 -4407
rect 53273 -4436 53947 -4407
rect 31047 -4848 31094 -4483
rect 31101 -4848 31148 -4537
rect 33209 -4848 33942 -4436
rect 34391 -4848 34438 -4483
rect 34445 -4848 34492 -4537
rect 36553 -4848 37286 -4436
rect 37735 -4848 37782 -4483
rect 37789 -4848 37836 -4537
rect 39897 -4848 40630 -4436
rect 41079 -4848 41126 -4483
rect 41133 -4848 41180 -4537
rect 43241 -4848 43974 -4436
rect 44423 -4848 44470 -4483
rect 44477 -4848 44524 -4537
rect 46585 -4848 47318 -4436
rect 47767 -4848 47814 -4483
rect 47821 -4848 47868 -4537
rect 49929 -4848 50662 -4436
rect 51111 -4848 51158 -4483
rect 51165 -4848 51212 -4537
rect 53273 -4848 54006 -4436
rect 54455 -4848 54502 -4483
rect 54509 -4848 54556 -4537
rect 3131 -6087 5022 -6022
rect 6475 -6087 8366 -6022
rect 9819 -6087 11710 -6022
rect 13163 -6087 15054 -6022
rect 16507 -6087 18398 -6022
rect 19851 -6087 21742 -6022
rect 23195 -6087 24232 -6022
rect 3722 -6147 5022 -6087
rect 7066 -6147 8366 -6087
rect 10410 -6147 11710 -6087
rect 13754 -6147 15054 -6087
rect 17098 -6147 18398 -6087
rect 20442 -6147 21742 -6087
rect 23786 -6147 24232 -6087
rect 3751 -6152 5022 -6147
rect 7095 -6152 8366 -6147
rect 10439 -6152 11710 -6147
rect 13783 -6152 15054 -6147
rect 17127 -6152 18398 -6147
rect 20471 -6152 21742 -6147
rect 23815 -6152 24232 -6147
rect 3875 -6170 5022 -6152
rect 7219 -6170 8366 -6152
rect 10563 -6170 11710 -6152
rect 13907 -6170 15054 -6152
rect 17251 -6170 18398 -6152
rect 20595 -6170 21742 -6152
rect 23939 -6170 24377 -6152
rect 4313 -6181 5022 -6170
rect 7657 -6181 8366 -6170
rect 11001 -6181 11710 -6170
rect 14345 -6181 15054 -6170
rect 17689 -6181 18398 -6170
rect 21033 -6181 21742 -6170
rect 4313 -6217 4987 -6181
rect 7657 -6217 8331 -6181
rect 11001 -6217 11675 -6181
rect 14345 -6217 15019 -6181
rect 17689 -6217 18363 -6181
rect 21033 -6217 21707 -6181
rect 25033 -6181 25086 -5067
rect 31016 -4943 31219 -4848
rect 33209 -4906 34563 -4848
rect 36553 -4906 37907 -4848
rect 39897 -4906 41251 -4848
rect 43241 -4906 44595 -4848
rect 46585 -4906 47939 -4848
rect 49929 -4906 51283 -4848
rect 53273 -4906 54627 -4848
rect 32636 -4943 34563 -4906
rect 35980 -4943 37907 -4906
rect 39324 -4943 41251 -4906
rect 42668 -4943 44595 -4906
rect 46012 -4943 47939 -4906
rect 49356 -4943 51283 -4906
rect 52700 -4943 54627 -4906
rect 31016 -5067 31721 -4943
rect 32636 -5067 35065 -4943
rect 35980 -5067 38409 -4943
rect 39324 -5067 41753 -4943
rect 42668 -5067 45097 -4943
rect 46012 -5067 48441 -4943
rect 49356 -5067 51785 -4943
rect 52700 -5067 55129 -4943
rect 31016 -6152 31774 -5067
rect 32636 -6022 35118 -5067
rect 35980 -6022 38462 -5067
rect 39324 -6022 41806 -5067
rect 42668 -6022 45150 -5067
rect 46012 -6022 48494 -5067
rect 49356 -6022 51838 -5067
rect 52700 -6022 55182 -5067
rect 33227 -6087 35118 -6022
rect 36571 -6087 38462 -6022
rect 39915 -6087 41806 -6022
rect 43259 -6087 45150 -6022
rect 46603 -6087 48494 -6022
rect 49947 -6087 51838 -6022
rect 53291 -6087 55182 -6022
rect 33818 -6147 35118 -6087
rect 37162 -6147 38462 -6087
rect 40506 -6147 41806 -6087
rect 43850 -6147 45150 -6087
rect 47194 -6147 48494 -6087
rect 50538 -6147 51838 -6087
rect 53882 -6147 55182 -6087
rect 33847 -6152 35118 -6147
rect 37191 -6152 38462 -6147
rect 40535 -6152 41806 -6147
rect 43879 -6152 45150 -6147
rect 47223 -6152 48494 -6147
rect 50567 -6152 51838 -6147
rect 53911 -6152 55182 -6147
rect 30627 -6170 31774 -6152
rect 33971 -6170 35118 -6152
rect 37315 -6170 38462 -6152
rect 40659 -6170 41806 -6152
rect 44003 -6170 45150 -6152
rect 47347 -6170 48494 -6152
rect 50691 -6170 51838 -6152
rect 54035 -6170 55182 -6152
rect 31065 -6181 31774 -6170
rect 34409 -6181 35118 -6170
rect 37753 -6181 38462 -6170
rect 41097 -6181 41806 -6170
rect 44441 -6181 45150 -6170
rect 47785 -6181 48494 -6170
rect 51129 -6181 51838 -6170
rect 54473 -6181 55182 -6170
rect 25033 -6217 25051 -6181
rect 31065 -6217 31739 -6181
rect 34409 -6217 35083 -6181
rect 37753 -6217 38427 -6181
rect 41097 -6217 41771 -6181
rect 44441 -6217 45115 -6181
rect 47785 -6217 48459 -6181
rect 51129 -6217 51803 -6181
rect 54473 -6217 55147 -6181
rect 4496 -6235 4987 -6217
rect 7840 -6235 8331 -6217
rect 11184 -6235 11675 -6217
rect 14528 -6235 15019 -6217
rect 17872 -6235 18363 -6217
rect 21216 -6235 21707 -6217
rect 24560 -6235 25051 -6217
rect 31248 -6235 31739 -6217
rect 34592 -6235 35083 -6217
rect 37936 -6235 38427 -6217
rect 41280 -6235 41771 -6217
rect 44624 -6235 45115 -6217
rect 47968 -6235 48459 -6217
rect 51312 -6235 51803 -6217
rect 54656 -6235 55147 -6217
<< error_s >>
rect 26752 -2965 26868 -2899
rect 26868 -3219 27254 -3153
rect 26604 -3232 26614 -3219
rect 26538 -3274 26614 -3232
rect 26666 -3274 27254 -3219
rect 26538 -3277 27254 -3274
rect 26538 -3514 26682 -3277
rect 26868 -3299 27254 -3277
rect 26792 -3385 27254 -3299
rect 26796 -3393 26996 -3385
rect 26812 -3397 26980 -3393
rect 26538 -3600 26712 -3514
rect 26738 -3574 26838 -3450
rect 26738 -3628 26740 -3574
rect 26423 -4371 26567 -4324
rect 26604 -4371 26621 -4270
rect 26423 -4382 27195 -4371
rect 26509 -4407 27195 -4382
rect 26521 -4436 27195 -4407
rect 26521 -4848 27254 -4436
rect 27703 -4848 27750 -4483
rect 27757 -4848 27804 -4537
rect 26521 -4906 27875 -4848
rect 25948 -4943 27875 -4906
rect 25948 -5067 28377 -4943
rect 25948 -6022 28430 -5067
rect 29292 -6022 29756 -4906
rect 26539 -6087 28430 -6022
rect 27130 -6147 28430 -6087
rect 27159 -6152 28430 -6147
rect 27283 -6170 28430 -6152
rect 27721 -6181 28430 -6170
rect 27721 -6217 28395 -6181
rect 27904 -6235 28395 -6217
<< error_ps >>
rect 29882 -3514 30026 -3274
rect 30212 -3299 30598 -3153
rect 30136 -3385 30598 -3299
rect 29882 -3600 30056 -3514
rect 2540 -6022 2720 -4906
rect 24232 -4943 24531 -4848
rect 29883 -4436 30539 -4371
rect 29883 -4848 30598 -4436
rect 29883 -4906 31016 -4848
rect 24232 -6152 25033 -4943
rect 24377 -6217 25033 -6152
rect 29756 -6022 31016 -4906
rect 29883 -6087 31016 -6022
rect 30474 -6147 31016 -6087
rect 30503 -6152 31016 -6147
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use icell8scs  x1
timestamp 1717439242
transform 1 0 0 0 1 0
box 0 -6337 28496 458
use icell8scs  x2
timestamp 1717439242
transform 1 0 26752 0 1 0
box 0 -6337 28496 458
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
