magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< nwell >>
rect -358 -132787 358 132787
<< mvpmos >>
rect -100 131690 100 132490
rect -100 130654 100 131454
rect -100 129618 100 130418
rect -100 128582 100 129382
rect -100 127546 100 128346
rect -100 126510 100 127310
rect -100 125474 100 126274
rect -100 124438 100 125238
rect -100 123402 100 124202
rect -100 122366 100 123166
rect -100 121330 100 122130
rect -100 120294 100 121094
rect -100 119258 100 120058
rect -100 118222 100 119022
rect -100 117186 100 117986
rect -100 116150 100 116950
rect -100 115114 100 115914
rect -100 114078 100 114878
rect -100 113042 100 113842
rect -100 112006 100 112806
rect -100 110970 100 111770
rect -100 109934 100 110734
rect -100 108898 100 109698
rect -100 107862 100 108662
rect -100 106826 100 107626
rect -100 105790 100 106590
rect -100 104754 100 105554
rect -100 103718 100 104518
rect -100 102682 100 103482
rect -100 101646 100 102446
rect -100 100610 100 101410
rect -100 99574 100 100374
rect -100 98538 100 99338
rect -100 97502 100 98302
rect -100 96466 100 97266
rect -100 95430 100 96230
rect -100 94394 100 95194
rect -100 93358 100 94158
rect -100 92322 100 93122
rect -100 91286 100 92086
rect -100 90250 100 91050
rect -100 89214 100 90014
rect -100 88178 100 88978
rect -100 87142 100 87942
rect -100 86106 100 86906
rect -100 85070 100 85870
rect -100 84034 100 84834
rect -100 82998 100 83798
rect -100 81962 100 82762
rect -100 80926 100 81726
rect -100 79890 100 80690
rect -100 78854 100 79654
rect -100 77818 100 78618
rect -100 76782 100 77582
rect -100 75746 100 76546
rect -100 74710 100 75510
rect -100 73674 100 74474
rect -100 72638 100 73438
rect -100 71602 100 72402
rect -100 70566 100 71366
rect -100 69530 100 70330
rect -100 68494 100 69294
rect -100 67458 100 68258
rect -100 66422 100 67222
rect -100 65386 100 66186
rect -100 64350 100 65150
rect -100 63314 100 64114
rect -100 62278 100 63078
rect -100 61242 100 62042
rect -100 60206 100 61006
rect -100 59170 100 59970
rect -100 58134 100 58934
rect -100 57098 100 57898
rect -100 56062 100 56862
rect -100 55026 100 55826
rect -100 53990 100 54790
rect -100 52954 100 53754
rect -100 51918 100 52718
rect -100 50882 100 51682
rect -100 49846 100 50646
rect -100 48810 100 49610
rect -100 47774 100 48574
rect -100 46738 100 47538
rect -100 45702 100 46502
rect -100 44666 100 45466
rect -100 43630 100 44430
rect -100 42594 100 43394
rect -100 41558 100 42358
rect -100 40522 100 41322
rect -100 39486 100 40286
rect -100 38450 100 39250
rect -100 37414 100 38214
rect -100 36378 100 37178
rect -100 35342 100 36142
rect -100 34306 100 35106
rect -100 33270 100 34070
rect -100 32234 100 33034
rect -100 31198 100 31998
rect -100 30162 100 30962
rect -100 29126 100 29926
rect -100 28090 100 28890
rect -100 27054 100 27854
rect -100 26018 100 26818
rect -100 24982 100 25782
rect -100 23946 100 24746
rect -100 22910 100 23710
rect -100 21874 100 22674
rect -100 20838 100 21638
rect -100 19802 100 20602
rect -100 18766 100 19566
rect -100 17730 100 18530
rect -100 16694 100 17494
rect -100 15658 100 16458
rect -100 14622 100 15422
rect -100 13586 100 14386
rect -100 12550 100 13350
rect -100 11514 100 12314
rect -100 10478 100 11278
rect -100 9442 100 10242
rect -100 8406 100 9206
rect -100 7370 100 8170
rect -100 6334 100 7134
rect -100 5298 100 6098
rect -100 4262 100 5062
rect -100 3226 100 4026
rect -100 2190 100 2990
rect -100 1154 100 1954
rect -100 118 100 918
rect -100 -918 100 -118
rect -100 -1954 100 -1154
rect -100 -2990 100 -2190
rect -100 -4026 100 -3226
rect -100 -5062 100 -4262
rect -100 -6098 100 -5298
rect -100 -7134 100 -6334
rect -100 -8170 100 -7370
rect -100 -9206 100 -8406
rect -100 -10242 100 -9442
rect -100 -11278 100 -10478
rect -100 -12314 100 -11514
rect -100 -13350 100 -12550
rect -100 -14386 100 -13586
rect -100 -15422 100 -14622
rect -100 -16458 100 -15658
rect -100 -17494 100 -16694
rect -100 -18530 100 -17730
rect -100 -19566 100 -18766
rect -100 -20602 100 -19802
rect -100 -21638 100 -20838
rect -100 -22674 100 -21874
rect -100 -23710 100 -22910
rect -100 -24746 100 -23946
rect -100 -25782 100 -24982
rect -100 -26818 100 -26018
rect -100 -27854 100 -27054
rect -100 -28890 100 -28090
rect -100 -29926 100 -29126
rect -100 -30962 100 -30162
rect -100 -31998 100 -31198
rect -100 -33034 100 -32234
rect -100 -34070 100 -33270
rect -100 -35106 100 -34306
rect -100 -36142 100 -35342
rect -100 -37178 100 -36378
rect -100 -38214 100 -37414
rect -100 -39250 100 -38450
rect -100 -40286 100 -39486
rect -100 -41322 100 -40522
rect -100 -42358 100 -41558
rect -100 -43394 100 -42594
rect -100 -44430 100 -43630
rect -100 -45466 100 -44666
rect -100 -46502 100 -45702
rect -100 -47538 100 -46738
rect -100 -48574 100 -47774
rect -100 -49610 100 -48810
rect -100 -50646 100 -49846
rect -100 -51682 100 -50882
rect -100 -52718 100 -51918
rect -100 -53754 100 -52954
rect -100 -54790 100 -53990
rect -100 -55826 100 -55026
rect -100 -56862 100 -56062
rect -100 -57898 100 -57098
rect -100 -58934 100 -58134
rect -100 -59970 100 -59170
rect -100 -61006 100 -60206
rect -100 -62042 100 -61242
rect -100 -63078 100 -62278
rect -100 -64114 100 -63314
rect -100 -65150 100 -64350
rect -100 -66186 100 -65386
rect -100 -67222 100 -66422
rect -100 -68258 100 -67458
rect -100 -69294 100 -68494
rect -100 -70330 100 -69530
rect -100 -71366 100 -70566
rect -100 -72402 100 -71602
rect -100 -73438 100 -72638
rect -100 -74474 100 -73674
rect -100 -75510 100 -74710
rect -100 -76546 100 -75746
rect -100 -77582 100 -76782
rect -100 -78618 100 -77818
rect -100 -79654 100 -78854
rect -100 -80690 100 -79890
rect -100 -81726 100 -80926
rect -100 -82762 100 -81962
rect -100 -83798 100 -82998
rect -100 -84834 100 -84034
rect -100 -85870 100 -85070
rect -100 -86906 100 -86106
rect -100 -87942 100 -87142
rect -100 -88978 100 -88178
rect -100 -90014 100 -89214
rect -100 -91050 100 -90250
rect -100 -92086 100 -91286
rect -100 -93122 100 -92322
rect -100 -94158 100 -93358
rect -100 -95194 100 -94394
rect -100 -96230 100 -95430
rect -100 -97266 100 -96466
rect -100 -98302 100 -97502
rect -100 -99338 100 -98538
rect -100 -100374 100 -99574
rect -100 -101410 100 -100610
rect -100 -102446 100 -101646
rect -100 -103482 100 -102682
rect -100 -104518 100 -103718
rect -100 -105554 100 -104754
rect -100 -106590 100 -105790
rect -100 -107626 100 -106826
rect -100 -108662 100 -107862
rect -100 -109698 100 -108898
rect -100 -110734 100 -109934
rect -100 -111770 100 -110970
rect -100 -112806 100 -112006
rect -100 -113842 100 -113042
rect -100 -114878 100 -114078
rect -100 -115914 100 -115114
rect -100 -116950 100 -116150
rect -100 -117986 100 -117186
rect -100 -119022 100 -118222
rect -100 -120058 100 -119258
rect -100 -121094 100 -120294
rect -100 -122130 100 -121330
rect -100 -123166 100 -122366
rect -100 -124202 100 -123402
rect -100 -125238 100 -124438
rect -100 -126274 100 -125474
rect -100 -127310 100 -126510
rect -100 -128346 100 -127546
rect -100 -129382 100 -128582
rect -100 -130418 100 -129618
rect -100 -131454 100 -130654
rect -100 -132490 100 -131690
<< mvpdiff >>
rect -158 132478 -100 132490
rect -158 131702 -146 132478
rect -112 131702 -100 132478
rect -158 131690 -100 131702
rect 100 132478 158 132490
rect 100 131702 112 132478
rect 146 131702 158 132478
rect 100 131690 158 131702
rect -158 131442 -100 131454
rect -158 130666 -146 131442
rect -112 130666 -100 131442
rect -158 130654 -100 130666
rect 100 131442 158 131454
rect 100 130666 112 131442
rect 146 130666 158 131442
rect 100 130654 158 130666
rect -158 130406 -100 130418
rect -158 129630 -146 130406
rect -112 129630 -100 130406
rect -158 129618 -100 129630
rect 100 130406 158 130418
rect 100 129630 112 130406
rect 146 129630 158 130406
rect 100 129618 158 129630
rect -158 129370 -100 129382
rect -158 128594 -146 129370
rect -112 128594 -100 129370
rect -158 128582 -100 128594
rect 100 129370 158 129382
rect 100 128594 112 129370
rect 146 128594 158 129370
rect 100 128582 158 128594
rect -158 128334 -100 128346
rect -158 127558 -146 128334
rect -112 127558 -100 128334
rect -158 127546 -100 127558
rect 100 128334 158 128346
rect 100 127558 112 128334
rect 146 127558 158 128334
rect 100 127546 158 127558
rect -158 127298 -100 127310
rect -158 126522 -146 127298
rect -112 126522 -100 127298
rect -158 126510 -100 126522
rect 100 127298 158 127310
rect 100 126522 112 127298
rect 146 126522 158 127298
rect 100 126510 158 126522
rect -158 126262 -100 126274
rect -158 125486 -146 126262
rect -112 125486 -100 126262
rect -158 125474 -100 125486
rect 100 126262 158 126274
rect 100 125486 112 126262
rect 146 125486 158 126262
rect 100 125474 158 125486
rect -158 125226 -100 125238
rect -158 124450 -146 125226
rect -112 124450 -100 125226
rect -158 124438 -100 124450
rect 100 125226 158 125238
rect 100 124450 112 125226
rect 146 124450 158 125226
rect 100 124438 158 124450
rect -158 124190 -100 124202
rect -158 123414 -146 124190
rect -112 123414 -100 124190
rect -158 123402 -100 123414
rect 100 124190 158 124202
rect 100 123414 112 124190
rect 146 123414 158 124190
rect 100 123402 158 123414
rect -158 123154 -100 123166
rect -158 122378 -146 123154
rect -112 122378 -100 123154
rect -158 122366 -100 122378
rect 100 123154 158 123166
rect 100 122378 112 123154
rect 146 122378 158 123154
rect 100 122366 158 122378
rect -158 122118 -100 122130
rect -158 121342 -146 122118
rect -112 121342 -100 122118
rect -158 121330 -100 121342
rect 100 122118 158 122130
rect 100 121342 112 122118
rect 146 121342 158 122118
rect 100 121330 158 121342
rect -158 121082 -100 121094
rect -158 120306 -146 121082
rect -112 120306 -100 121082
rect -158 120294 -100 120306
rect 100 121082 158 121094
rect 100 120306 112 121082
rect 146 120306 158 121082
rect 100 120294 158 120306
rect -158 120046 -100 120058
rect -158 119270 -146 120046
rect -112 119270 -100 120046
rect -158 119258 -100 119270
rect 100 120046 158 120058
rect 100 119270 112 120046
rect 146 119270 158 120046
rect 100 119258 158 119270
rect -158 119010 -100 119022
rect -158 118234 -146 119010
rect -112 118234 -100 119010
rect -158 118222 -100 118234
rect 100 119010 158 119022
rect 100 118234 112 119010
rect 146 118234 158 119010
rect 100 118222 158 118234
rect -158 117974 -100 117986
rect -158 117198 -146 117974
rect -112 117198 -100 117974
rect -158 117186 -100 117198
rect 100 117974 158 117986
rect 100 117198 112 117974
rect 146 117198 158 117974
rect 100 117186 158 117198
rect -158 116938 -100 116950
rect -158 116162 -146 116938
rect -112 116162 -100 116938
rect -158 116150 -100 116162
rect 100 116938 158 116950
rect 100 116162 112 116938
rect 146 116162 158 116938
rect 100 116150 158 116162
rect -158 115902 -100 115914
rect -158 115126 -146 115902
rect -112 115126 -100 115902
rect -158 115114 -100 115126
rect 100 115902 158 115914
rect 100 115126 112 115902
rect 146 115126 158 115902
rect 100 115114 158 115126
rect -158 114866 -100 114878
rect -158 114090 -146 114866
rect -112 114090 -100 114866
rect -158 114078 -100 114090
rect 100 114866 158 114878
rect 100 114090 112 114866
rect 146 114090 158 114866
rect 100 114078 158 114090
rect -158 113830 -100 113842
rect -158 113054 -146 113830
rect -112 113054 -100 113830
rect -158 113042 -100 113054
rect 100 113830 158 113842
rect 100 113054 112 113830
rect 146 113054 158 113830
rect 100 113042 158 113054
rect -158 112794 -100 112806
rect -158 112018 -146 112794
rect -112 112018 -100 112794
rect -158 112006 -100 112018
rect 100 112794 158 112806
rect 100 112018 112 112794
rect 146 112018 158 112794
rect 100 112006 158 112018
rect -158 111758 -100 111770
rect -158 110982 -146 111758
rect -112 110982 -100 111758
rect -158 110970 -100 110982
rect 100 111758 158 111770
rect 100 110982 112 111758
rect 146 110982 158 111758
rect 100 110970 158 110982
rect -158 110722 -100 110734
rect -158 109946 -146 110722
rect -112 109946 -100 110722
rect -158 109934 -100 109946
rect 100 110722 158 110734
rect 100 109946 112 110722
rect 146 109946 158 110722
rect 100 109934 158 109946
rect -158 109686 -100 109698
rect -158 108910 -146 109686
rect -112 108910 -100 109686
rect -158 108898 -100 108910
rect 100 109686 158 109698
rect 100 108910 112 109686
rect 146 108910 158 109686
rect 100 108898 158 108910
rect -158 108650 -100 108662
rect -158 107874 -146 108650
rect -112 107874 -100 108650
rect -158 107862 -100 107874
rect 100 108650 158 108662
rect 100 107874 112 108650
rect 146 107874 158 108650
rect 100 107862 158 107874
rect -158 107614 -100 107626
rect -158 106838 -146 107614
rect -112 106838 -100 107614
rect -158 106826 -100 106838
rect 100 107614 158 107626
rect 100 106838 112 107614
rect 146 106838 158 107614
rect 100 106826 158 106838
rect -158 106578 -100 106590
rect -158 105802 -146 106578
rect -112 105802 -100 106578
rect -158 105790 -100 105802
rect 100 106578 158 106590
rect 100 105802 112 106578
rect 146 105802 158 106578
rect 100 105790 158 105802
rect -158 105542 -100 105554
rect -158 104766 -146 105542
rect -112 104766 -100 105542
rect -158 104754 -100 104766
rect 100 105542 158 105554
rect 100 104766 112 105542
rect 146 104766 158 105542
rect 100 104754 158 104766
rect -158 104506 -100 104518
rect -158 103730 -146 104506
rect -112 103730 -100 104506
rect -158 103718 -100 103730
rect 100 104506 158 104518
rect 100 103730 112 104506
rect 146 103730 158 104506
rect 100 103718 158 103730
rect -158 103470 -100 103482
rect -158 102694 -146 103470
rect -112 102694 -100 103470
rect -158 102682 -100 102694
rect 100 103470 158 103482
rect 100 102694 112 103470
rect 146 102694 158 103470
rect 100 102682 158 102694
rect -158 102434 -100 102446
rect -158 101658 -146 102434
rect -112 101658 -100 102434
rect -158 101646 -100 101658
rect 100 102434 158 102446
rect 100 101658 112 102434
rect 146 101658 158 102434
rect 100 101646 158 101658
rect -158 101398 -100 101410
rect -158 100622 -146 101398
rect -112 100622 -100 101398
rect -158 100610 -100 100622
rect 100 101398 158 101410
rect 100 100622 112 101398
rect 146 100622 158 101398
rect 100 100610 158 100622
rect -158 100362 -100 100374
rect -158 99586 -146 100362
rect -112 99586 -100 100362
rect -158 99574 -100 99586
rect 100 100362 158 100374
rect 100 99586 112 100362
rect 146 99586 158 100362
rect 100 99574 158 99586
rect -158 99326 -100 99338
rect -158 98550 -146 99326
rect -112 98550 -100 99326
rect -158 98538 -100 98550
rect 100 99326 158 99338
rect 100 98550 112 99326
rect 146 98550 158 99326
rect 100 98538 158 98550
rect -158 98290 -100 98302
rect -158 97514 -146 98290
rect -112 97514 -100 98290
rect -158 97502 -100 97514
rect 100 98290 158 98302
rect 100 97514 112 98290
rect 146 97514 158 98290
rect 100 97502 158 97514
rect -158 97254 -100 97266
rect -158 96478 -146 97254
rect -112 96478 -100 97254
rect -158 96466 -100 96478
rect 100 97254 158 97266
rect 100 96478 112 97254
rect 146 96478 158 97254
rect 100 96466 158 96478
rect -158 96218 -100 96230
rect -158 95442 -146 96218
rect -112 95442 -100 96218
rect -158 95430 -100 95442
rect 100 96218 158 96230
rect 100 95442 112 96218
rect 146 95442 158 96218
rect 100 95430 158 95442
rect -158 95182 -100 95194
rect -158 94406 -146 95182
rect -112 94406 -100 95182
rect -158 94394 -100 94406
rect 100 95182 158 95194
rect 100 94406 112 95182
rect 146 94406 158 95182
rect 100 94394 158 94406
rect -158 94146 -100 94158
rect -158 93370 -146 94146
rect -112 93370 -100 94146
rect -158 93358 -100 93370
rect 100 94146 158 94158
rect 100 93370 112 94146
rect 146 93370 158 94146
rect 100 93358 158 93370
rect -158 93110 -100 93122
rect -158 92334 -146 93110
rect -112 92334 -100 93110
rect -158 92322 -100 92334
rect 100 93110 158 93122
rect 100 92334 112 93110
rect 146 92334 158 93110
rect 100 92322 158 92334
rect -158 92074 -100 92086
rect -158 91298 -146 92074
rect -112 91298 -100 92074
rect -158 91286 -100 91298
rect 100 92074 158 92086
rect 100 91298 112 92074
rect 146 91298 158 92074
rect 100 91286 158 91298
rect -158 91038 -100 91050
rect -158 90262 -146 91038
rect -112 90262 -100 91038
rect -158 90250 -100 90262
rect 100 91038 158 91050
rect 100 90262 112 91038
rect 146 90262 158 91038
rect 100 90250 158 90262
rect -158 90002 -100 90014
rect -158 89226 -146 90002
rect -112 89226 -100 90002
rect -158 89214 -100 89226
rect 100 90002 158 90014
rect 100 89226 112 90002
rect 146 89226 158 90002
rect 100 89214 158 89226
rect -158 88966 -100 88978
rect -158 88190 -146 88966
rect -112 88190 -100 88966
rect -158 88178 -100 88190
rect 100 88966 158 88978
rect 100 88190 112 88966
rect 146 88190 158 88966
rect 100 88178 158 88190
rect -158 87930 -100 87942
rect -158 87154 -146 87930
rect -112 87154 -100 87930
rect -158 87142 -100 87154
rect 100 87930 158 87942
rect 100 87154 112 87930
rect 146 87154 158 87930
rect 100 87142 158 87154
rect -158 86894 -100 86906
rect -158 86118 -146 86894
rect -112 86118 -100 86894
rect -158 86106 -100 86118
rect 100 86894 158 86906
rect 100 86118 112 86894
rect 146 86118 158 86894
rect 100 86106 158 86118
rect -158 85858 -100 85870
rect -158 85082 -146 85858
rect -112 85082 -100 85858
rect -158 85070 -100 85082
rect 100 85858 158 85870
rect 100 85082 112 85858
rect 146 85082 158 85858
rect 100 85070 158 85082
rect -158 84822 -100 84834
rect -158 84046 -146 84822
rect -112 84046 -100 84822
rect -158 84034 -100 84046
rect 100 84822 158 84834
rect 100 84046 112 84822
rect 146 84046 158 84822
rect 100 84034 158 84046
rect -158 83786 -100 83798
rect -158 83010 -146 83786
rect -112 83010 -100 83786
rect -158 82998 -100 83010
rect 100 83786 158 83798
rect 100 83010 112 83786
rect 146 83010 158 83786
rect 100 82998 158 83010
rect -158 82750 -100 82762
rect -158 81974 -146 82750
rect -112 81974 -100 82750
rect -158 81962 -100 81974
rect 100 82750 158 82762
rect 100 81974 112 82750
rect 146 81974 158 82750
rect 100 81962 158 81974
rect -158 81714 -100 81726
rect -158 80938 -146 81714
rect -112 80938 -100 81714
rect -158 80926 -100 80938
rect 100 81714 158 81726
rect 100 80938 112 81714
rect 146 80938 158 81714
rect 100 80926 158 80938
rect -158 80678 -100 80690
rect -158 79902 -146 80678
rect -112 79902 -100 80678
rect -158 79890 -100 79902
rect 100 80678 158 80690
rect 100 79902 112 80678
rect 146 79902 158 80678
rect 100 79890 158 79902
rect -158 79642 -100 79654
rect -158 78866 -146 79642
rect -112 78866 -100 79642
rect -158 78854 -100 78866
rect 100 79642 158 79654
rect 100 78866 112 79642
rect 146 78866 158 79642
rect 100 78854 158 78866
rect -158 78606 -100 78618
rect -158 77830 -146 78606
rect -112 77830 -100 78606
rect -158 77818 -100 77830
rect 100 78606 158 78618
rect 100 77830 112 78606
rect 146 77830 158 78606
rect 100 77818 158 77830
rect -158 77570 -100 77582
rect -158 76794 -146 77570
rect -112 76794 -100 77570
rect -158 76782 -100 76794
rect 100 77570 158 77582
rect 100 76794 112 77570
rect 146 76794 158 77570
rect 100 76782 158 76794
rect -158 76534 -100 76546
rect -158 75758 -146 76534
rect -112 75758 -100 76534
rect -158 75746 -100 75758
rect 100 76534 158 76546
rect 100 75758 112 76534
rect 146 75758 158 76534
rect 100 75746 158 75758
rect -158 75498 -100 75510
rect -158 74722 -146 75498
rect -112 74722 -100 75498
rect -158 74710 -100 74722
rect 100 75498 158 75510
rect 100 74722 112 75498
rect 146 74722 158 75498
rect 100 74710 158 74722
rect -158 74462 -100 74474
rect -158 73686 -146 74462
rect -112 73686 -100 74462
rect -158 73674 -100 73686
rect 100 74462 158 74474
rect 100 73686 112 74462
rect 146 73686 158 74462
rect 100 73674 158 73686
rect -158 73426 -100 73438
rect -158 72650 -146 73426
rect -112 72650 -100 73426
rect -158 72638 -100 72650
rect 100 73426 158 73438
rect 100 72650 112 73426
rect 146 72650 158 73426
rect 100 72638 158 72650
rect -158 72390 -100 72402
rect -158 71614 -146 72390
rect -112 71614 -100 72390
rect -158 71602 -100 71614
rect 100 72390 158 72402
rect 100 71614 112 72390
rect 146 71614 158 72390
rect 100 71602 158 71614
rect -158 71354 -100 71366
rect -158 70578 -146 71354
rect -112 70578 -100 71354
rect -158 70566 -100 70578
rect 100 71354 158 71366
rect 100 70578 112 71354
rect 146 70578 158 71354
rect 100 70566 158 70578
rect -158 70318 -100 70330
rect -158 69542 -146 70318
rect -112 69542 -100 70318
rect -158 69530 -100 69542
rect 100 70318 158 70330
rect 100 69542 112 70318
rect 146 69542 158 70318
rect 100 69530 158 69542
rect -158 69282 -100 69294
rect -158 68506 -146 69282
rect -112 68506 -100 69282
rect -158 68494 -100 68506
rect 100 69282 158 69294
rect 100 68506 112 69282
rect 146 68506 158 69282
rect 100 68494 158 68506
rect -158 68246 -100 68258
rect -158 67470 -146 68246
rect -112 67470 -100 68246
rect -158 67458 -100 67470
rect 100 68246 158 68258
rect 100 67470 112 68246
rect 146 67470 158 68246
rect 100 67458 158 67470
rect -158 67210 -100 67222
rect -158 66434 -146 67210
rect -112 66434 -100 67210
rect -158 66422 -100 66434
rect 100 67210 158 67222
rect 100 66434 112 67210
rect 146 66434 158 67210
rect 100 66422 158 66434
rect -158 66174 -100 66186
rect -158 65398 -146 66174
rect -112 65398 -100 66174
rect -158 65386 -100 65398
rect 100 66174 158 66186
rect 100 65398 112 66174
rect 146 65398 158 66174
rect 100 65386 158 65398
rect -158 65138 -100 65150
rect -158 64362 -146 65138
rect -112 64362 -100 65138
rect -158 64350 -100 64362
rect 100 65138 158 65150
rect 100 64362 112 65138
rect 146 64362 158 65138
rect 100 64350 158 64362
rect -158 64102 -100 64114
rect -158 63326 -146 64102
rect -112 63326 -100 64102
rect -158 63314 -100 63326
rect 100 64102 158 64114
rect 100 63326 112 64102
rect 146 63326 158 64102
rect 100 63314 158 63326
rect -158 63066 -100 63078
rect -158 62290 -146 63066
rect -112 62290 -100 63066
rect -158 62278 -100 62290
rect 100 63066 158 63078
rect 100 62290 112 63066
rect 146 62290 158 63066
rect 100 62278 158 62290
rect -158 62030 -100 62042
rect -158 61254 -146 62030
rect -112 61254 -100 62030
rect -158 61242 -100 61254
rect 100 62030 158 62042
rect 100 61254 112 62030
rect 146 61254 158 62030
rect 100 61242 158 61254
rect -158 60994 -100 61006
rect -158 60218 -146 60994
rect -112 60218 -100 60994
rect -158 60206 -100 60218
rect 100 60994 158 61006
rect 100 60218 112 60994
rect 146 60218 158 60994
rect 100 60206 158 60218
rect -158 59958 -100 59970
rect -158 59182 -146 59958
rect -112 59182 -100 59958
rect -158 59170 -100 59182
rect 100 59958 158 59970
rect 100 59182 112 59958
rect 146 59182 158 59958
rect 100 59170 158 59182
rect -158 58922 -100 58934
rect -158 58146 -146 58922
rect -112 58146 -100 58922
rect -158 58134 -100 58146
rect 100 58922 158 58934
rect 100 58146 112 58922
rect 146 58146 158 58922
rect 100 58134 158 58146
rect -158 57886 -100 57898
rect -158 57110 -146 57886
rect -112 57110 -100 57886
rect -158 57098 -100 57110
rect 100 57886 158 57898
rect 100 57110 112 57886
rect 146 57110 158 57886
rect 100 57098 158 57110
rect -158 56850 -100 56862
rect -158 56074 -146 56850
rect -112 56074 -100 56850
rect -158 56062 -100 56074
rect 100 56850 158 56862
rect 100 56074 112 56850
rect 146 56074 158 56850
rect 100 56062 158 56074
rect -158 55814 -100 55826
rect -158 55038 -146 55814
rect -112 55038 -100 55814
rect -158 55026 -100 55038
rect 100 55814 158 55826
rect 100 55038 112 55814
rect 146 55038 158 55814
rect 100 55026 158 55038
rect -158 54778 -100 54790
rect -158 54002 -146 54778
rect -112 54002 -100 54778
rect -158 53990 -100 54002
rect 100 54778 158 54790
rect 100 54002 112 54778
rect 146 54002 158 54778
rect 100 53990 158 54002
rect -158 53742 -100 53754
rect -158 52966 -146 53742
rect -112 52966 -100 53742
rect -158 52954 -100 52966
rect 100 53742 158 53754
rect 100 52966 112 53742
rect 146 52966 158 53742
rect 100 52954 158 52966
rect -158 52706 -100 52718
rect -158 51930 -146 52706
rect -112 51930 -100 52706
rect -158 51918 -100 51930
rect 100 52706 158 52718
rect 100 51930 112 52706
rect 146 51930 158 52706
rect 100 51918 158 51930
rect -158 51670 -100 51682
rect -158 50894 -146 51670
rect -112 50894 -100 51670
rect -158 50882 -100 50894
rect 100 51670 158 51682
rect 100 50894 112 51670
rect 146 50894 158 51670
rect 100 50882 158 50894
rect -158 50634 -100 50646
rect -158 49858 -146 50634
rect -112 49858 -100 50634
rect -158 49846 -100 49858
rect 100 50634 158 50646
rect 100 49858 112 50634
rect 146 49858 158 50634
rect 100 49846 158 49858
rect -158 49598 -100 49610
rect -158 48822 -146 49598
rect -112 48822 -100 49598
rect -158 48810 -100 48822
rect 100 49598 158 49610
rect 100 48822 112 49598
rect 146 48822 158 49598
rect 100 48810 158 48822
rect -158 48562 -100 48574
rect -158 47786 -146 48562
rect -112 47786 -100 48562
rect -158 47774 -100 47786
rect 100 48562 158 48574
rect 100 47786 112 48562
rect 146 47786 158 48562
rect 100 47774 158 47786
rect -158 47526 -100 47538
rect -158 46750 -146 47526
rect -112 46750 -100 47526
rect -158 46738 -100 46750
rect 100 47526 158 47538
rect 100 46750 112 47526
rect 146 46750 158 47526
rect 100 46738 158 46750
rect -158 46490 -100 46502
rect -158 45714 -146 46490
rect -112 45714 -100 46490
rect -158 45702 -100 45714
rect 100 46490 158 46502
rect 100 45714 112 46490
rect 146 45714 158 46490
rect 100 45702 158 45714
rect -158 45454 -100 45466
rect -158 44678 -146 45454
rect -112 44678 -100 45454
rect -158 44666 -100 44678
rect 100 45454 158 45466
rect 100 44678 112 45454
rect 146 44678 158 45454
rect 100 44666 158 44678
rect -158 44418 -100 44430
rect -158 43642 -146 44418
rect -112 43642 -100 44418
rect -158 43630 -100 43642
rect 100 44418 158 44430
rect 100 43642 112 44418
rect 146 43642 158 44418
rect 100 43630 158 43642
rect -158 43382 -100 43394
rect -158 42606 -146 43382
rect -112 42606 -100 43382
rect -158 42594 -100 42606
rect 100 43382 158 43394
rect 100 42606 112 43382
rect 146 42606 158 43382
rect 100 42594 158 42606
rect -158 42346 -100 42358
rect -158 41570 -146 42346
rect -112 41570 -100 42346
rect -158 41558 -100 41570
rect 100 42346 158 42358
rect 100 41570 112 42346
rect 146 41570 158 42346
rect 100 41558 158 41570
rect -158 41310 -100 41322
rect -158 40534 -146 41310
rect -112 40534 -100 41310
rect -158 40522 -100 40534
rect 100 41310 158 41322
rect 100 40534 112 41310
rect 146 40534 158 41310
rect 100 40522 158 40534
rect -158 40274 -100 40286
rect -158 39498 -146 40274
rect -112 39498 -100 40274
rect -158 39486 -100 39498
rect 100 40274 158 40286
rect 100 39498 112 40274
rect 146 39498 158 40274
rect 100 39486 158 39498
rect -158 39238 -100 39250
rect -158 38462 -146 39238
rect -112 38462 -100 39238
rect -158 38450 -100 38462
rect 100 39238 158 39250
rect 100 38462 112 39238
rect 146 38462 158 39238
rect 100 38450 158 38462
rect -158 38202 -100 38214
rect -158 37426 -146 38202
rect -112 37426 -100 38202
rect -158 37414 -100 37426
rect 100 38202 158 38214
rect 100 37426 112 38202
rect 146 37426 158 38202
rect 100 37414 158 37426
rect -158 37166 -100 37178
rect -158 36390 -146 37166
rect -112 36390 -100 37166
rect -158 36378 -100 36390
rect 100 37166 158 37178
rect 100 36390 112 37166
rect 146 36390 158 37166
rect 100 36378 158 36390
rect -158 36130 -100 36142
rect -158 35354 -146 36130
rect -112 35354 -100 36130
rect -158 35342 -100 35354
rect 100 36130 158 36142
rect 100 35354 112 36130
rect 146 35354 158 36130
rect 100 35342 158 35354
rect -158 35094 -100 35106
rect -158 34318 -146 35094
rect -112 34318 -100 35094
rect -158 34306 -100 34318
rect 100 35094 158 35106
rect 100 34318 112 35094
rect 146 34318 158 35094
rect 100 34306 158 34318
rect -158 34058 -100 34070
rect -158 33282 -146 34058
rect -112 33282 -100 34058
rect -158 33270 -100 33282
rect 100 34058 158 34070
rect 100 33282 112 34058
rect 146 33282 158 34058
rect 100 33270 158 33282
rect -158 33022 -100 33034
rect -158 32246 -146 33022
rect -112 32246 -100 33022
rect -158 32234 -100 32246
rect 100 33022 158 33034
rect 100 32246 112 33022
rect 146 32246 158 33022
rect 100 32234 158 32246
rect -158 31986 -100 31998
rect -158 31210 -146 31986
rect -112 31210 -100 31986
rect -158 31198 -100 31210
rect 100 31986 158 31998
rect 100 31210 112 31986
rect 146 31210 158 31986
rect 100 31198 158 31210
rect -158 30950 -100 30962
rect -158 30174 -146 30950
rect -112 30174 -100 30950
rect -158 30162 -100 30174
rect 100 30950 158 30962
rect 100 30174 112 30950
rect 146 30174 158 30950
rect 100 30162 158 30174
rect -158 29914 -100 29926
rect -158 29138 -146 29914
rect -112 29138 -100 29914
rect -158 29126 -100 29138
rect 100 29914 158 29926
rect 100 29138 112 29914
rect 146 29138 158 29914
rect 100 29126 158 29138
rect -158 28878 -100 28890
rect -158 28102 -146 28878
rect -112 28102 -100 28878
rect -158 28090 -100 28102
rect 100 28878 158 28890
rect 100 28102 112 28878
rect 146 28102 158 28878
rect 100 28090 158 28102
rect -158 27842 -100 27854
rect -158 27066 -146 27842
rect -112 27066 -100 27842
rect -158 27054 -100 27066
rect 100 27842 158 27854
rect 100 27066 112 27842
rect 146 27066 158 27842
rect 100 27054 158 27066
rect -158 26806 -100 26818
rect -158 26030 -146 26806
rect -112 26030 -100 26806
rect -158 26018 -100 26030
rect 100 26806 158 26818
rect 100 26030 112 26806
rect 146 26030 158 26806
rect 100 26018 158 26030
rect -158 25770 -100 25782
rect -158 24994 -146 25770
rect -112 24994 -100 25770
rect -158 24982 -100 24994
rect 100 25770 158 25782
rect 100 24994 112 25770
rect 146 24994 158 25770
rect 100 24982 158 24994
rect -158 24734 -100 24746
rect -158 23958 -146 24734
rect -112 23958 -100 24734
rect -158 23946 -100 23958
rect 100 24734 158 24746
rect 100 23958 112 24734
rect 146 23958 158 24734
rect 100 23946 158 23958
rect -158 23698 -100 23710
rect -158 22922 -146 23698
rect -112 22922 -100 23698
rect -158 22910 -100 22922
rect 100 23698 158 23710
rect 100 22922 112 23698
rect 146 22922 158 23698
rect 100 22910 158 22922
rect -158 22662 -100 22674
rect -158 21886 -146 22662
rect -112 21886 -100 22662
rect -158 21874 -100 21886
rect 100 22662 158 22674
rect 100 21886 112 22662
rect 146 21886 158 22662
rect 100 21874 158 21886
rect -158 21626 -100 21638
rect -158 20850 -146 21626
rect -112 20850 -100 21626
rect -158 20838 -100 20850
rect 100 21626 158 21638
rect 100 20850 112 21626
rect 146 20850 158 21626
rect 100 20838 158 20850
rect -158 20590 -100 20602
rect -158 19814 -146 20590
rect -112 19814 -100 20590
rect -158 19802 -100 19814
rect 100 20590 158 20602
rect 100 19814 112 20590
rect 146 19814 158 20590
rect 100 19802 158 19814
rect -158 19554 -100 19566
rect -158 18778 -146 19554
rect -112 18778 -100 19554
rect -158 18766 -100 18778
rect 100 19554 158 19566
rect 100 18778 112 19554
rect 146 18778 158 19554
rect 100 18766 158 18778
rect -158 18518 -100 18530
rect -158 17742 -146 18518
rect -112 17742 -100 18518
rect -158 17730 -100 17742
rect 100 18518 158 18530
rect 100 17742 112 18518
rect 146 17742 158 18518
rect 100 17730 158 17742
rect -158 17482 -100 17494
rect -158 16706 -146 17482
rect -112 16706 -100 17482
rect -158 16694 -100 16706
rect 100 17482 158 17494
rect 100 16706 112 17482
rect 146 16706 158 17482
rect 100 16694 158 16706
rect -158 16446 -100 16458
rect -158 15670 -146 16446
rect -112 15670 -100 16446
rect -158 15658 -100 15670
rect 100 16446 158 16458
rect 100 15670 112 16446
rect 146 15670 158 16446
rect 100 15658 158 15670
rect -158 15410 -100 15422
rect -158 14634 -146 15410
rect -112 14634 -100 15410
rect -158 14622 -100 14634
rect 100 15410 158 15422
rect 100 14634 112 15410
rect 146 14634 158 15410
rect 100 14622 158 14634
rect -158 14374 -100 14386
rect -158 13598 -146 14374
rect -112 13598 -100 14374
rect -158 13586 -100 13598
rect 100 14374 158 14386
rect 100 13598 112 14374
rect 146 13598 158 14374
rect 100 13586 158 13598
rect -158 13338 -100 13350
rect -158 12562 -146 13338
rect -112 12562 -100 13338
rect -158 12550 -100 12562
rect 100 13338 158 13350
rect 100 12562 112 13338
rect 146 12562 158 13338
rect 100 12550 158 12562
rect -158 12302 -100 12314
rect -158 11526 -146 12302
rect -112 11526 -100 12302
rect -158 11514 -100 11526
rect 100 12302 158 12314
rect 100 11526 112 12302
rect 146 11526 158 12302
rect 100 11514 158 11526
rect -158 11266 -100 11278
rect -158 10490 -146 11266
rect -112 10490 -100 11266
rect -158 10478 -100 10490
rect 100 11266 158 11278
rect 100 10490 112 11266
rect 146 10490 158 11266
rect 100 10478 158 10490
rect -158 10230 -100 10242
rect -158 9454 -146 10230
rect -112 9454 -100 10230
rect -158 9442 -100 9454
rect 100 10230 158 10242
rect 100 9454 112 10230
rect 146 9454 158 10230
rect 100 9442 158 9454
rect -158 9194 -100 9206
rect -158 8418 -146 9194
rect -112 8418 -100 9194
rect -158 8406 -100 8418
rect 100 9194 158 9206
rect 100 8418 112 9194
rect 146 8418 158 9194
rect 100 8406 158 8418
rect -158 8158 -100 8170
rect -158 7382 -146 8158
rect -112 7382 -100 8158
rect -158 7370 -100 7382
rect 100 8158 158 8170
rect 100 7382 112 8158
rect 146 7382 158 8158
rect 100 7370 158 7382
rect -158 7122 -100 7134
rect -158 6346 -146 7122
rect -112 6346 -100 7122
rect -158 6334 -100 6346
rect 100 7122 158 7134
rect 100 6346 112 7122
rect 146 6346 158 7122
rect 100 6334 158 6346
rect -158 6086 -100 6098
rect -158 5310 -146 6086
rect -112 5310 -100 6086
rect -158 5298 -100 5310
rect 100 6086 158 6098
rect 100 5310 112 6086
rect 146 5310 158 6086
rect 100 5298 158 5310
rect -158 5050 -100 5062
rect -158 4274 -146 5050
rect -112 4274 -100 5050
rect -158 4262 -100 4274
rect 100 5050 158 5062
rect 100 4274 112 5050
rect 146 4274 158 5050
rect 100 4262 158 4274
rect -158 4014 -100 4026
rect -158 3238 -146 4014
rect -112 3238 -100 4014
rect -158 3226 -100 3238
rect 100 4014 158 4026
rect 100 3238 112 4014
rect 146 3238 158 4014
rect 100 3226 158 3238
rect -158 2978 -100 2990
rect -158 2202 -146 2978
rect -112 2202 -100 2978
rect -158 2190 -100 2202
rect 100 2978 158 2990
rect 100 2202 112 2978
rect 146 2202 158 2978
rect 100 2190 158 2202
rect -158 1942 -100 1954
rect -158 1166 -146 1942
rect -112 1166 -100 1942
rect -158 1154 -100 1166
rect 100 1942 158 1954
rect 100 1166 112 1942
rect 146 1166 158 1942
rect 100 1154 158 1166
rect -158 906 -100 918
rect -158 130 -146 906
rect -112 130 -100 906
rect -158 118 -100 130
rect 100 906 158 918
rect 100 130 112 906
rect 146 130 158 906
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -906 -146 -130
rect -112 -906 -100 -130
rect -158 -918 -100 -906
rect 100 -130 158 -118
rect 100 -906 112 -130
rect 146 -906 158 -130
rect 100 -918 158 -906
rect -158 -1166 -100 -1154
rect -158 -1942 -146 -1166
rect -112 -1942 -100 -1166
rect -158 -1954 -100 -1942
rect 100 -1166 158 -1154
rect 100 -1942 112 -1166
rect 146 -1942 158 -1166
rect 100 -1954 158 -1942
rect -158 -2202 -100 -2190
rect -158 -2978 -146 -2202
rect -112 -2978 -100 -2202
rect -158 -2990 -100 -2978
rect 100 -2202 158 -2190
rect 100 -2978 112 -2202
rect 146 -2978 158 -2202
rect 100 -2990 158 -2978
rect -158 -3238 -100 -3226
rect -158 -4014 -146 -3238
rect -112 -4014 -100 -3238
rect -158 -4026 -100 -4014
rect 100 -3238 158 -3226
rect 100 -4014 112 -3238
rect 146 -4014 158 -3238
rect 100 -4026 158 -4014
rect -158 -4274 -100 -4262
rect -158 -5050 -146 -4274
rect -112 -5050 -100 -4274
rect -158 -5062 -100 -5050
rect 100 -4274 158 -4262
rect 100 -5050 112 -4274
rect 146 -5050 158 -4274
rect 100 -5062 158 -5050
rect -158 -5310 -100 -5298
rect -158 -6086 -146 -5310
rect -112 -6086 -100 -5310
rect -158 -6098 -100 -6086
rect 100 -5310 158 -5298
rect 100 -6086 112 -5310
rect 146 -6086 158 -5310
rect 100 -6098 158 -6086
rect -158 -6346 -100 -6334
rect -158 -7122 -146 -6346
rect -112 -7122 -100 -6346
rect -158 -7134 -100 -7122
rect 100 -6346 158 -6334
rect 100 -7122 112 -6346
rect 146 -7122 158 -6346
rect 100 -7134 158 -7122
rect -158 -7382 -100 -7370
rect -158 -8158 -146 -7382
rect -112 -8158 -100 -7382
rect -158 -8170 -100 -8158
rect 100 -7382 158 -7370
rect 100 -8158 112 -7382
rect 146 -8158 158 -7382
rect 100 -8170 158 -8158
rect -158 -8418 -100 -8406
rect -158 -9194 -146 -8418
rect -112 -9194 -100 -8418
rect -158 -9206 -100 -9194
rect 100 -8418 158 -8406
rect 100 -9194 112 -8418
rect 146 -9194 158 -8418
rect 100 -9206 158 -9194
rect -158 -9454 -100 -9442
rect -158 -10230 -146 -9454
rect -112 -10230 -100 -9454
rect -158 -10242 -100 -10230
rect 100 -9454 158 -9442
rect 100 -10230 112 -9454
rect 146 -10230 158 -9454
rect 100 -10242 158 -10230
rect -158 -10490 -100 -10478
rect -158 -11266 -146 -10490
rect -112 -11266 -100 -10490
rect -158 -11278 -100 -11266
rect 100 -10490 158 -10478
rect 100 -11266 112 -10490
rect 146 -11266 158 -10490
rect 100 -11278 158 -11266
rect -158 -11526 -100 -11514
rect -158 -12302 -146 -11526
rect -112 -12302 -100 -11526
rect -158 -12314 -100 -12302
rect 100 -11526 158 -11514
rect 100 -12302 112 -11526
rect 146 -12302 158 -11526
rect 100 -12314 158 -12302
rect -158 -12562 -100 -12550
rect -158 -13338 -146 -12562
rect -112 -13338 -100 -12562
rect -158 -13350 -100 -13338
rect 100 -12562 158 -12550
rect 100 -13338 112 -12562
rect 146 -13338 158 -12562
rect 100 -13350 158 -13338
rect -158 -13598 -100 -13586
rect -158 -14374 -146 -13598
rect -112 -14374 -100 -13598
rect -158 -14386 -100 -14374
rect 100 -13598 158 -13586
rect 100 -14374 112 -13598
rect 146 -14374 158 -13598
rect 100 -14386 158 -14374
rect -158 -14634 -100 -14622
rect -158 -15410 -146 -14634
rect -112 -15410 -100 -14634
rect -158 -15422 -100 -15410
rect 100 -14634 158 -14622
rect 100 -15410 112 -14634
rect 146 -15410 158 -14634
rect 100 -15422 158 -15410
rect -158 -15670 -100 -15658
rect -158 -16446 -146 -15670
rect -112 -16446 -100 -15670
rect -158 -16458 -100 -16446
rect 100 -15670 158 -15658
rect 100 -16446 112 -15670
rect 146 -16446 158 -15670
rect 100 -16458 158 -16446
rect -158 -16706 -100 -16694
rect -158 -17482 -146 -16706
rect -112 -17482 -100 -16706
rect -158 -17494 -100 -17482
rect 100 -16706 158 -16694
rect 100 -17482 112 -16706
rect 146 -17482 158 -16706
rect 100 -17494 158 -17482
rect -158 -17742 -100 -17730
rect -158 -18518 -146 -17742
rect -112 -18518 -100 -17742
rect -158 -18530 -100 -18518
rect 100 -17742 158 -17730
rect 100 -18518 112 -17742
rect 146 -18518 158 -17742
rect 100 -18530 158 -18518
rect -158 -18778 -100 -18766
rect -158 -19554 -146 -18778
rect -112 -19554 -100 -18778
rect -158 -19566 -100 -19554
rect 100 -18778 158 -18766
rect 100 -19554 112 -18778
rect 146 -19554 158 -18778
rect 100 -19566 158 -19554
rect -158 -19814 -100 -19802
rect -158 -20590 -146 -19814
rect -112 -20590 -100 -19814
rect -158 -20602 -100 -20590
rect 100 -19814 158 -19802
rect 100 -20590 112 -19814
rect 146 -20590 158 -19814
rect 100 -20602 158 -20590
rect -158 -20850 -100 -20838
rect -158 -21626 -146 -20850
rect -112 -21626 -100 -20850
rect -158 -21638 -100 -21626
rect 100 -20850 158 -20838
rect 100 -21626 112 -20850
rect 146 -21626 158 -20850
rect 100 -21638 158 -21626
rect -158 -21886 -100 -21874
rect -158 -22662 -146 -21886
rect -112 -22662 -100 -21886
rect -158 -22674 -100 -22662
rect 100 -21886 158 -21874
rect 100 -22662 112 -21886
rect 146 -22662 158 -21886
rect 100 -22674 158 -22662
rect -158 -22922 -100 -22910
rect -158 -23698 -146 -22922
rect -112 -23698 -100 -22922
rect -158 -23710 -100 -23698
rect 100 -22922 158 -22910
rect 100 -23698 112 -22922
rect 146 -23698 158 -22922
rect 100 -23710 158 -23698
rect -158 -23958 -100 -23946
rect -158 -24734 -146 -23958
rect -112 -24734 -100 -23958
rect -158 -24746 -100 -24734
rect 100 -23958 158 -23946
rect 100 -24734 112 -23958
rect 146 -24734 158 -23958
rect 100 -24746 158 -24734
rect -158 -24994 -100 -24982
rect -158 -25770 -146 -24994
rect -112 -25770 -100 -24994
rect -158 -25782 -100 -25770
rect 100 -24994 158 -24982
rect 100 -25770 112 -24994
rect 146 -25770 158 -24994
rect 100 -25782 158 -25770
rect -158 -26030 -100 -26018
rect -158 -26806 -146 -26030
rect -112 -26806 -100 -26030
rect -158 -26818 -100 -26806
rect 100 -26030 158 -26018
rect 100 -26806 112 -26030
rect 146 -26806 158 -26030
rect 100 -26818 158 -26806
rect -158 -27066 -100 -27054
rect -158 -27842 -146 -27066
rect -112 -27842 -100 -27066
rect -158 -27854 -100 -27842
rect 100 -27066 158 -27054
rect 100 -27842 112 -27066
rect 146 -27842 158 -27066
rect 100 -27854 158 -27842
rect -158 -28102 -100 -28090
rect -158 -28878 -146 -28102
rect -112 -28878 -100 -28102
rect -158 -28890 -100 -28878
rect 100 -28102 158 -28090
rect 100 -28878 112 -28102
rect 146 -28878 158 -28102
rect 100 -28890 158 -28878
rect -158 -29138 -100 -29126
rect -158 -29914 -146 -29138
rect -112 -29914 -100 -29138
rect -158 -29926 -100 -29914
rect 100 -29138 158 -29126
rect 100 -29914 112 -29138
rect 146 -29914 158 -29138
rect 100 -29926 158 -29914
rect -158 -30174 -100 -30162
rect -158 -30950 -146 -30174
rect -112 -30950 -100 -30174
rect -158 -30962 -100 -30950
rect 100 -30174 158 -30162
rect 100 -30950 112 -30174
rect 146 -30950 158 -30174
rect 100 -30962 158 -30950
rect -158 -31210 -100 -31198
rect -158 -31986 -146 -31210
rect -112 -31986 -100 -31210
rect -158 -31998 -100 -31986
rect 100 -31210 158 -31198
rect 100 -31986 112 -31210
rect 146 -31986 158 -31210
rect 100 -31998 158 -31986
rect -158 -32246 -100 -32234
rect -158 -33022 -146 -32246
rect -112 -33022 -100 -32246
rect -158 -33034 -100 -33022
rect 100 -32246 158 -32234
rect 100 -33022 112 -32246
rect 146 -33022 158 -32246
rect 100 -33034 158 -33022
rect -158 -33282 -100 -33270
rect -158 -34058 -146 -33282
rect -112 -34058 -100 -33282
rect -158 -34070 -100 -34058
rect 100 -33282 158 -33270
rect 100 -34058 112 -33282
rect 146 -34058 158 -33282
rect 100 -34070 158 -34058
rect -158 -34318 -100 -34306
rect -158 -35094 -146 -34318
rect -112 -35094 -100 -34318
rect -158 -35106 -100 -35094
rect 100 -34318 158 -34306
rect 100 -35094 112 -34318
rect 146 -35094 158 -34318
rect 100 -35106 158 -35094
rect -158 -35354 -100 -35342
rect -158 -36130 -146 -35354
rect -112 -36130 -100 -35354
rect -158 -36142 -100 -36130
rect 100 -35354 158 -35342
rect 100 -36130 112 -35354
rect 146 -36130 158 -35354
rect 100 -36142 158 -36130
rect -158 -36390 -100 -36378
rect -158 -37166 -146 -36390
rect -112 -37166 -100 -36390
rect -158 -37178 -100 -37166
rect 100 -36390 158 -36378
rect 100 -37166 112 -36390
rect 146 -37166 158 -36390
rect 100 -37178 158 -37166
rect -158 -37426 -100 -37414
rect -158 -38202 -146 -37426
rect -112 -38202 -100 -37426
rect -158 -38214 -100 -38202
rect 100 -37426 158 -37414
rect 100 -38202 112 -37426
rect 146 -38202 158 -37426
rect 100 -38214 158 -38202
rect -158 -38462 -100 -38450
rect -158 -39238 -146 -38462
rect -112 -39238 -100 -38462
rect -158 -39250 -100 -39238
rect 100 -38462 158 -38450
rect 100 -39238 112 -38462
rect 146 -39238 158 -38462
rect 100 -39250 158 -39238
rect -158 -39498 -100 -39486
rect -158 -40274 -146 -39498
rect -112 -40274 -100 -39498
rect -158 -40286 -100 -40274
rect 100 -39498 158 -39486
rect 100 -40274 112 -39498
rect 146 -40274 158 -39498
rect 100 -40286 158 -40274
rect -158 -40534 -100 -40522
rect -158 -41310 -146 -40534
rect -112 -41310 -100 -40534
rect -158 -41322 -100 -41310
rect 100 -40534 158 -40522
rect 100 -41310 112 -40534
rect 146 -41310 158 -40534
rect 100 -41322 158 -41310
rect -158 -41570 -100 -41558
rect -158 -42346 -146 -41570
rect -112 -42346 -100 -41570
rect -158 -42358 -100 -42346
rect 100 -41570 158 -41558
rect 100 -42346 112 -41570
rect 146 -42346 158 -41570
rect 100 -42358 158 -42346
rect -158 -42606 -100 -42594
rect -158 -43382 -146 -42606
rect -112 -43382 -100 -42606
rect -158 -43394 -100 -43382
rect 100 -42606 158 -42594
rect 100 -43382 112 -42606
rect 146 -43382 158 -42606
rect 100 -43394 158 -43382
rect -158 -43642 -100 -43630
rect -158 -44418 -146 -43642
rect -112 -44418 -100 -43642
rect -158 -44430 -100 -44418
rect 100 -43642 158 -43630
rect 100 -44418 112 -43642
rect 146 -44418 158 -43642
rect 100 -44430 158 -44418
rect -158 -44678 -100 -44666
rect -158 -45454 -146 -44678
rect -112 -45454 -100 -44678
rect -158 -45466 -100 -45454
rect 100 -44678 158 -44666
rect 100 -45454 112 -44678
rect 146 -45454 158 -44678
rect 100 -45466 158 -45454
rect -158 -45714 -100 -45702
rect -158 -46490 -146 -45714
rect -112 -46490 -100 -45714
rect -158 -46502 -100 -46490
rect 100 -45714 158 -45702
rect 100 -46490 112 -45714
rect 146 -46490 158 -45714
rect 100 -46502 158 -46490
rect -158 -46750 -100 -46738
rect -158 -47526 -146 -46750
rect -112 -47526 -100 -46750
rect -158 -47538 -100 -47526
rect 100 -46750 158 -46738
rect 100 -47526 112 -46750
rect 146 -47526 158 -46750
rect 100 -47538 158 -47526
rect -158 -47786 -100 -47774
rect -158 -48562 -146 -47786
rect -112 -48562 -100 -47786
rect -158 -48574 -100 -48562
rect 100 -47786 158 -47774
rect 100 -48562 112 -47786
rect 146 -48562 158 -47786
rect 100 -48574 158 -48562
rect -158 -48822 -100 -48810
rect -158 -49598 -146 -48822
rect -112 -49598 -100 -48822
rect -158 -49610 -100 -49598
rect 100 -48822 158 -48810
rect 100 -49598 112 -48822
rect 146 -49598 158 -48822
rect 100 -49610 158 -49598
rect -158 -49858 -100 -49846
rect -158 -50634 -146 -49858
rect -112 -50634 -100 -49858
rect -158 -50646 -100 -50634
rect 100 -49858 158 -49846
rect 100 -50634 112 -49858
rect 146 -50634 158 -49858
rect 100 -50646 158 -50634
rect -158 -50894 -100 -50882
rect -158 -51670 -146 -50894
rect -112 -51670 -100 -50894
rect -158 -51682 -100 -51670
rect 100 -50894 158 -50882
rect 100 -51670 112 -50894
rect 146 -51670 158 -50894
rect 100 -51682 158 -51670
rect -158 -51930 -100 -51918
rect -158 -52706 -146 -51930
rect -112 -52706 -100 -51930
rect -158 -52718 -100 -52706
rect 100 -51930 158 -51918
rect 100 -52706 112 -51930
rect 146 -52706 158 -51930
rect 100 -52718 158 -52706
rect -158 -52966 -100 -52954
rect -158 -53742 -146 -52966
rect -112 -53742 -100 -52966
rect -158 -53754 -100 -53742
rect 100 -52966 158 -52954
rect 100 -53742 112 -52966
rect 146 -53742 158 -52966
rect 100 -53754 158 -53742
rect -158 -54002 -100 -53990
rect -158 -54778 -146 -54002
rect -112 -54778 -100 -54002
rect -158 -54790 -100 -54778
rect 100 -54002 158 -53990
rect 100 -54778 112 -54002
rect 146 -54778 158 -54002
rect 100 -54790 158 -54778
rect -158 -55038 -100 -55026
rect -158 -55814 -146 -55038
rect -112 -55814 -100 -55038
rect -158 -55826 -100 -55814
rect 100 -55038 158 -55026
rect 100 -55814 112 -55038
rect 146 -55814 158 -55038
rect 100 -55826 158 -55814
rect -158 -56074 -100 -56062
rect -158 -56850 -146 -56074
rect -112 -56850 -100 -56074
rect -158 -56862 -100 -56850
rect 100 -56074 158 -56062
rect 100 -56850 112 -56074
rect 146 -56850 158 -56074
rect 100 -56862 158 -56850
rect -158 -57110 -100 -57098
rect -158 -57886 -146 -57110
rect -112 -57886 -100 -57110
rect -158 -57898 -100 -57886
rect 100 -57110 158 -57098
rect 100 -57886 112 -57110
rect 146 -57886 158 -57110
rect 100 -57898 158 -57886
rect -158 -58146 -100 -58134
rect -158 -58922 -146 -58146
rect -112 -58922 -100 -58146
rect -158 -58934 -100 -58922
rect 100 -58146 158 -58134
rect 100 -58922 112 -58146
rect 146 -58922 158 -58146
rect 100 -58934 158 -58922
rect -158 -59182 -100 -59170
rect -158 -59958 -146 -59182
rect -112 -59958 -100 -59182
rect -158 -59970 -100 -59958
rect 100 -59182 158 -59170
rect 100 -59958 112 -59182
rect 146 -59958 158 -59182
rect 100 -59970 158 -59958
rect -158 -60218 -100 -60206
rect -158 -60994 -146 -60218
rect -112 -60994 -100 -60218
rect -158 -61006 -100 -60994
rect 100 -60218 158 -60206
rect 100 -60994 112 -60218
rect 146 -60994 158 -60218
rect 100 -61006 158 -60994
rect -158 -61254 -100 -61242
rect -158 -62030 -146 -61254
rect -112 -62030 -100 -61254
rect -158 -62042 -100 -62030
rect 100 -61254 158 -61242
rect 100 -62030 112 -61254
rect 146 -62030 158 -61254
rect 100 -62042 158 -62030
rect -158 -62290 -100 -62278
rect -158 -63066 -146 -62290
rect -112 -63066 -100 -62290
rect -158 -63078 -100 -63066
rect 100 -62290 158 -62278
rect 100 -63066 112 -62290
rect 146 -63066 158 -62290
rect 100 -63078 158 -63066
rect -158 -63326 -100 -63314
rect -158 -64102 -146 -63326
rect -112 -64102 -100 -63326
rect -158 -64114 -100 -64102
rect 100 -63326 158 -63314
rect 100 -64102 112 -63326
rect 146 -64102 158 -63326
rect 100 -64114 158 -64102
rect -158 -64362 -100 -64350
rect -158 -65138 -146 -64362
rect -112 -65138 -100 -64362
rect -158 -65150 -100 -65138
rect 100 -64362 158 -64350
rect 100 -65138 112 -64362
rect 146 -65138 158 -64362
rect 100 -65150 158 -65138
rect -158 -65398 -100 -65386
rect -158 -66174 -146 -65398
rect -112 -66174 -100 -65398
rect -158 -66186 -100 -66174
rect 100 -65398 158 -65386
rect 100 -66174 112 -65398
rect 146 -66174 158 -65398
rect 100 -66186 158 -66174
rect -158 -66434 -100 -66422
rect -158 -67210 -146 -66434
rect -112 -67210 -100 -66434
rect -158 -67222 -100 -67210
rect 100 -66434 158 -66422
rect 100 -67210 112 -66434
rect 146 -67210 158 -66434
rect 100 -67222 158 -67210
rect -158 -67470 -100 -67458
rect -158 -68246 -146 -67470
rect -112 -68246 -100 -67470
rect -158 -68258 -100 -68246
rect 100 -67470 158 -67458
rect 100 -68246 112 -67470
rect 146 -68246 158 -67470
rect 100 -68258 158 -68246
rect -158 -68506 -100 -68494
rect -158 -69282 -146 -68506
rect -112 -69282 -100 -68506
rect -158 -69294 -100 -69282
rect 100 -68506 158 -68494
rect 100 -69282 112 -68506
rect 146 -69282 158 -68506
rect 100 -69294 158 -69282
rect -158 -69542 -100 -69530
rect -158 -70318 -146 -69542
rect -112 -70318 -100 -69542
rect -158 -70330 -100 -70318
rect 100 -69542 158 -69530
rect 100 -70318 112 -69542
rect 146 -70318 158 -69542
rect 100 -70330 158 -70318
rect -158 -70578 -100 -70566
rect -158 -71354 -146 -70578
rect -112 -71354 -100 -70578
rect -158 -71366 -100 -71354
rect 100 -70578 158 -70566
rect 100 -71354 112 -70578
rect 146 -71354 158 -70578
rect 100 -71366 158 -71354
rect -158 -71614 -100 -71602
rect -158 -72390 -146 -71614
rect -112 -72390 -100 -71614
rect -158 -72402 -100 -72390
rect 100 -71614 158 -71602
rect 100 -72390 112 -71614
rect 146 -72390 158 -71614
rect 100 -72402 158 -72390
rect -158 -72650 -100 -72638
rect -158 -73426 -146 -72650
rect -112 -73426 -100 -72650
rect -158 -73438 -100 -73426
rect 100 -72650 158 -72638
rect 100 -73426 112 -72650
rect 146 -73426 158 -72650
rect 100 -73438 158 -73426
rect -158 -73686 -100 -73674
rect -158 -74462 -146 -73686
rect -112 -74462 -100 -73686
rect -158 -74474 -100 -74462
rect 100 -73686 158 -73674
rect 100 -74462 112 -73686
rect 146 -74462 158 -73686
rect 100 -74474 158 -74462
rect -158 -74722 -100 -74710
rect -158 -75498 -146 -74722
rect -112 -75498 -100 -74722
rect -158 -75510 -100 -75498
rect 100 -74722 158 -74710
rect 100 -75498 112 -74722
rect 146 -75498 158 -74722
rect 100 -75510 158 -75498
rect -158 -75758 -100 -75746
rect -158 -76534 -146 -75758
rect -112 -76534 -100 -75758
rect -158 -76546 -100 -76534
rect 100 -75758 158 -75746
rect 100 -76534 112 -75758
rect 146 -76534 158 -75758
rect 100 -76546 158 -76534
rect -158 -76794 -100 -76782
rect -158 -77570 -146 -76794
rect -112 -77570 -100 -76794
rect -158 -77582 -100 -77570
rect 100 -76794 158 -76782
rect 100 -77570 112 -76794
rect 146 -77570 158 -76794
rect 100 -77582 158 -77570
rect -158 -77830 -100 -77818
rect -158 -78606 -146 -77830
rect -112 -78606 -100 -77830
rect -158 -78618 -100 -78606
rect 100 -77830 158 -77818
rect 100 -78606 112 -77830
rect 146 -78606 158 -77830
rect 100 -78618 158 -78606
rect -158 -78866 -100 -78854
rect -158 -79642 -146 -78866
rect -112 -79642 -100 -78866
rect -158 -79654 -100 -79642
rect 100 -78866 158 -78854
rect 100 -79642 112 -78866
rect 146 -79642 158 -78866
rect 100 -79654 158 -79642
rect -158 -79902 -100 -79890
rect -158 -80678 -146 -79902
rect -112 -80678 -100 -79902
rect -158 -80690 -100 -80678
rect 100 -79902 158 -79890
rect 100 -80678 112 -79902
rect 146 -80678 158 -79902
rect 100 -80690 158 -80678
rect -158 -80938 -100 -80926
rect -158 -81714 -146 -80938
rect -112 -81714 -100 -80938
rect -158 -81726 -100 -81714
rect 100 -80938 158 -80926
rect 100 -81714 112 -80938
rect 146 -81714 158 -80938
rect 100 -81726 158 -81714
rect -158 -81974 -100 -81962
rect -158 -82750 -146 -81974
rect -112 -82750 -100 -81974
rect -158 -82762 -100 -82750
rect 100 -81974 158 -81962
rect 100 -82750 112 -81974
rect 146 -82750 158 -81974
rect 100 -82762 158 -82750
rect -158 -83010 -100 -82998
rect -158 -83786 -146 -83010
rect -112 -83786 -100 -83010
rect -158 -83798 -100 -83786
rect 100 -83010 158 -82998
rect 100 -83786 112 -83010
rect 146 -83786 158 -83010
rect 100 -83798 158 -83786
rect -158 -84046 -100 -84034
rect -158 -84822 -146 -84046
rect -112 -84822 -100 -84046
rect -158 -84834 -100 -84822
rect 100 -84046 158 -84034
rect 100 -84822 112 -84046
rect 146 -84822 158 -84046
rect 100 -84834 158 -84822
rect -158 -85082 -100 -85070
rect -158 -85858 -146 -85082
rect -112 -85858 -100 -85082
rect -158 -85870 -100 -85858
rect 100 -85082 158 -85070
rect 100 -85858 112 -85082
rect 146 -85858 158 -85082
rect 100 -85870 158 -85858
rect -158 -86118 -100 -86106
rect -158 -86894 -146 -86118
rect -112 -86894 -100 -86118
rect -158 -86906 -100 -86894
rect 100 -86118 158 -86106
rect 100 -86894 112 -86118
rect 146 -86894 158 -86118
rect 100 -86906 158 -86894
rect -158 -87154 -100 -87142
rect -158 -87930 -146 -87154
rect -112 -87930 -100 -87154
rect -158 -87942 -100 -87930
rect 100 -87154 158 -87142
rect 100 -87930 112 -87154
rect 146 -87930 158 -87154
rect 100 -87942 158 -87930
rect -158 -88190 -100 -88178
rect -158 -88966 -146 -88190
rect -112 -88966 -100 -88190
rect -158 -88978 -100 -88966
rect 100 -88190 158 -88178
rect 100 -88966 112 -88190
rect 146 -88966 158 -88190
rect 100 -88978 158 -88966
rect -158 -89226 -100 -89214
rect -158 -90002 -146 -89226
rect -112 -90002 -100 -89226
rect -158 -90014 -100 -90002
rect 100 -89226 158 -89214
rect 100 -90002 112 -89226
rect 146 -90002 158 -89226
rect 100 -90014 158 -90002
rect -158 -90262 -100 -90250
rect -158 -91038 -146 -90262
rect -112 -91038 -100 -90262
rect -158 -91050 -100 -91038
rect 100 -90262 158 -90250
rect 100 -91038 112 -90262
rect 146 -91038 158 -90262
rect 100 -91050 158 -91038
rect -158 -91298 -100 -91286
rect -158 -92074 -146 -91298
rect -112 -92074 -100 -91298
rect -158 -92086 -100 -92074
rect 100 -91298 158 -91286
rect 100 -92074 112 -91298
rect 146 -92074 158 -91298
rect 100 -92086 158 -92074
rect -158 -92334 -100 -92322
rect -158 -93110 -146 -92334
rect -112 -93110 -100 -92334
rect -158 -93122 -100 -93110
rect 100 -92334 158 -92322
rect 100 -93110 112 -92334
rect 146 -93110 158 -92334
rect 100 -93122 158 -93110
rect -158 -93370 -100 -93358
rect -158 -94146 -146 -93370
rect -112 -94146 -100 -93370
rect -158 -94158 -100 -94146
rect 100 -93370 158 -93358
rect 100 -94146 112 -93370
rect 146 -94146 158 -93370
rect 100 -94158 158 -94146
rect -158 -94406 -100 -94394
rect -158 -95182 -146 -94406
rect -112 -95182 -100 -94406
rect -158 -95194 -100 -95182
rect 100 -94406 158 -94394
rect 100 -95182 112 -94406
rect 146 -95182 158 -94406
rect 100 -95194 158 -95182
rect -158 -95442 -100 -95430
rect -158 -96218 -146 -95442
rect -112 -96218 -100 -95442
rect -158 -96230 -100 -96218
rect 100 -95442 158 -95430
rect 100 -96218 112 -95442
rect 146 -96218 158 -95442
rect 100 -96230 158 -96218
rect -158 -96478 -100 -96466
rect -158 -97254 -146 -96478
rect -112 -97254 -100 -96478
rect -158 -97266 -100 -97254
rect 100 -96478 158 -96466
rect 100 -97254 112 -96478
rect 146 -97254 158 -96478
rect 100 -97266 158 -97254
rect -158 -97514 -100 -97502
rect -158 -98290 -146 -97514
rect -112 -98290 -100 -97514
rect -158 -98302 -100 -98290
rect 100 -97514 158 -97502
rect 100 -98290 112 -97514
rect 146 -98290 158 -97514
rect 100 -98302 158 -98290
rect -158 -98550 -100 -98538
rect -158 -99326 -146 -98550
rect -112 -99326 -100 -98550
rect -158 -99338 -100 -99326
rect 100 -98550 158 -98538
rect 100 -99326 112 -98550
rect 146 -99326 158 -98550
rect 100 -99338 158 -99326
rect -158 -99586 -100 -99574
rect -158 -100362 -146 -99586
rect -112 -100362 -100 -99586
rect -158 -100374 -100 -100362
rect 100 -99586 158 -99574
rect 100 -100362 112 -99586
rect 146 -100362 158 -99586
rect 100 -100374 158 -100362
rect -158 -100622 -100 -100610
rect -158 -101398 -146 -100622
rect -112 -101398 -100 -100622
rect -158 -101410 -100 -101398
rect 100 -100622 158 -100610
rect 100 -101398 112 -100622
rect 146 -101398 158 -100622
rect 100 -101410 158 -101398
rect -158 -101658 -100 -101646
rect -158 -102434 -146 -101658
rect -112 -102434 -100 -101658
rect -158 -102446 -100 -102434
rect 100 -101658 158 -101646
rect 100 -102434 112 -101658
rect 146 -102434 158 -101658
rect 100 -102446 158 -102434
rect -158 -102694 -100 -102682
rect -158 -103470 -146 -102694
rect -112 -103470 -100 -102694
rect -158 -103482 -100 -103470
rect 100 -102694 158 -102682
rect 100 -103470 112 -102694
rect 146 -103470 158 -102694
rect 100 -103482 158 -103470
rect -158 -103730 -100 -103718
rect -158 -104506 -146 -103730
rect -112 -104506 -100 -103730
rect -158 -104518 -100 -104506
rect 100 -103730 158 -103718
rect 100 -104506 112 -103730
rect 146 -104506 158 -103730
rect 100 -104518 158 -104506
rect -158 -104766 -100 -104754
rect -158 -105542 -146 -104766
rect -112 -105542 -100 -104766
rect -158 -105554 -100 -105542
rect 100 -104766 158 -104754
rect 100 -105542 112 -104766
rect 146 -105542 158 -104766
rect 100 -105554 158 -105542
rect -158 -105802 -100 -105790
rect -158 -106578 -146 -105802
rect -112 -106578 -100 -105802
rect -158 -106590 -100 -106578
rect 100 -105802 158 -105790
rect 100 -106578 112 -105802
rect 146 -106578 158 -105802
rect 100 -106590 158 -106578
rect -158 -106838 -100 -106826
rect -158 -107614 -146 -106838
rect -112 -107614 -100 -106838
rect -158 -107626 -100 -107614
rect 100 -106838 158 -106826
rect 100 -107614 112 -106838
rect 146 -107614 158 -106838
rect 100 -107626 158 -107614
rect -158 -107874 -100 -107862
rect -158 -108650 -146 -107874
rect -112 -108650 -100 -107874
rect -158 -108662 -100 -108650
rect 100 -107874 158 -107862
rect 100 -108650 112 -107874
rect 146 -108650 158 -107874
rect 100 -108662 158 -108650
rect -158 -108910 -100 -108898
rect -158 -109686 -146 -108910
rect -112 -109686 -100 -108910
rect -158 -109698 -100 -109686
rect 100 -108910 158 -108898
rect 100 -109686 112 -108910
rect 146 -109686 158 -108910
rect 100 -109698 158 -109686
rect -158 -109946 -100 -109934
rect -158 -110722 -146 -109946
rect -112 -110722 -100 -109946
rect -158 -110734 -100 -110722
rect 100 -109946 158 -109934
rect 100 -110722 112 -109946
rect 146 -110722 158 -109946
rect 100 -110734 158 -110722
rect -158 -110982 -100 -110970
rect -158 -111758 -146 -110982
rect -112 -111758 -100 -110982
rect -158 -111770 -100 -111758
rect 100 -110982 158 -110970
rect 100 -111758 112 -110982
rect 146 -111758 158 -110982
rect 100 -111770 158 -111758
rect -158 -112018 -100 -112006
rect -158 -112794 -146 -112018
rect -112 -112794 -100 -112018
rect -158 -112806 -100 -112794
rect 100 -112018 158 -112006
rect 100 -112794 112 -112018
rect 146 -112794 158 -112018
rect 100 -112806 158 -112794
rect -158 -113054 -100 -113042
rect -158 -113830 -146 -113054
rect -112 -113830 -100 -113054
rect -158 -113842 -100 -113830
rect 100 -113054 158 -113042
rect 100 -113830 112 -113054
rect 146 -113830 158 -113054
rect 100 -113842 158 -113830
rect -158 -114090 -100 -114078
rect -158 -114866 -146 -114090
rect -112 -114866 -100 -114090
rect -158 -114878 -100 -114866
rect 100 -114090 158 -114078
rect 100 -114866 112 -114090
rect 146 -114866 158 -114090
rect 100 -114878 158 -114866
rect -158 -115126 -100 -115114
rect -158 -115902 -146 -115126
rect -112 -115902 -100 -115126
rect -158 -115914 -100 -115902
rect 100 -115126 158 -115114
rect 100 -115902 112 -115126
rect 146 -115902 158 -115126
rect 100 -115914 158 -115902
rect -158 -116162 -100 -116150
rect -158 -116938 -146 -116162
rect -112 -116938 -100 -116162
rect -158 -116950 -100 -116938
rect 100 -116162 158 -116150
rect 100 -116938 112 -116162
rect 146 -116938 158 -116162
rect 100 -116950 158 -116938
rect -158 -117198 -100 -117186
rect -158 -117974 -146 -117198
rect -112 -117974 -100 -117198
rect -158 -117986 -100 -117974
rect 100 -117198 158 -117186
rect 100 -117974 112 -117198
rect 146 -117974 158 -117198
rect 100 -117986 158 -117974
rect -158 -118234 -100 -118222
rect -158 -119010 -146 -118234
rect -112 -119010 -100 -118234
rect -158 -119022 -100 -119010
rect 100 -118234 158 -118222
rect 100 -119010 112 -118234
rect 146 -119010 158 -118234
rect 100 -119022 158 -119010
rect -158 -119270 -100 -119258
rect -158 -120046 -146 -119270
rect -112 -120046 -100 -119270
rect -158 -120058 -100 -120046
rect 100 -119270 158 -119258
rect 100 -120046 112 -119270
rect 146 -120046 158 -119270
rect 100 -120058 158 -120046
rect -158 -120306 -100 -120294
rect -158 -121082 -146 -120306
rect -112 -121082 -100 -120306
rect -158 -121094 -100 -121082
rect 100 -120306 158 -120294
rect 100 -121082 112 -120306
rect 146 -121082 158 -120306
rect 100 -121094 158 -121082
rect -158 -121342 -100 -121330
rect -158 -122118 -146 -121342
rect -112 -122118 -100 -121342
rect -158 -122130 -100 -122118
rect 100 -121342 158 -121330
rect 100 -122118 112 -121342
rect 146 -122118 158 -121342
rect 100 -122130 158 -122118
rect -158 -122378 -100 -122366
rect -158 -123154 -146 -122378
rect -112 -123154 -100 -122378
rect -158 -123166 -100 -123154
rect 100 -122378 158 -122366
rect 100 -123154 112 -122378
rect 146 -123154 158 -122378
rect 100 -123166 158 -123154
rect -158 -123414 -100 -123402
rect -158 -124190 -146 -123414
rect -112 -124190 -100 -123414
rect -158 -124202 -100 -124190
rect 100 -123414 158 -123402
rect 100 -124190 112 -123414
rect 146 -124190 158 -123414
rect 100 -124202 158 -124190
rect -158 -124450 -100 -124438
rect -158 -125226 -146 -124450
rect -112 -125226 -100 -124450
rect -158 -125238 -100 -125226
rect 100 -124450 158 -124438
rect 100 -125226 112 -124450
rect 146 -125226 158 -124450
rect 100 -125238 158 -125226
rect -158 -125486 -100 -125474
rect -158 -126262 -146 -125486
rect -112 -126262 -100 -125486
rect -158 -126274 -100 -126262
rect 100 -125486 158 -125474
rect 100 -126262 112 -125486
rect 146 -126262 158 -125486
rect 100 -126274 158 -126262
rect -158 -126522 -100 -126510
rect -158 -127298 -146 -126522
rect -112 -127298 -100 -126522
rect -158 -127310 -100 -127298
rect 100 -126522 158 -126510
rect 100 -127298 112 -126522
rect 146 -127298 158 -126522
rect 100 -127310 158 -127298
rect -158 -127558 -100 -127546
rect -158 -128334 -146 -127558
rect -112 -128334 -100 -127558
rect -158 -128346 -100 -128334
rect 100 -127558 158 -127546
rect 100 -128334 112 -127558
rect 146 -128334 158 -127558
rect 100 -128346 158 -128334
rect -158 -128594 -100 -128582
rect -158 -129370 -146 -128594
rect -112 -129370 -100 -128594
rect -158 -129382 -100 -129370
rect 100 -128594 158 -128582
rect 100 -129370 112 -128594
rect 146 -129370 158 -128594
rect 100 -129382 158 -129370
rect -158 -129630 -100 -129618
rect -158 -130406 -146 -129630
rect -112 -130406 -100 -129630
rect -158 -130418 -100 -130406
rect 100 -129630 158 -129618
rect 100 -130406 112 -129630
rect 146 -130406 158 -129630
rect 100 -130418 158 -130406
rect -158 -130666 -100 -130654
rect -158 -131442 -146 -130666
rect -112 -131442 -100 -130666
rect -158 -131454 -100 -131442
rect 100 -130666 158 -130654
rect 100 -131442 112 -130666
rect 146 -131442 158 -130666
rect 100 -131454 158 -131442
rect -158 -131702 -100 -131690
rect -158 -132478 -146 -131702
rect -112 -132478 -100 -131702
rect -158 -132490 -100 -132478
rect 100 -131702 158 -131690
rect 100 -132478 112 -131702
rect 146 -132478 158 -131702
rect 100 -132490 158 -132478
<< mvpdiffc >>
rect -146 131702 -112 132478
rect 112 131702 146 132478
rect -146 130666 -112 131442
rect 112 130666 146 131442
rect -146 129630 -112 130406
rect 112 129630 146 130406
rect -146 128594 -112 129370
rect 112 128594 146 129370
rect -146 127558 -112 128334
rect 112 127558 146 128334
rect -146 126522 -112 127298
rect 112 126522 146 127298
rect -146 125486 -112 126262
rect 112 125486 146 126262
rect -146 124450 -112 125226
rect 112 124450 146 125226
rect -146 123414 -112 124190
rect 112 123414 146 124190
rect -146 122378 -112 123154
rect 112 122378 146 123154
rect -146 121342 -112 122118
rect 112 121342 146 122118
rect -146 120306 -112 121082
rect 112 120306 146 121082
rect -146 119270 -112 120046
rect 112 119270 146 120046
rect -146 118234 -112 119010
rect 112 118234 146 119010
rect -146 117198 -112 117974
rect 112 117198 146 117974
rect -146 116162 -112 116938
rect 112 116162 146 116938
rect -146 115126 -112 115902
rect 112 115126 146 115902
rect -146 114090 -112 114866
rect 112 114090 146 114866
rect -146 113054 -112 113830
rect 112 113054 146 113830
rect -146 112018 -112 112794
rect 112 112018 146 112794
rect -146 110982 -112 111758
rect 112 110982 146 111758
rect -146 109946 -112 110722
rect 112 109946 146 110722
rect -146 108910 -112 109686
rect 112 108910 146 109686
rect -146 107874 -112 108650
rect 112 107874 146 108650
rect -146 106838 -112 107614
rect 112 106838 146 107614
rect -146 105802 -112 106578
rect 112 105802 146 106578
rect -146 104766 -112 105542
rect 112 104766 146 105542
rect -146 103730 -112 104506
rect 112 103730 146 104506
rect -146 102694 -112 103470
rect 112 102694 146 103470
rect -146 101658 -112 102434
rect 112 101658 146 102434
rect -146 100622 -112 101398
rect 112 100622 146 101398
rect -146 99586 -112 100362
rect 112 99586 146 100362
rect -146 98550 -112 99326
rect 112 98550 146 99326
rect -146 97514 -112 98290
rect 112 97514 146 98290
rect -146 96478 -112 97254
rect 112 96478 146 97254
rect -146 95442 -112 96218
rect 112 95442 146 96218
rect -146 94406 -112 95182
rect 112 94406 146 95182
rect -146 93370 -112 94146
rect 112 93370 146 94146
rect -146 92334 -112 93110
rect 112 92334 146 93110
rect -146 91298 -112 92074
rect 112 91298 146 92074
rect -146 90262 -112 91038
rect 112 90262 146 91038
rect -146 89226 -112 90002
rect 112 89226 146 90002
rect -146 88190 -112 88966
rect 112 88190 146 88966
rect -146 87154 -112 87930
rect 112 87154 146 87930
rect -146 86118 -112 86894
rect 112 86118 146 86894
rect -146 85082 -112 85858
rect 112 85082 146 85858
rect -146 84046 -112 84822
rect 112 84046 146 84822
rect -146 83010 -112 83786
rect 112 83010 146 83786
rect -146 81974 -112 82750
rect 112 81974 146 82750
rect -146 80938 -112 81714
rect 112 80938 146 81714
rect -146 79902 -112 80678
rect 112 79902 146 80678
rect -146 78866 -112 79642
rect 112 78866 146 79642
rect -146 77830 -112 78606
rect 112 77830 146 78606
rect -146 76794 -112 77570
rect 112 76794 146 77570
rect -146 75758 -112 76534
rect 112 75758 146 76534
rect -146 74722 -112 75498
rect 112 74722 146 75498
rect -146 73686 -112 74462
rect 112 73686 146 74462
rect -146 72650 -112 73426
rect 112 72650 146 73426
rect -146 71614 -112 72390
rect 112 71614 146 72390
rect -146 70578 -112 71354
rect 112 70578 146 71354
rect -146 69542 -112 70318
rect 112 69542 146 70318
rect -146 68506 -112 69282
rect 112 68506 146 69282
rect -146 67470 -112 68246
rect 112 67470 146 68246
rect -146 66434 -112 67210
rect 112 66434 146 67210
rect -146 65398 -112 66174
rect 112 65398 146 66174
rect -146 64362 -112 65138
rect 112 64362 146 65138
rect -146 63326 -112 64102
rect 112 63326 146 64102
rect -146 62290 -112 63066
rect 112 62290 146 63066
rect -146 61254 -112 62030
rect 112 61254 146 62030
rect -146 60218 -112 60994
rect 112 60218 146 60994
rect -146 59182 -112 59958
rect 112 59182 146 59958
rect -146 58146 -112 58922
rect 112 58146 146 58922
rect -146 57110 -112 57886
rect 112 57110 146 57886
rect -146 56074 -112 56850
rect 112 56074 146 56850
rect -146 55038 -112 55814
rect 112 55038 146 55814
rect -146 54002 -112 54778
rect 112 54002 146 54778
rect -146 52966 -112 53742
rect 112 52966 146 53742
rect -146 51930 -112 52706
rect 112 51930 146 52706
rect -146 50894 -112 51670
rect 112 50894 146 51670
rect -146 49858 -112 50634
rect 112 49858 146 50634
rect -146 48822 -112 49598
rect 112 48822 146 49598
rect -146 47786 -112 48562
rect 112 47786 146 48562
rect -146 46750 -112 47526
rect 112 46750 146 47526
rect -146 45714 -112 46490
rect 112 45714 146 46490
rect -146 44678 -112 45454
rect 112 44678 146 45454
rect -146 43642 -112 44418
rect 112 43642 146 44418
rect -146 42606 -112 43382
rect 112 42606 146 43382
rect -146 41570 -112 42346
rect 112 41570 146 42346
rect -146 40534 -112 41310
rect 112 40534 146 41310
rect -146 39498 -112 40274
rect 112 39498 146 40274
rect -146 38462 -112 39238
rect 112 38462 146 39238
rect -146 37426 -112 38202
rect 112 37426 146 38202
rect -146 36390 -112 37166
rect 112 36390 146 37166
rect -146 35354 -112 36130
rect 112 35354 146 36130
rect -146 34318 -112 35094
rect 112 34318 146 35094
rect -146 33282 -112 34058
rect 112 33282 146 34058
rect -146 32246 -112 33022
rect 112 32246 146 33022
rect -146 31210 -112 31986
rect 112 31210 146 31986
rect -146 30174 -112 30950
rect 112 30174 146 30950
rect -146 29138 -112 29914
rect 112 29138 146 29914
rect -146 28102 -112 28878
rect 112 28102 146 28878
rect -146 27066 -112 27842
rect 112 27066 146 27842
rect -146 26030 -112 26806
rect 112 26030 146 26806
rect -146 24994 -112 25770
rect 112 24994 146 25770
rect -146 23958 -112 24734
rect 112 23958 146 24734
rect -146 22922 -112 23698
rect 112 22922 146 23698
rect -146 21886 -112 22662
rect 112 21886 146 22662
rect -146 20850 -112 21626
rect 112 20850 146 21626
rect -146 19814 -112 20590
rect 112 19814 146 20590
rect -146 18778 -112 19554
rect 112 18778 146 19554
rect -146 17742 -112 18518
rect 112 17742 146 18518
rect -146 16706 -112 17482
rect 112 16706 146 17482
rect -146 15670 -112 16446
rect 112 15670 146 16446
rect -146 14634 -112 15410
rect 112 14634 146 15410
rect -146 13598 -112 14374
rect 112 13598 146 14374
rect -146 12562 -112 13338
rect 112 12562 146 13338
rect -146 11526 -112 12302
rect 112 11526 146 12302
rect -146 10490 -112 11266
rect 112 10490 146 11266
rect -146 9454 -112 10230
rect 112 9454 146 10230
rect -146 8418 -112 9194
rect 112 8418 146 9194
rect -146 7382 -112 8158
rect 112 7382 146 8158
rect -146 6346 -112 7122
rect 112 6346 146 7122
rect -146 5310 -112 6086
rect 112 5310 146 6086
rect -146 4274 -112 5050
rect 112 4274 146 5050
rect -146 3238 -112 4014
rect 112 3238 146 4014
rect -146 2202 -112 2978
rect 112 2202 146 2978
rect -146 1166 -112 1942
rect 112 1166 146 1942
rect -146 130 -112 906
rect 112 130 146 906
rect -146 -906 -112 -130
rect 112 -906 146 -130
rect -146 -1942 -112 -1166
rect 112 -1942 146 -1166
rect -146 -2978 -112 -2202
rect 112 -2978 146 -2202
rect -146 -4014 -112 -3238
rect 112 -4014 146 -3238
rect -146 -5050 -112 -4274
rect 112 -5050 146 -4274
rect -146 -6086 -112 -5310
rect 112 -6086 146 -5310
rect -146 -7122 -112 -6346
rect 112 -7122 146 -6346
rect -146 -8158 -112 -7382
rect 112 -8158 146 -7382
rect -146 -9194 -112 -8418
rect 112 -9194 146 -8418
rect -146 -10230 -112 -9454
rect 112 -10230 146 -9454
rect -146 -11266 -112 -10490
rect 112 -11266 146 -10490
rect -146 -12302 -112 -11526
rect 112 -12302 146 -11526
rect -146 -13338 -112 -12562
rect 112 -13338 146 -12562
rect -146 -14374 -112 -13598
rect 112 -14374 146 -13598
rect -146 -15410 -112 -14634
rect 112 -15410 146 -14634
rect -146 -16446 -112 -15670
rect 112 -16446 146 -15670
rect -146 -17482 -112 -16706
rect 112 -17482 146 -16706
rect -146 -18518 -112 -17742
rect 112 -18518 146 -17742
rect -146 -19554 -112 -18778
rect 112 -19554 146 -18778
rect -146 -20590 -112 -19814
rect 112 -20590 146 -19814
rect -146 -21626 -112 -20850
rect 112 -21626 146 -20850
rect -146 -22662 -112 -21886
rect 112 -22662 146 -21886
rect -146 -23698 -112 -22922
rect 112 -23698 146 -22922
rect -146 -24734 -112 -23958
rect 112 -24734 146 -23958
rect -146 -25770 -112 -24994
rect 112 -25770 146 -24994
rect -146 -26806 -112 -26030
rect 112 -26806 146 -26030
rect -146 -27842 -112 -27066
rect 112 -27842 146 -27066
rect -146 -28878 -112 -28102
rect 112 -28878 146 -28102
rect -146 -29914 -112 -29138
rect 112 -29914 146 -29138
rect -146 -30950 -112 -30174
rect 112 -30950 146 -30174
rect -146 -31986 -112 -31210
rect 112 -31986 146 -31210
rect -146 -33022 -112 -32246
rect 112 -33022 146 -32246
rect -146 -34058 -112 -33282
rect 112 -34058 146 -33282
rect -146 -35094 -112 -34318
rect 112 -35094 146 -34318
rect -146 -36130 -112 -35354
rect 112 -36130 146 -35354
rect -146 -37166 -112 -36390
rect 112 -37166 146 -36390
rect -146 -38202 -112 -37426
rect 112 -38202 146 -37426
rect -146 -39238 -112 -38462
rect 112 -39238 146 -38462
rect -146 -40274 -112 -39498
rect 112 -40274 146 -39498
rect -146 -41310 -112 -40534
rect 112 -41310 146 -40534
rect -146 -42346 -112 -41570
rect 112 -42346 146 -41570
rect -146 -43382 -112 -42606
rect 112 -43382 146 -42606
rect -146 -44418 -112 -43642
rect 112 -44418 146 -43642
rect -146 -45454 -112 -44678
rect 112 -45454 146 -44678
rect -146 -46490 -112 -45714
rect 112 -46490 146 -45714
rect -146 -47526 -112 -46750
rect 112 -47526 146 -46750
rect -146 -48562 -112 -47786
rect 112 -48562 146 -47786
rect -146 -49598 -112 -48822
rect 112 -49598 146 -48822
rect -146 -50634 -112 -49858
rect 112 -50634 146 -49858
rect -146 -51670 -112 -50894
rect 112 -51670 146 -50894
rect -146 -52706 -112 -51930
rect 112 -52706 146 -51930
rect -146 -53742 -112 -52966
rect 112 -53742 146 -52966
rect -146 -54778 -112 -54002
rect 112 -54778 146 -54002
rect -146 -55814 -112 -55038
rect 112 -55814 146 -55038
rect -146 -56850 -112 -56074
rect 112 -56850 146 -56074
rect -146 -57886 -112 -57110
rect 112 -57886 146 -57110
rect -146 -58922 -112 -58146
rect 112 -58922 146 -58146
rect -146 -59958 -112 -59182
rect 112 -59958 146 -59182
rect -146 -60994 -112 -60218
rect 112 -60994 146 -60218
rect -146 -62030 -112 -61254
rect 112 -62030 146 -61254
rect -146 -63066 -112 -62290
rect 112 -63066 146 -62290
rect -146 -64102 -112 -63326
rect 112 -64102 146 -63326
rect -146 -65138 -112 -64362
rect 112 -65138 146 -64362
rect -146 -66174 -112 -65398
rect 112 -66174 146 -65398
rect -146 -67210 -112 -66434
rect 112 -67210 146 -66434
rect -146 -68246 -112 -67470
rect 112 -68246 146 -67470
rect -146 -69282 -112 -68506
rect 112 -69282 146 -68506
rect -146 -70318 -112 -69542
rect 112 -70318 146 -69542
rect -146 -71354 -112 -70578
rect 112 -71354 146 -70578
rect -146 -72390 -112 -71614
rect 112 -72390 146 -71614
rect -146 -73426 -112 -72650
rect 112 -73426 146 -72650
rect -146 -74462 -112 -73686
rect 112 -74462 146 -73686
rect -146 -75498 -112 -74722
rect 112 -75498 146 -74722
rect -146 -76534 -112 -75758
rect 112 -76534 146 -75758
rect -146 -77570 -112 -76794
rect 112 -77570 146 -76794
rect -146 -78606 -112 -77830
rect 112 -78606 146 -77830
rect -146 -79642 -112 -78866
rect 112 -79642 146 -78866
rect -146 -80678 -112 -79902
rect 112 -80678 146 -79902
rect -146 -81714 -112 -80938
rect 112 -81714 146 -80938
rect -146 -82750 -112 -81974
rect 112 -82750 146 -81974
rect -146 -83786 -112 -83010
rect 112 -83786 146 -83010
rect -146 -84822 -112 -84046
rect 112 -84822 146 -84046
rect -146 -85858 -112 -85082
rect 112 -85858 146 -85082
rect -146 -86894 -112 -86118
rect 112 -86894 146 -86118
rect -146 -87930 -112 -87154
rect 112 -87930 146 -87154
rect -146 -88966 -112 -88190
rect 112 -88966 146 -88190
rect -146 -90002 -112 -89226
rect 112 -90002 146 -89226
rect -146 -91038 -112 -90262
rect 112 -91038 146 -90262
rect -146 -92074 -112 -91298
rect 112 -92074 146 -91298
rect -146 -93110 -112 -92334
rect 112 -93110 146 -92334
rect -146 -94146 -112 -93370
rect 112 -94146 146 -93370
rect -146 -95182 -112 -94406
rect 112 -95182 146 -94406
rect -146 -96218 -112 -95442
rect 112 -96218 146 -95442
rect -146 -97254 -112 -96478
rect 112 -97254 146 -96478
rect -146 -98290 -112 -97514
rect 112 -98290 146 -97514
rect -146 -99326 -112 -98550
rect 112 -99326 146 -98550
rect -146 -100362 -112 -99586
rect 112 -100362 146 -99586
rect -146 -101398 -112 -100622
rect 112 -101398 146 -100622
rect -146 -102434 -112 -101658
rect 112 -102434 146 -101658
rect -146 -103470 -112 -102694
rect 112 -103470 146 -102694
rect -146 -104506 -112 -103730
rect 112 -104506 146 -103730
rect -146 -105542 -112 -104766
rect 112 -105542 146 -104766
rect -146 -106578 -112 -105802
rect 112 -106578 146 -105802
rect -146 -107614 -112 -106838
rect 112 -107614 146 -106838
rect -146 -108650 -112 -107874
rect 112 -108650 146 -107874
rect -146 -109686 -112 -108910
rect 112 -109686 146 -108910
rect -146 -110722 -112 -109946
rect 112 -110722 146 -109946
rect -146 -111758 -112 -110982
rect 112 -111758 146 -110982
rect -146 -112794 -112 -112018
rect 112 -112794 146 -112018
rect -146 -113830 -112 -113054
rect 112 -113830 146 -113054
rect -146 -114866 -112 -114090
rect 112 -114866 146 -114090
rect -146 -115902 -112 -115126
rect 112 -115902 146 -115126
rect -146 -116938 -112 -116162
rect 112 -116938 146 -116162
rect -146 -117974 -112 -117198
rect 112 -117974 146 -117198
rect -146 -119010 -112 -118234
rect 112 -119010 146 -118234
rect -146 -120046 -112 -119270
rect 112 -120046 146 -119270
rect -146 -121082 -112 -120306
rect 112 -121082 146 -120306
rect -146 -122118 -112 -121342
rect 112 -122118 146 -121342
rect -146 -123154 -112 -122378
rect 112 -123154 146 -122378
rect -146 -124190 -112 -123414
rect 112 -124190 146 -123414
rect -146 -125226 -112 -124450
rect 112 -125226 146 -124450
rect -146 -126262 -112 -125486
rect 112 -126262 146 -125486
rect -146 -127298 -112 -126522
rect 112 -127298 146 -126522
rect -146 -128334 -112 -127558
rect 112 -128334 146 -127558
rect -146 -129370 -112 -128594
rect 112 -129370 146 -128594
rect -146 -130406 -112 -129630
rect 112 -130406 146 -129630
rect -146 -131442 -112 -130666
rect 112 -131442 146 -130666
rect -146 -132478 -112 -131702
rect 112 -132478 146 -131702
<< mvnsubdiff >>
rect -292 132709 292 132721
rect -292 132675 -184 132709
rect 184 132675 292 132709
rect -292 132663 292 132675
rect -292 132613 -234 132663
rect -292 -132613 -280 132613
rect -246 -132613 -234 132613
rect 234 132613 292 132663
rect -292 -132663 -234 -132613
rect 234 -132613 246 132613
rect 280 -132613 292 132613
rect 234 -132663 292 -132613
rect -292 -132675 292 -132663
rect -292 -132709 -184 -132675
rect 184 -132709 292 -132675
rect -292 -132721 292 -132709
<< mvnsubdiffcont >>
rect -184 132675 184 132709
rect -280 -132613 -246 132613
rect 246 -132613 280 132613
rect -184 -132709 184 -132675
<< poly >>
rect -100 132571 100 132587
rect -100 132537 -84 132571
rect 84 132537 100 132571
rect -100 132490 100 132537
rect -100 131643 100 131690
rect -100 131609 -84 131643
rect 84 131609 100 131643
rect -100 131593 100 131609
rect -100 131535 100 131551
rect -100 131501 -84 131535
rect 84 131501 100 131535
rect -100 131454 100 131501
rect -100 130607 100 130654
rect -100 130573 -84 130607
rect 84 130573 100 130607
rect -100 130557 100 130573
rect -100 130499 100 130515
rect -100 130465 -84 130499
rect 84 130465 100 130499
rect -100 130418 100 130465
rect -100 129571 100 129618
rect -100 129537 -84 129571
rect 84 129537 100 129571
rect -100 129521 100 129537
rect -100 129463 100 129479
rect -100 129429 -84 129463
rect 84 129429 100 129463
rect -100 129382 100 129429
rect -100 128535 100 128582
rect -100 128501 -84 128535
rect 84 128501 100 128535
rect -100 128485 100 128501
rect -100 128427 100 128443
rect -100 128393 -84 128427
rect 84 128393 100 128427
rect -100 128346 100 128393
rect -100 127499 100 127546
rect -100 127465 -84 127499
rect 84 127465 100 127499
rect -100 127449 100 127465
rect -100 127391 100 127407
rect -100 127357 -84 127391
rect 84 127357 100 127391
rect -100 127310 100 127357
rect -100 126463 100 126510
rect -100 126429 -84 126463
rect 84 126429 100 126463
rect -100 126413 100 126429
rect -100 126355 100 126371
rect -100 126321 -84 126355
rect 84 126321 100 126355
rect -100 126274 100 126321
rect -100 125427 100 125474
rect -100 125393 -84 125427
rect 84 125393 100 125427
rect -100 125377 100 125393
rect -100 125319 100 125335
rect -100 125285 -84 125319
rect 84 125285 100 125319
rect -100 125238 100 125285
rect -100 124391 100 124438
rect -100 124357 -84 124391
rect 84 124357 100 124391
rect -100 124341 100 124357
rect -100 124283 100 124299
rect -100 124249 -84 124283
rect 84 124249 100 124283
rect -100 124202 100 124249
rect -100 123355 100 123402
rect -100 123321 -84 123355
rect 84 123321 100 123355
rect -100 123305 100 123321
rect -100 123247 100 123263
rect -100 123213 -84 123247
rect 84 123213 100 123247
rect -100 123166 100 123213
rect -100 122319 100 122366
rect -100 122285 -84 122319
rect 84 122285 100 122319
rect -100 122269 100 122285
rect -100 122211 100 122227
rect -100 122177 -84 122211
rect 84 122177 100 122211
rect -100 122130 100 122177
rect -100 121283 100 121330
rect -100 121249 -84 121283
rect 84 121249 100 121283
rect -100 121233 100 121249
rect -100 121175 100 121191
rect -100 121141 -84 121175
rect 84 121141 100 121175
rect -100 121094 100 121141
rect -100 120247 100 120294
rect -100 120213 -84 120247
rect 84 120213 100 120247
rect -100 120197 100 120213
rect -100 120139 100 120155
rect -100 120105 -84 120139
rect 84 120105 100 120139
rect -100 120058 100 120105
rect -100 119211 100 119258
rect -100 119177 -84 119211
rect 84 119177 100 119211
rect -100 119161 100 119177
rect -100 119103 100 119119
rect -100 119069 -84 119103
rect 84 119069 100 119103
rect -100 119022 100 119069
rect -100 118175 100 118222
rect -100 118141 -84 118175
rect 84 118141 100 118175
rect -100 118125 100 118141
rect -100 118067 100 118083
rect -100 118033 -84 118067
rect 84 118033 100 118067
rect -100 117986 100 118033
rect -100 117139 100 117186
rect -100 117105 -84 117139
rect 84 117105 100 117139
rect -100 117089 100 117105
rect -100 117031 100 117047
rect -100 116997 -84 117031
rect 84 116997 100 117031
rect -100 116950 100 116997
rect -100 116103 100 116150
rect -100 116069 -84 116103
rect 84 116069 100 116103
rect -100 116053 100 116069
rect -100 115995 100 116011
rect -100 115961 -84 115995
rect 84 115961 100 115995
rect -100 115914 100 115961
rect -100 115067 100 115114
rect -100 115033 -84 115067
rect 84 115033 100 115067
rect -100 115017 100 115033
rect -100 114959 100 114975
rect -100 114925 -84 114959
rect 84 114925 100 114959
rect -100 114878 100 114925
rect -100 114031 100 114078
rect -100 113997 -84 114031
rect 84 113997 100 114031
rect -100 113981 100 113997
rect -100 113923 100 113939
rect -100 113889 -84 113923
rect 84 113889 100 113923
rect -100 113842 100 113889
rect -100 112995 100 113042
rect -100 112961 -84 112995
rect 84 112961 100 112995
rect -100 112945 100 112961
rect -100 112887 100 112903
rect -100 112853 -84 112887
rect 84 112853 100 112887
rect -100 112806 100 112853
rect -100 111959 100 112006
rect -100 111925 -84 111959
rect 84 111925 100 111959
rect -100 111909 100 111925
rect -100 111851 100 111867
rect -100 111817 -84 111851
rect 84 111817 100 111851
rect -100 111770 100 111817
rect -100 110923 100 110970
rect -100 110889 -84 110923
rect 84 110889 100 110923
rect -100 110873 100 110889
rect -100 110815 100 110831
rect -100 110781 -84 110815
rect 84 110781 100 110815
rect -100 110734 100 110781
rect -100 109887 100 109934
rect -100 109853 -84 109887
rect 84 109853 100 109887
rect -100 109837 100 109853
rect -100 109779 100 109795
rect -100 109745 -84 109779
rect 84 109745 100 109779
rect -100 109698 100 109745
rect -100 108851 100 108898
rect -100 108817 -84 108851
rect 84 108817 100 108851
rect -100 108801 100 108817
rect -100 108743 100 108759
rect -100 108709 -84 108743
rect 84 108709 100 108743
rect -100 108662 100 108709
rect -100 107815 100 107862
rect -100 107781 -84 107815
rect 84 107781 100 107815
rect -100 107765 100 107781
rect -100 107707 100 107723
rect -100 107673 -84 107707
rect 84 107673 100 107707
rect -100 107626 100 107673
rect -100 106779 100 106826
rect -100 106745 -84 106779
rect 84 106745 100 106779
rect -100 106729 100 106745
rect -100 106671 100 106687
rect -100 106637 -84 106671
rect 84 106637 100 106671
rect -100 106590 100 106637
rect -100 105743 100 105790
rect -100 105709 -84 105743
rect 84 105709 100 105743
rect -100 105693 100 105709
rect -100 105635 100 105651
rect -100 105601 -84 105635
rect 84 105601 100 105635
rect -100 105554 100 105601
rect -100 104707 100 104754
rect -100 104673 -84 104707
rect 84 104673 100 104707
rect -100 104657 100 104673
rect -100 104599 100 104615
rect -100 104565 -84 104599
rect 84 104565 100 104599
rect -100 104518 100 104565
rect -100 103671 100 103718
rect -100 103637 -84 103671
rect 84 103637 100 103671
rect -100 103621 100 103637
rect -100 103563 100 103579
rect -100 103529 -84 103563
rect 84 103529 100 103563
rect -100 103482 100 103529
rect -100 102635 100 102682
rect -100 102601 -84 102635
rect 84 102601 100 102635
rect -100 102585 100 102601
rect -100 102527 100 102543
rect -100 102493 -84 102527
rect 84 102493 100 102527
rect -100 102446 100 102493
rect -100 101599 100 101646
rect -100 101565 -84 101599
rect 84 101565 100 101599
rect -100 101549 100 101565
rect -100 101491 100 101507
rect -100 101457 -84 101491
rect 84 101457 100 101491
rect -100 101410 100 101457
rect -100 100563 100 100610
rect -100 100529 -84 100563
rect 84 100529 100 100563
rect -100 100513 100 100529
rect -100 100455 100 100471
rect -100 100421 -84 100455
rect 84 100421 100 100455
rect -100 100374 100 100421
rect -100 99527 100 99574
rect -100 99493 -84 99527
rect 84 99493 100 99527
rect -100 99477 100 99493
rect -100 99419 100 99435
rect -100 99385 -84 99419
rect 84 99385 100 99419
rect -100 99338 100 99385
rect -100 98491 100 98538
rect -100 98457 -84 98491
rect 84 98457 100 98491
rect -100 98441 100 98457
rect -100 98383 100 98399
rect -100 98349 -84 98383
rect 84 98349 100 98383
rect -100 98302 100 98349
rect -100 97455 100 97502
rect -100 97421 -84 97455
rect 84 97421 100 97455
rect -100 97405 100 97421
rect -100 97347 100 97363
rect -100 97313 -84 97347
rect 84 97313 100 97347
rect -100 97266 100 97313
rect -100 96419 100 96466
rect -100 96385 -84 96419
rect 84 96385 100 96419
rect -100 96369 100 96385
rect -100 96311 100 96327
rect -100 96277 -84 96311
rect 84 96277 100 96311
rect -100 96230 100 96277
rect -100 95383 100 95430
rect -100 95349 -84 95383
rect 84 95349 100 95383
rect -100 95333 100 95349
rect -100 95275 100 95291
rect -100 95241 -84 95275
rect 84 95241 100 95275
rect -100 95194 100 95241
rect -100 94347 100 94394
rect -100 94313 -84 94347
rect 84 94313 100 94347
rect -100 94297 100 94313
rect -100 94239 100 94255
rect -100 94205 -84 94239
rect 84 94205 100 94239
rect -100 94158 100 94205
rect -100 93311 100 93358
rect -100 93277 -84 93311
rect 84 93277 100 93311
rect -100 93261 100 93277
rect -100 93203 100 93219
rect -100 93169 -84 93203
rect 84 93169 100 93203
rect -100 93122 100 93169
rect -100 92275 100 92322
rect -100 92241 -84 92275
rect 84 92241 100 92275
rect -100 92225 100 92241
rect -100 92167 100 92183
rect -100 92133 -84 92167
rect 84 92133 100 92167
rect -100 92086 100 92133
rect -100 91239 100 91286
rect -100 91205 -84 91239
rect 84 91205 100 91239
rect -100 91189 100 91205
rect -100 91131 100 91147
rect -100 91097 -84 91131
rect 84 91097 100 91131
rect -100 91050 100 91097
rect -100 90203 100 90250
rect -100 90169 -84 90203
rect 84 90169 100 90203
rect -100 90153 100 90169
rect -100 90095 100 90111
rect -100 90061 -84 90095
rect 84 90061 100 90095
rect -100 90014 100 90061
rect -100 89167 100 89214
rect -100 89133 -84 89167
rect 84 89133 100 89167
rect -100 89117 100 89133
rect -100 89059 100 89075
rect -100 89025 -84 89059
rect 84 89025 100 89059
rect -100 88978 100 89025
rect -100 88131 100 88178
rect -100 88097 -84 88131
rect 84 88097 100 88131
rect -100 88081 100 88097
rect -100 88023 100 88039
rect -100 87989 -84 88023
rect 84 87989 100 88023
rect -100 87942 100 87989
rect -100 87095 100 87142
rect -100 87061 -84 87095
rect 84 87061 100 87095
rect -100 87045 100 87061
rect -100 86987 100 87003
rect -100 86953 -84 86987
rect 84 86953 100 86987
rect -100 86906 100 86953
rect -100 86059 100 86106
rect -100 86025 -84 86059
rect 84 86025 100 86059
rect -100 86009 100 86025
rect -100 85951 100 85967
rect -100 85917 -84 85951
rect 84 85917 100 85951
rect -100 85870 100 85917
rect -100 85023 100 85070
rect -100 84989 -84 85023
rect 84 84989 100 85023
rect -100 84973 100 84989
rect -100 84915 100 84931
rect -100 84881 -84 84915
rect 84 84881 100 84915
rect -100 84834 100 84881
rect -100 83987 100 84034
rect -100 83953 -84 83987
rect 84 83953 100 83987
rect -100 83937 100 83953
rect -100 83879 100 83895
rect -100 83845 -84 83879
rect 84 83845 100 83879
rect -100 83798 100 83845
rect -100 82951 100 82998
rect -100 82917 -84 82951
rect 84 82917 100 82951
rect -100 82901 100 82917
rect -100 82843 100 82859
rect -100 82809 -84 82843
rect 84 82809 100 82843
rect -100 82762 100 82809
rect -100 81915 100 81962
rect -100 81881 -84 81915
rect 84 81881 100 81915
rect -100 81865 100 81881
rect -100 81807 100 81823
rect -100 81773 -84 81807
rect 84 81773 100 81807
rect -100 81726 100 81773
rect -100 80879 100 80926
rect -100 80845 -84 80879
rect 84 80845 100 80879
rect -100 80829 100 80845
rect -100 80771 100 80787
rect -100 80737 -84 80771
rect 84 80737 100 80771
rect -100 80690 100 80737
rect -100 79843 100 79890
rect -100 79809 -84 79843
rect 84 79809 100 79843
rect -100 79793 100 79809
rect -100 79735 100 79751
rect -100 79701 -84 79735
rect 84 79701 100 79735
rect -100 79654 100 79701
rect -100 78807 100 78854
rect -100 78773 -84 78807
rect 84 78773 100 78807
rect -100 78757 100 78773
rect -100 78699 100 78715
rect -100 78665 -84 78699
rect 84 78665 100 78699
rect -100 78618 100 78665
rect -100 77771 100 77818
rect -100 77737 -84 77771
rect 84 77737 100 77771
rect -100 77721 100 77737
rect -100 77663 100 77679
rect -100 77629 -84 77663
rect 84 77629 100 77663
rect -100 77582 100 77629
rect -100 76735 100 76782
rect -100 76701 -84 76735
rect 84 76701 100 76735
rect -100 76685 100 76701
rect -100 76627 100 76643
rect -100 76593 -84 76627
rect 84 76593 100 76627
rect -100 76546 100 76593
rect -100 75699 100 75746
rect -100 75665 -84 75699
rect 84 75665 100 75699
rect -100 75649 100 75665
rect -100 75591 100 75607
rect -100 75557 -84 75591
rect 84 75557 100 75591
rect -100 75510 100 75557
rect -100 74663 100 74710
rect -100 74629 -84 74663
rect 84 74629 100 74663
rect -100 74613 100 74629
rect -100 74555 100 74571
rect -100 74521 -84 74555
rect 84 74521 100 74555
rect -100 74474 100 74521
rect -100 73627 100 73674
rect -100 73593 -84 73627
rect 84 73593 100 73627
rect -100 73577 100 73593
rect -100 73519 100 73535
rect -100 73485 -84 73519
rect 84 73485 100 73519
rect -100 73438 100 73485
rect -100 72591 100 72638
rect -100 72557 -84 72591
rect 84 72557 100 72591
rect -100 72541 100 72557
rect -100 72483 100 72499
rect -100 72449 -84 72483
rect 84 72449 100 72483
rect -100 72402 100 72449
rect -100 71555 100 71602
rect -100 71521 -84 71555
rect 84 71521 100 71555
rect -100 71505 100 71521
rect -100 71447 100 71463
rect -100 71413 -84 71447
rect 84 71413 100 71447
rect -100 71366 100 71413
rect -100 70519 100 70566
rect -100 70485 -84 70519
rect 84 70485 100 70519
rect -100 70469 100 70485
rect -100 70411 100 70427
rect -100 70377 -84 70411
rect 84 70377 100 70411
rect -100 70330 100 70377
rect -100 69483 100 69530
rect -100 69449 -84 69483
rect 84 69449 100 69483
rect -100 69433 100 69449
rect -100 69375 100 69391
rect -100 69341 -84 69375
rect 84 69341 100 69375
rect -100 69294 100 69341
rect -100 68447 100 68494
rect -100 68413 -84 68447
rect 84 68413 100 68447
rect -100 68397 100 68413
rect -100 68339 100 68355
rect -100 68305 -84 68339
rect 84 68305 100 68339
rect -100 68258 100 68305
rect -100 67411 100 67458
rect -100 67377 -84 67411
rect 84 67377 100 67411
rect -100 67361 100 67377
rect -100 67303 100 67319
rect -100 67269 -84 67303
rect 84 67269 100 67303
rect -100 67222 100 67269
rect -100 66375 100 66422
rect -100 66341 -84 66375
rect 84 66341 100 66375
rect -100 66325 100 66341
rect -100 66267 100 66283
rect -100 66233 -84 66267
rect 84 66233 100 66267
rect -100 66186 100 66233
rect -100 65339 100 65386
rect -100 65305 -84 65339
rect 84 65305 100 65339
rect -100 65289 100 65305
rect -100 65231 100 65247
rect -100 65197 -84 65231
rect 84 65197 100 65231
rect -100 65150 100 65197
rect -100 64303 100 64350
rect -100 64269 -84 64303
rect 84 64269 100 64303
rect -100 64253 100 64269
rect -100 64195 100 64211
rect -100 64161 -84 64195
rect 84 64161 100 64195
rect -100 64114 100 64161
rect -100 63267 100 63314
rect -100 63233 -84 63267
rect 84 63233 100 63267
rect -100 63217 100 63233
rect -100 63159 100 63175
rect -100 63125 -84 63159
rect 84 63125 100 63159
rect -100 63078 100 63125
rect -100 62231 100 62278
rect -100 62197 -84 62231
rect 84 62197 100 62231
rect -100 62181 100 62197
rect -100 62123 100 62139
rect -100 62089 -84 62123
rect 84 62089 100 62123
rect -100 62042 100 62089
rect -100 61195 100 61242
rect -100 61161 -84 61195
rect 84 61161 100 61195
rect -100 61145 100 61161
rect -100 61087 100 61103
rect -100 61053 -84 61087
rect 84 61053 100 61087
rect -100 61006 100 61053
rect -100 60159 100 60206
rect -100 60125 -84 60159
rect 84 60125 100 60159
rect -100 60109 100 60125
rect -100 60051 100 60067
rect -100 60017 -84 60051
rect 84 60017 100 60051
rect -100 59970 100 60017
rect -100 59123 100 59170
rect -100 59089 -84 59123
rect 84 59089 100 59123
rect -100 59073 100 59089
rect -100 59015 100 59031
rect -100 58981 -84 59015
rect 84 58981 100 59015
rect -100 58934 100 58981
rect -100 58087 100 58134
rect -100 58053 -84 58087
rect 84 58053 100 58087
rect -100 58037 100 58053
rect -100 57979 100 57995
rect -100 57945 -84 57979
rect 84 57945 100 57979
rect -100 57898 100 57945
rect -100 57051 100 57098
rect -100 57017 -84 57051
rect 84 57017 100 57051
rect -100 57001 100 57017
rect -100 56943 100 56959
rect -100 56909 -84 56943
rect 84 56909 100 56943
rect -100 56862 100 56909
rect -100 56015 100 56062
rect -100 55981 -84 56015
rect 84 55981 100 56015
rect -100 55965 100 55981
rect -100 55907 100 55923
rect -100 55873 -84 55907
rect 84 55873 100 55907
rect -100 55826 100 55873
rect -100 54979 100 55026
rect -100 54945 -84 54979
rect 84 54945 100 54979
rect -100 54929 100 54945
rect -100 54871 100 54887
rect -100 54837 -84 54871
rect 84 54837 100 54871
rect -100 54790 100 54837
rect -100 53943 100 53990
rect -100 53909 -84 53943
rect 84 53909 100 53943
rect -100 53893 100 53909
rect -100 53835 100 53851
rect -100 53801 -84 53835
rect 84 53801 100 53835
rect -100 53754 100 53801
rect -100 52907 100 52954
rect -100 52873 -84 52907
rect 84 52873 100 52907
rect -100 52857 100 52873
rect -100 52799 100 52815
rect -100 52765 -84 52799
rect 84 52765 100 52799
rect -100 52718 100 52765
rect -100 51871 100 51918
rect -100 51837 -84 51871
rect 84 51837 100 51871
rect -100 51821 100 51837
rect -100 51763 100 51779
rect -100 51729 -84 51763
rect 84 51729 100 51763
rect -100 51682 100 51729
rect -100 50835 100 50882
rect -100 50801 -84 50835
rect 84 50801 100 50835
rect -100 50785 100 50801
rect -100 50727 100 50743
rect -100 50693 -84 50727
rect 84 50693 100 50727
rect -100 50646 100 50693
rect -100 49799 100 49846
rect -100 49765 -84 49799
rect 84 49765 100 49799
rect -100 49749 100 49765
rect -100 49691 100 49707
rect -100 49657 -84 49691
rect 84 49657 100 49691
rect -100 49610 100 49657
rect -100 48763 100 48810
rect -100 48729 -84 48763
rect 84 48729 100 48763
rect -100 48713 100 48729
rect -100 48655 100 48671
rect -100 48621 -84 48655
rect 84 48621 100 48655
rect -100 48574 100 48621
rect -100 47727 100 47774
rect -100 47693 -84 47727
rect 84 47693 100 47727
rect -100 47677 100 47693
rect -100 47619 100 47635
rect -100 47585 -84 47619
rect 84 47585 100 47619
rect -100 47538 100 47585
rect -100 46691 100 46738
rect -100 46657 -84 46691
rect 84 46657 100 46691
rect -100 46641 100 46657
rect -100 46583 100 46599
rect -100 46549 -84 46583
rect 84 46549 100 46583
rect -100 46502 100 46549
rect -100 45655 100 45702
rect -100 45621 -84 45655
rect 84 45621 100 45655
rect -100 45605 100 45621
rect -100 45547 100 45563
rect -100 45513 -84 45547
rect 84 45513 100 45547
rect -100 45466 100 45513
rect -100 44619 100 44666
rect -100 44585 -84 44619
rect 84 44585 100 44619
rect -100 44569 100 44585
rect -100 44511 100 44527
rect -100 44477 -84 44511
rect 84 44477 100 44511
rect -100 44430 100 44477
rect -100 43583 100 43630
rect -100 43549 -84 43583
rect 84 43549 100 43583
rect -100 43533 100 43549
rect -100 43475 100 43491
rect -100 43441 -84 43475
rect 84 43441 100 43475
rect -100 43394 100 43441
rect -100 42547 100 42594
rect -100 42513 -84 42547
rect 84 42513 100 42547
rect -100 42497 100 42513
rect -100 42439 100 42455
rect -100 42405 -84 42439
rect 84 42405 100 42439
rect -100 42358 100 42405
rect -100 41511 100 41558
rect -100 41477 -84 41511
rect 84 41477 100 41511
rect -100 41461 100 41477
rect -100 41403 100 41419
rect -100 41369 -84 41403
rect 84 41369 100 41403
rect -100 41322 100 41369
rect -100 40475 100 40522
rect -100 40441 -84 40475
rect 84 40441 100 40475
rect -100 40425 100 40441
rect -100 40367 100 40383
rect -100 40333 -84 40367
rect 84 40333 100 40367
rect -100 40286 100 40333
rect -100 39439 100 39486
rect -100 39405 -84 39439
rect 84 39405 100 39439
rect -100 39389 100 39405
rect -100 39331 100 39347
rect -100 39297 -84 39331
rect 84 39297 100 39331
rect -100 39250 100 39297
rect -100 38403 100 38450
rect -100 38369 -84 38403
rect 84 38369 100 38403
rect -100 38353 100 38369
rect -100 38295 100 38311
rect -100 38261 -84 38295
rect 84 38261 100 38295
rect -100 38214 100 38261
rect -100 37367 100 37414
rect -100 37333 -84 37367
rect 84 37333 100 37367
rect -100 37317 100 37333
rect -100 37259 100 37275
rect -100 37225 -84 37259
rect 84 37225 100 37259
rect -100 37178 100 37225
rect -100 36331 100 36378
rect -100 36297 -84 36331
rect 84 36297 100 36331
rect -100 36281 100 36297
rect -100 36223 100 36239
rect -100 36189 -84 36223
rect 84 36189 100 36223
rect -100 36142 100 36189
rect -100 35295 100 35342
rect -100 35261 -84 35295
rect 84 35261 100 35295
rect -100 35245 100 35261
rect -100 35187 100 35203
rect -100 35153 -84 35187
rect 84 35153 100 35187
rect -100 35106 100 35153
rect -100 34259 100 34306
rect -100 34225 -84 34259
rect 84 34225 100 34259
rect -100 34209 100 34225
rect -100 34151 100 34167
rect -100 34117 -84 34151
rect 84 34117 100 34151
rect -100 34070 100 34117
rect -100 33223 100 33270
rect -100 33189 -84 33223
rect 84 33189 100 33223
rect -100 33173 100 33189
rect -100 33115 100 33131
rect -100 33081 -84 33115
rect 84 33081 100 33115
rect -100 33034 100 33081
rect -100 32187 100 32234
rect -100 32153 -84 32187
rect 84 32153 100 32187
rect -100 32137 100 32153
rect -100 32079 100 32095
rect -100 32045 -84 32079
rect 84 32045 100 32079
rect -100 31998 100 32045
rect -100 31151 100 31198
rect -100 31117 -84 31151
rect 84 31117 100 31151
rect -100 31101 100 31117
rect -100 31043 100 31059
rect -100 31009 -84 31043
rect 84 31009 100 31043
rect -100 30962 100 31009
rect -100 30115 100 30162
rect -100 30081 -84 30115
rect 84 30081 100 30115
rect -100 30065 100 30081
rect -100 30007 100 30023
rect -100 29973 -84 30007
rect 84 29973 100 30007
rect -100 29926 100 29973
rect -100 29079 100 29126
rect -100 29045 -84 29079
rect 84 29045 100 29079
rect -100 29029 100 29045
rect -100 28971 100 28987
rect -100 28937 -84 28971
rect 84 28937 100 28971
rect -100 28890 100 28937
rect -100 28043 100 28090
rect -100 28009 -84 28043
rect 84 28009 100 28043
rect -100 27993 100 28009
rect -100 27935 100 27951
rect -100 27901 -84 27935
rect 84 27901 100 27935
rect -100 27854 100 27901
rect -100 27007 100 27054
rect -100 26973 -84 27007
rect 84 26973 100 27007
rect -100 26957 100 26973
rect -100 26899 100 26915
rect -100 26865 -84 26899
rect 84 26865 100 26899
rect -100 26818 100 26865
rect -100 25971 100 26018
rect -100 25937 -84 25971
rect 84 25937 100 25971
rect -100 25921 100 25937
rect -100 25863 100 25879
rect -100 25829 -84 25863
rect 84 25829 100 25863
rect -100 25782 100 25829
rect -100 24935 100 24982
rect -100 24901 -84 24935
rect 84 24901 100 24935
rect -100 24885 100 24901
rect -100 24827 100 24843
rect -100 24793 -84 24827
rect 84 24793 100 24827
rect -100 24746 100 24793
rect -100 23899 100 23946
rect -100 23865 -84 23899
rect 84 23865 100 23899
rect -100 23849 100 23865
rect -100 23791 100 23807
rect -100 23757 -84 23791
rect 84 23757 100 23791
rect -100 23710 100 23757
rect -100 22863 100 22910
rect -100 22829 -84 22863
rect 84 22829 100 22863
rect -100 22813 100 22829
rect -100 22755 100 22771
rect -100 22721 -84 22755
rect 84 22721 100 22755
rect -100 22674 100 22721
rect -100 21827 100 21874
rect -100 21793 -84 21827
rect 84 21793 100 21827
rect -100 21777 100 21793
rect -100 21719 100 21735
rect -100 21685 -84 21719
rect 84 21685 100 21719
rect -100 21638 100 21685
rect -100 20791 100 20838
rect -100 20757 -84 20791
rect 84 20757 100 20791
rect -100 20741 100 20757
rect -100 20683 100 20699
rect -100 20649 -84 20683
rect 84 20649 100 20683
rect -100 20602 100 20649
rect -100 19755 100 19802
rect -100 19721 -84 19755
rect 84 19721 100 19755
rect -100 19705 100 19721
rect -100 19647 100 19663
rect -100 19613 -84 19647
rect 84 19613 100 19647
rect -100 19566 100 19613
rect -100 18719 100 18766
rect -100 18685 -84 18719
rect 84 18685 100 18719
rect -100 18669 100 18685
rect -100 18611 100 18627
rect -100 18577 -84 18611
rect 84 18577 100 18611
rect -100 18530 100 18577
rect -100 17683 100 17730
rect -100 17649 -84 17683
rect 84 17649 100 17683
rect -100 17633 100 17649
rect -100 17575 100 17591
rect -100 17541 -84 17575
rect 84 17541 100 17575
rect -100 17494 100 17541
rect -100 16647 100 16694
rect -100 16613 -84 16647
rect 84 16613 100 16647
rect -100 16597 100 16613
rect -100 16539 100 16555
rect -100 16505 -84 16539
rect 84 16505 100 16539
rect -100 16458 100 16505
rect -100 15611 100 15658
rect -100 15577 -84 15611
rect 84 15577 100 15611
rect -100 15561 100 15577
rect -100 15503 100 15519
rect -100 15469 -84 15503
rect 84 15469 100 15503
rect -100 15422 100 15469
rect -100 14575 100 14622
rect -100 14541 -84 14575
rect 84 14541 100 14575
rect -100 14525 100 14541
rect -100 14467 100 14483
rect -100 14433 -84 14467
rect 84 14433 100 14467
rect -100 14386 100 14433
rect -100 13539 100 13586
rect -100 13505 -84 13539
rect 84 13505 100 13539
rect -100 13489 100 13505
rect -100 13431 100 13447
rect -100 13397 -84 13431
rect 84 13397 100 13431
rect -100 13350 100 13397
rect -100 12503 100 12550
rect -100 12469 -84 12503
rect 84 12469 100 12503
rect -100 12453 100 12469
rect -100 12395 100 12411
rect -100 12361 -84 12395
rect 84 12361 100 12395
rect -100 12314 100 12361
rect -100 11467 100 11514
rect -100 11433 -84 11467
rect 84 11433 100 11467
rect -100 11417 100 11433
rect -100 11359 100 11375
rect -100 11325 -84 11359
rect 84 11325 100 11359
rect -100 11278 100 11325
rect -100 10431 100 10478
rect -100 10397 -84 10431
rect 84 10397 100 10431
rect -100 10381 100 10397
rect -100 10323 100 10339
rect -100 10289 -84 10323
rect 84 10289 100 10323
rect -100 10242 100 10289
rect -100 9395 100 9442
rect -100 9361 -84 9395
rect 84 9361 100 9395
rect -100 9345 100 9361
rect -100 9287 100 9303
rect -100 9253 -84 9287
rect 84 9253 100 9287
rect -100 9206 100 9253
rect -100 8359 100 8406
rect -100 8325 -84 8359
rect 84 8325 100 8359
rect -100 8309 100 8325
rect -100 8251 100 8267
rect -100 8217 -84 8251
rect 84 8217 100 8251
rect -100 8170 100 8217
rect -100 7323 100 7370
rect -100 7289 -84 7323
rect 84 7289 100 7323
rect -100 7273 100 7289
rect -100 7215 100 7231
rect -100 7181 -84 7215
rect 84 7181 100 7215
rect -100 7134 100 7181
rect -100 6287 100 6334
rect -100 6253 -84 6287
rect 84 6253 100 6287
rect -100 6237 100 6253
rect -100 6179 100 6195
rect -100 6145 -84 6179
rect 84 6145 100 6179
rect -100 6098 100 6145
rect -100 5251 100 5298
rect -100 5217 -84 5251
rect 84 5217 100 5251
rect -100 5201 100 5217
rect -100 5143 100 5159
rect -100 5109 -84 5143
rect 84 5109 100 5143
rect -100 5062 100 5109
rect -100 4215 100 4262
rect -100 4181 -84 4215
rect 84 4181 100 4215
rect -100 4165 100 4181
rect -100 4107 100 4123
rect -100 4073 -84 4107
rect 84 4073 100 4107
rect -100 4026 100 4073
rect -100 3179 100 3226
rect -100 3145 -84 3179
rect 84 3145 100 3179
rect -100 3129 100 3145
rect -100 3071 100 3087
rect -100 3037 -84 3071
rect 84 3037 100 3071
rect -100 2990 100 3037
rect -100 2143 100 2190
rect -100 2109 -84 2143
rect 84 2109 100 2143
rect -100 2093 100 2109
rect -100 2035 100 2051
rect -100 2001 -84 2035
rect 84 2001 100 2035
rect -100 1954 100 2001
rect -100 1107 100 1154
rect -100 1073 -84 1107
rect 84 1073 100 1107
rect -100 1057 100 1073
rect -100 999 100 1015
rect -100 965 -84 999
rect 84 965 100 999
rect -100 918 100 965
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -965 100 -918
rect -100 -999 -84 -965
rect 84 -999 100 -965
rect -100 -1015 100 -999
rect -100 -1073 100 -1057
rect -100 -1107 -84 -1073
rect 84 -1107 100 -1073
rect -100 -1154 100 -1107
rect -100 -2001 100 -1954
rect -100 -2035 -84 -2001
rect 84 -2035 100 -2001
rect -100 -2051 100 -2035
rect -100 -2109 100 -2093
rect -100 -2143 -84 -2109
rect 84 -2143 100 -2109
rect -100 -2190 100 -2143
rect -100 -3037 100 -2990
rect -100 -3071 -84 -3037
rect 84 -3071 100 -3037
rect -100 -3087 100 -3071
rect -100 -3145 100 -3129
rect -100 -3179 -84 -3145
rect 84 -3179 100 -3145
rect -100 -3226 100 -3179
rect -100 -4073 100 -4026
rect -100 -4107 -84 -4073
rect 84 -4107 100 -4073
rect -100 -4123 100 -4107
rect -100 -4181 100 -4165
rect -100 -4215 -84 -4181
rect 84 -4215 100 -4181
rect -100 -4262 100 -4215
rect -100 -5109 100 -5062
rect -100 -5143 -84 -5109
rect 84 -5143 100 -5109
rect -100 -5159 100 -5143
rect -100 -5217 100 -5201
rect -100 -5251 -84 -5217
rect 84 -5251 100 -5217
rect -100 -5298 100 -5251
rect -100 -6145 100 -6098
rect -100 -6179 -84 -6145
rect 84 -6179 100 -6145
rect -100 -6195 100 -6179
rect -100 -6253 100 -6237
rect -100 -6287 -84 -6253
rect 84 -6287 100 -6253
rect -100 -6334 100 -6287
rect -100 -7181 100 -7134
rect -100 -7215 -84 -7181
rect 84 -7215 100 -7181
rect -100 -7231 100 -7215
rect -100 -7289 100 -7273
rect -100 -7323 -84 -7289
rect 84 -7323 100 -7289
rect -100 -7370 100 -7323
rect -100 -8217 100 -8170
rect -100 -8251 -84 -8217
rect 84 -8251 100 -8217
rect -100 -8267 100 -8251
rect -100 -8325 100 -8309
rect -100 -8359 -84 -8325
rect 84 -8359 100 -8325
rect -100 -8406 100 -8359
rect -100 -9253 100 -9206
rect -100 -9287 -84 -9253
rect 84 -9287 100 -9253
rect -100 -9303 100 -9287
rect -100 -9361 100 -9345
rect -100 -9395 -84 -9361
rect 84 -9395 100 -9361
rect -100 -9442 100 -9395
rect -100 -10289 100 -10242
rect -100 -10323 -84 -10289
rect 84 -10323 100 -10289
rect -100 -10339 100 -10323
rect -100 -10397 100 -10381
rect -100 -10431 -84 -10397
rect 84 -10431 100 -10397
rect -100 -10478 100 -10431
rect -100 -11325 100 -11278
rect -100 -11359 -84 -11325
rect 84 -11359 100 -11325
rect -100 -11375 100 -11359
rect -100 -11433 100 -11417
rect -100 -11467 -84 -11433
rect 84 -11467 100 -11433
rect -100 -11514 100 -11467
rect -100 -12361 100 -12314
rect -100 -12395 -84 -12361
rect 84 -12395 100 -12361
rect -100 -12411 100 -12395
rect -100 -12469 100 -12453
rect -100 -12503 -84 -12469
rect 84 -12503 100 -12469
rect -100 -12550 100 -12503
rect -100 -13397 100 -13350
rect -100 -13431 -84 -13397
rect 84 -13431 100 -13397
rect -100 -13447 100 -13431
rect -100 -13505 100 -13489
rect -100 -13539 -84 -13505
rect 84 -13539 100 -13505
rect -100 -13586 100 -13539
rect -100 -14433 100 -14386
rect -100 -14467 -84 -14433
rect 84 -14467 100 -14433
rect -100 -14483 100 -14467
rect -100 -14541 100 -14525
rect -100 -14575 -84 -14541
rect 84 -14575 100 -14541
rect -100 -14622 100 -14575
rect -100 -15469 100 -15422
rect -100 -15503 -84 -15469
rect 84 -15503 100 -15469
rect -100 -15519 100 -15503
rect -100 -15577 100 -15561
rect -100 -15611 -84 -15577
rect 84 -15611 100 -15577
rect -100 -15658 100 -15611
rect -100 -16505 100 -16458
rect -100 -16539 -84 -16505
rect 84 -16539 100 -16505
rect -100 -16555 100 -16539
rect -100 -16613 100 -16597
rect -100 -16647 -84 -16613
rect 84 -16647 100 -16613
rect -100 -16694 100 -16647
rect -100 -17541 100 -17494
rect -100 -17575 -84 -17541
rect 84 -17575 100 -17541
rect -100 -17591 100 -17575
rect -100 -17649 100 -17633
rect -100 -17683 -84 -17649
rect 84 -17683 100 -17649
rect -100 -17730 100 -17683
rect -100 -18577 100 -18530
rect -100 -18611 -84 -18577
rect 84 -18611 100 -18577
rect -100 -18627 100 -18611
rect -100 -18685 100 -18669
rect -100 -18719 -84 -18685
rect 84 -18719 100 -18685
rect -100 -18766 100 -18719
rect -100 -19613 100 -19566
rect -100 -19647 -84 -19613
rect 84 -19647 100 -19613
rect -100 -19663 100 -19647
rect -100 -19721 100 -19705
rect -100 -19755 -84 -19721
rect 84 -19755 100 -19721
rect -100 -19802 100 -19755
rect -100 -20649 100 -20602
rect -100 -20683 -84 -20649
rect 84 -20683 100 -20649
rect -100 -20699 100 -20683
rect -100 -20757 100 -20741
rect -100 -20791 -84 -20757
rect 84 -20791 100 -20757
rect -100 -20838 100 -20791
rect -100 -21685 100 -21638
rect -100 -21719 -84 -21685
rect 84 -21719 100 -21685
rect -100 -21735 100 -21719
rect -100 -21793 100 -21777
rect -100 -21827 -84 -21793
rect 84 -21827 100 -21793
rect -100 -21874 100 -21827
rect -100 -22721 100 -22674
rect -100 -22755 -84 -22721
rect 84 -22755 100 -22721
rect -100 -22771 100 -22755
rect -100 -22829 100 -22813
rect -100 -22863 -84 -22829
rect 84 -22863 100 -22829
rect -100 -22910 100 -22863
rect -100 -23757 100 -23710
rect -100 -23791 -84 -23757
rect 84 -23791 100 -23757
rect -100 -23807 100 -23791
rect -100 -23865 100 -23849
rect -100 -23899 -84 -23865
rect 84 -23899 100 -23865
rect -100 -23946 100 -23899
rect -100 -24793 100 -24746
rect -100 -24827 -84 -24793
rect 84 -24827 100 -24793
rect -100 -24843 100 -24827
rect -100 -24901 100 -24885
rect -100 -24935 -84 -24901
rect 84 -24935 100 -24901
rect -100 -24982 100 -24935
rect -100 -25829 100 -25782
rect -100 -25863 -84 -25829
rect 84 -25863 100 -25829
rect -100 -25879 100 -25863
rect -100 -25937 100 -25921
rect -100 -25971 -84 -25937
rect 84 -25971 100 -25937
rect -100 -26018 100 -25971
rect -100 -26865 100 -26818
rect -100 -26899 -84 -26865
rect 84 -26899 100 -26865
rect -100 -26915 100 -26899
rect -100 -26973 100 -26957
rect -100 -27007 -84 -26973
rect 84 -27007 100 -26973
rect -100 -27054 100 -27007
rect -100 -27901 100 -27854
rect -100 -27935 -84 -27901
rect 84 -27935 100 -27901
rect -100 -27951 100 -27935
rect -100 -28009 100 -27993
rect -100 -28043 -84 -28009
rect 84 -28043 100 -28009
rect -100 -28090 100 -28043
rect -100 -28937 100 -28890
rect -100 -28971 -84 -28937
rect 84 -28971 100 -28937
rect -100 -28987 100 -28971
rect -100 -29045 100 -29029
rect -100 -29079 -84 -29045
rect 84 -29079 100 -29045
rect -100 -29126 100 -29079
rect -100 -29973 100 -29926
rect -100 -30007 -84 -29973
rect 84 -30007 100 -29973
rect -100 -30023 100 -30007
rect -100 -30081 100 -30065
rect -100 -30115 -84 -30081
rect 84 -30115 100 -30081
rect -100 -30162 100 -30115
rect -100 -31009 100 -30962
rect -100 -31043 -84 -31009
rect 84 -31043 100 -31009
rect -100 -31059 100 -31043
rect -100 -31117 100 -31101
rect -100 -31151 -84 -31117
rect 84 -31151 100 -31117
rect -100 -31198 100 -31151
rect -100 -32045 100 -31998
rect -100 -32079 -84 -32045
rect 84 -32079 100 -32045
rect -100 -32095 100 -32079
rect -100 -32153 100 -32137
rect -100 -32187 -84 -32153
rect 84 -32187 100 -32153
rect -100 -32234 100 -32187
rect -100 -33081 100 -33034
rect -100 -33115 -84 -33081
rect 84 -33115 100 -33081
rect -100 -33131 100 -33115
rect -100 -33189 100 -33173
rect -100 -33223 -84 -33189
rect 84 -33223 100 -33189
rect -100 -33270 100 -33223
rect -100 -34117 100 -34070
rect -100 -34151 -84 -34117
rect 84 -34151 100 -34117
rect -100 -34167 100 -34151
rect -100 -34225 100 -34209
rect -100 -34259 -84 -34225
rect 84 -34259 100 -34225
rect -100 -34306 100 -34259
rect -100 -35153 100 -35106
rect -100 -35187 -84 -35153
rect 84 -35187 100 -35153
rect -100 -35203 100 -35187
rect -100 -35261 100 -35245
rect -100 -35295 -84 -35261
rect 84 -35295 100 -35261
rect -100 -35342 100 -35295
rect -100 -36189 100 -36142
rect -100 -36223 -84 -36189
rect 84 -36223 100 -36189
rect -100 -36239 100 -36223
rect -100 -36297 100 -36281
rect -100 -36331 -84 -36297
rect 84 -36331 100 -36297
rect -100 -36378 100 -36331
rect -100 -37225 100 -37178
rect -100 -37259 -84 -37225
rect 84 -37259 100 -37225
rect -100 -37275 100 -37259
rect -100 -37333 100 -37317
rect -100 -37367 -84 -37333
rect 84 -37367 100 -37333
rect -100 -37414 100 -37367
rect -100 -38261 100 -38214
rect -100 -38295 -84 -38261
rect 84 -38295 100 -38261
rect -100 -38311 100 -38295
rect -100 -38369 100 -38353
rect -100 -38403 -84 -38369
rect 84 -38403 100 -38369
rect -100 -38450 100 -38403
rect -100 -39297 100 -39250
rect -100 -39331 -84 -39297
rect 84 -39331 100 -39297
rect -100 -39347 100 -39331
rect -100 -39405 100 -39389
rect -100 -39439 -84 -39405
rect 84 -39439 100 -39405
rect -100 -39486 100 -39439
rect -100 -40333 100 -40286
rect -100 -40367 -84 -40333
rect 84 -40367 100 -40333
rect -100 -40383 100 -40367
rect -100 -40441 100 -40425
rect -100 -40475 -84 -40441
rect 84 -40475 100 -40441
rect -100 -40522 100 -40475
rect -100 -41369 100 -41322
rect -100 -41403 -84 -41369
rect 84 -41403 100 -41369
rect -100 -41419 100 -41403
rect -100 -41477 100 -41461
rect -100 -41511 -84 -41477
rect 84 -41511 100 -41477
rect -100 -41558 100 -41511
rect -100 -42405 100 -42358
rect -100 -42439 -84 -42405
rect 84 -42439 100 -42405
rect -100 -42455 100 -42439
rect -100 -42513 100 -42497
rect -100 -42547 -84 -42513
rect 84 -42547 100 -42513
rect -100 -42594 100 -42547
rect -100 -43441 100 -43394
rect -100 -43475 -84 -43441
rect 84 -43475 100 -43441
rect -100 -43491 100 -43475
rect -100 -43549 100 -43533
rect -100 -43583 -84 -43549
rect 84 -43583 100 -43549
rect -100 -43630 100 -43583
rect -100 -44477 100 -44430
rect -100 -44511 -84 -44477
rect 84 -44511 100 -44477
rect -100 -44527 100 -44511
rect -100 -44585 100 -44569
rect -100 -44619 -84 -44585
rect 84 -44619 100 -44585
rect -100 -44666 100 -44619
rect -100 -45513 100 -45466
rect -100 -45547 -84 -45513
rect 84 -45547 100 -45513
rect -100 -45563 100 -45547
rect -100 -45621 100 -45605
rect -100 -45655 -84 -45621
rect 84 -45655 100 -45621
rect -100 -45702 100 -45655
rect -100 -46549 100 -46502
rect -100 -46583 -84 -46549
rect 84 -46583 100 -46549
rect -100 -46599 100 -46583
rect -100 -46657 100 -46641
rect -100 -46691 -84 -46657
rect 84 -46691 100 -46657
rect -100 -46738 100 -46691
rect -100 -47585 100 -47538
rect -100 -47619 -84 -47585
rect 84 -47619 100 -47585
rect -100 -47635 100 -47619
rect -100 -47693 100 -47677
rect -100 -47727 -84 -47693
rect 84 -47727 100 -47693
rect -100 -47774 100 -47727
rect -100 -48621 100 -48574
rect -100 -48655 -84 -48621
rect 84 -48655 100 -48621
rect -100 -48671 100 -48655
rect -100 -48729 100 -48713
rect -100 -48763 -84 -48729
rect 84 -48763 100 -48729
rect -100 -48810 100 -48763
rect -100 -49657 100 -49610
rect -100 -49691 -84 -49657
rect 84 -49691 100 -49657
rect -100 -49707 100 -49691
rect -100 -49765 100 -49749
rect -100 -49799 -84 -49765
rect 84 -49799 100 -49765
rect -100 -49846 100 -49799
rect -100 -50693 100 -50646
rect -100 -50727 -84 -50693
rect 84 -50727 100 -50693
rect -100 -50743 100 -50727
rect -100 -50801 100 -50785
rect -100 -50835 -84 -50801
rect 84 -50835 100 -50801
rect -100 -50882 100 -50835
rect -100 -51729 100 -51682
rect -100 -51763 -84 -51729
rect 84 -51763 100 -51729
rect -100 -51779 100 -51763
rect -100 -51837 100 -51821
rect -100 -51871 -84 -51837
rect 84 -51871 100 -51837
rect -100 -51918 100 -51871
rect -100 -52765 100 -52718
rect -100 -52799 -84 -52765
rect 84 -52799 100 -52765
rect -100 -52815 100 -52799
rect -100 -52873 100 -52857
rect -100 -52907 -84 -52873
rect 84 -52907 100 -52873
rect -100 -52954 100 -52907
rect -100 -53801 100 -53754
rect -100 -53835 -84 -53801
rect 84 -53835 100 -53801
rect -100 -53851 100 -53835
rect -100 -53909 100 -53893
rect -100 -53943 -84 -53909
rect 84 -53943 100 -53909
rect -100 -53990 100 -53943
rect -100 -54837 100 -54790
rect -100 -54871 -84 -54837
rect 84 -54871 100 -54837
rect -100 -54887 100 -54871
rect -100 -54945 100 -54929
rect -100 -54979 -84 -54945
rect 84 -54979 100 -54945
rect -100 -55026 100 -54979
rect -100 -55873 100 -55826
rect -100 -55907 -84 -55873
rect 84 -55907 100 -55873
rect -100 -55923 100 -55907
rect -100 -55981 100 -55965
rect -100 -56015 -84 -55981
rect 84 -56015 100 -55981
rect -100 -56062 100 -56015
rect -100 -56909 100 -56862
rect -100 -56943 -84 -56909
rect 84 -56943 100 -56909
rect -100 -56959 100 -56943
rect -100 -57017 100 -57001
rect -100 -57051 -84 -57017
rect 84 -57051 100 -57017
rect -100 -57098 100 -57051
rect -100 -57945 100 -57898
rect -100 -57979 -84 -57945
rect 84 -57979 100 -57945
rect -100 -57995 100 -57979
rect -100 -58053 100 -58037
rect -100 -58087 -84 -58053
rect 84 -58087 100 -58053
rect -100 -58134 100 -58087
rect -100 -58981 100 -58934
rect -100 -59015 -84 -58981
rect 84 -59015 100 -58981
rect -100 -59031 100 -59015
rect -100 -59089 100 -59073
rect -100 -59123 -84 -59089
rect 84 -59123 100 -59089
rect -100 -59170 100 -59123
rect -100 -60017 100 -59970
rect -100 -60051 -84 -60017
rect 84 -60051 100 -60017
rect -100 -60067 100 -60051
rect -100 -60125 100 -60109
rect -100 -60159 -84 -60125
rect 84 -60159 100 -60125
rect -100 -60206 100 -60159
rect -100 -61053 100 -61006
rect -100 -61087 -84 -61053
rect 84 -61087 100 -61053
rect -100 -61103 100 -61087
rect -100 -61161 100 -61145
rect -100 -61195 -84 -61161
rect 84 -61195 100 -61161
rect -100 -61242 100 -61195
rect -100 -62089 100 -62042
rect -100 -62123 -84 -62089
rect 84 -62123 100 -62089
rect -100 -62139 100 -62123
rect -100 -62197 100 -62181
rect -100 -62231 -84 -62197
rect 84 -62231 100 -62197
rect -100 -62278 100 -62231
rect -100 -63125 100 -63078
rect -100 -63159 -84 -63125
rect 84 -63159 100 -63125
rect -100 -63175 100 -63159
rect -100 -63233 100 -63217
rect -100 -63267 -84 -63233
rect 84 -63267 100 -63233
rect -100 -63314 100 -63267
rect -100 -64161 100 -64114
rect -100 -64195 -84 -64161
rect 84 -64195 100 -64161
rect -100 -64211 100 -64195
rect -100 -64269 100 -64253
rect -100 -64303 -84 -64269
rect 84 -64303 100 -64269
rect -100 -64350 100 -64303
rect -100 -65197 100 -65150
rect -100 -65231 -84 -65197
rect 84 -65231 100 -65197
rect -100 -65247 100 -65231
rect -100 -65305 100 -65289
rect -100 -65339 -84 -65305
rect 84 -65339 100 -65305
rect -100 -65386 100 -65339
rect -100 -66233 100 -66186
rect -100 -66267 -84 -66233
rect 84 -66267 100 -66233
rect -100 -66283 100 -66267
rect -100 -66341 100 -66325
rect -100 -66375 -84 -66341
rect 84 -66375 100 -66341
rect -100 -66422 100 -66375
rect -100 -67269 100 -67222
rect -100 -67303 -84 -67269
rect 84 -67303 100 -67269
rect -100 -67319 100 -67303
rect -100 -67377 100 -67361
rect -100 -67411 -84 -67377
rect 84 -67411 100 -67377
rect -100 -67458 100 -67411
rect -100 -68305 100 -68258
rect -100 -68339 -84 -68305
rect 84 -68339 100 -68305
rect -100 -68355 100 -68339
rect -100 -68413 100 -68397
rect -100 -68447 -84 -68413
rect 84 -68447 100 -68413
rect -100 -68494 100 -68447
rect -100 -69341 100 -69294
rect -100 -69375 -84 -69341
rect 84 -69375 100 -69341
rect -100 -69391 100 -69375
rect -100 -69449 100 -69433
rect -100 -69483 -84 -69449
rect 84 -69483 100 -69449
rect -100 -69530 100 -69483
rect -100 -70377 100 -70330
rect -100 -70411 -84 -70377
rect 84 -70411 100 -70377
rect -100 -70427 100 -70411
rect -100 -70485 100 -70469
rect -100 -70519 -84 -70485
rect 84 -70519 100 -70485
rect -100 -70566 100 -70519
rect -100 -71413 100 -71366
rect -100 -71447 -84 -71413
rect 84 -71447 100 -71413
rect -100 -71463 100 -71447
rect -100 -71521 100 -71505
rect -100 -71555 -84 -71521
rect 84 -71555 100 -71521
rect -100 -71602 100 -71555
rect -100 -72449 100 -72402
rect -100 -72483 -84 -72449
rect 84 -72483 100 -72449
rect -100 -72499 100 -72483
rect -100 -72557 100 -72541
rect -100 -72591 -84 -72557
rect 84 -72591 100 -72557
rect -100 -72638 100 -72591
rect -100 -73485 100 -73438
rect -100 -73519 -84 -73485
rect 84 -73519 100 -73485
rect -100 -73535 100 -73519
rect -100 -73593 100 -73577
rect -100 -73627 -84 -73593
rect 84 -73627 100 -73593
rect -100 -73674 100 -73627
rect -100 -74521 100 -74474
rect -100 -74555 -84 -74521
rect 84 -74555 100 -74521
rect -100 -74571 100 -74555
rect -100 -74629 100 -74613
rect -100 -74663 -84 -74629
rect 84 -74663 100 -74629
rect -100 -74710 100 -74663
rect -100 -75557 100 -75510
rect -100 -75591 -84 -75557
rect 84 -75591 100 -75557
rect -100 -75607 100 -75591
rect -100 -75665 100 -75649
rect -100 -75699 -84 -75665
rect 84 -75699 100 -75665
rect -100 -75746 100 -75699
rect -100 -76593 100 -76546
rect -100 -76627 -84 -76593
rect 84 -76627 100 -76593
rect -100 -76643 100 -76627
rect -100 -76701 100 -76685
rect -100 -76735 -84 -76701
rect 84 -76735 100 -76701
rect -100 -76782 100 -76735
rect -100 -77629 100 -77582
rect -100 -77663 -84 -77629
rect 84 -77663 100 -77629
rect -100 -77679 100 -77663
rect -100 -77737 100 -77721
rect -100 -77771 -84 -77737
rect 84 -77771 100 -77737
rect -100 -77818 100 -77771
rect -100 -78665 100 -78618
rect -100 -78699 -84 -78665
rect 84 -78699 100 -78665
rect -100 -78715 100 -78699
rect -100 -78773 100 -78757
rect -100 -78807 -84 -78773
rect 84 -78807 100 -78773
rect -100 -78854 100 -78807
rect -100 -79701 100 -79654
rect -100 -79735 -84 -79701
rect 84 -79735 100 -79701
rect -100 -79751 100 -79735
rect -100 -79809 100 -79793
rect -100 -79843 -84 -79809
rect 84 -79843 100 -79809
rect -100 -79890 100 -79843
rect -100 -80737 100 -80690
rect -100 -80771 -84 -80737
rect 84 -80771 100 -80737
rect -100 -80787 100 -80771
rect -100 -80845 100 -80829
rect -100 -80879 -84 -80845
rect 84 -80879 100 -80845
rect -100 -80926 100 -80879
rect -100 -81773 100 -81726
rect -100 -81807 -84 -81773
rect 84 -81807 100 -81773
rect -100 -81823 100 -81807
rect -100 -81881 100 -81865
rect -100 -81915 -84 -81881
rect 84 -81915 100 -81881
rect -100 -81962 100 -81915
rect -100 -82809 100 -82762
rect -100 -82843 -84 -82809
rect 84 -82843 100 -82809
rect -100 -82859 100 -82843
rect -100 -82917 100 -82901
rect -100 -82951 -84 -82917
rect 84 -82951 100 -82917
rect -100 -82998 100 -82951
rect -100 -83845 100 -83798
rect -100 -83879 -84 -83845
rect 84 -83879 100 -83845
rect -100 -83895 100 -83879
rect -100 -83953 100 -83937
rect -100 -83987 -84 -83953
rect 84 -83987 100 -83953
rect -100 -84034 100 -83987
rect -100 -84881 100 -84834
rect -100 -84915 -84 -84881
rect 84 -84915 100 -84881
rect -100 -84931 100 -84915
rect -100 -84989 100 -84973
rect -100 -85023 -84 -84989
rect 84 -85023 100 -84989
rect -100 -85070 100 -85023
rect -100 -85917 100 -85870
rect -100 -85951 -84 -85917
rect 84 -85951 100 -85917
rect -100 -85967 100 -85951
rect -100 -86025 100 -86009
rect -100 -86059 -84 -86025
rect 84 -86059 100 -86025
rect -100 -86106 100 -86059
rect -100 -86953 100 -86906
rect -100 -86987 -84 -86953
rect 84 -86987 100 -86953
rect -100 -87003 100 -86987
rect -100 -87061 100 -87045
rect -100 -87095 -84 -87061
rect 84 -87095 100 -87061
rect -100 -87142 100 -87095
rect -100 -87989 100 -87942
rect -100 -88023 -84 -87989
rect 84 -88023 100 -87989
rect -100 -88039 100 -88023
rect -100 -88097 100 -88081
rect -100 -88131 -84 -88097
rect 84 -88131 100 -88097
rect -100 -88178 100 -88131
rect -100 -89025 100 -88978
rect -100 -89059 -84 -89025
rect 84 -89059 100 -89025
rect -100 -89075 100 -89059
rect -100 -89133 100 -89117
rect -100 -89167 -84 -89133
rect 84 -89167 100 -89133
rect -100 -89214 100 -89167
rect -100 -90061 100 -90014
rect -100 -90095 -84 -90061
rect 84 -90095 100 -90061
rect -100 -90111 100 -90095
rect -100 -90169 100 -90153
rect -100 -90203 -84 -90169
rect 84 -90203 100 -90169
rect -100 -90250 100 -90203
rect -100 -91097 100 -91050
rect -100 -91131 -84 -91097
rect 84 -91131 100 -91097
rect -100 -91147 100 -91131
rect -100 -91205 100 -91189
rect -100 -91239 -84 -91205
rect 84 -91239 100 -91205
rect -100 -91286 100 -91239
rect -100 -92133 100 -92086
rect -100 -92167 -84 -92133
rect 84 -92167 100 -92133
rect -100 -92183 100 -92167
rect -100 -92241 100 -92225
rect -100 -92275 -84 -92241
rect 84 -92275 100 -92241
rect -100 -92322 100 -92275
rect -100 -93169 100 -93122
rect -100 -93203 -84 -93169
rect 84 -93203 100 -93169
rect -100 -93219 100 -93203
rect -100 -93277 100 -93261
rect -100 -93311 -84 -93277
rect 84 -93311 100 -93277
rect -100 -93358 100 -93311
rect -100 -94205 100 -94158
rect -100 -94239 -84 -94205
rect 84 -94239 100 -94205
rect -100 -94255 100 -94239
rect -100 -94313 100 -94297
rect -100 -94347 -84 -94313
rect 84 -94347 100 -94313
rect -100 -94394 100 -94347
rect -100 -95241 100 -95194
rect -100 -95275 -84 -95241
rect 84 -95275 100 -95241
rect -100 -95291 100 -95275
rect -100 -95349 100 -95333
rect -100 -95383 -84 -95349
rect 84 -95383 100 -95349
rect -100 -95430 100 -95383
rect -100 -96277 100 -96230
rect -100 -96311 -84 -96277
rect 84 -96311 100 -96277
rect -100 -96327 100 -96311
rect -100 -96385 100 -96369
rect -100 -96419 -84 -96385
rect 84 -96419 100 -96385
rect -100 -96466 100 -96419
rect -100 -97313 100 -97266
rect -100 -97347 -84 -97313
rect 84 -97347 100 -97313
rect -100 -97363 100 -97347
rect -100 -97421 100 -97405
rect -100 -97455 -84 -97421
rect 84 -97455 100 -97421
rect -100 -97502 100 -97455
rect -100 -98349 100 -98302
rect -100 -98383 -84 -98349
rect 84 -98383 100 -98349
rect -100 -98399 100 -98383
rect -100 -98457 100 -98441
rect -100 -98491 -84 -98457
rect 84 -98491 100 -98457
rect -100 -98538 100 -98491
rect -100 -99385 100 -99338
rect -100 -99419 -84 -99385
rect 84 -99419 100 -99385
rect -100 -99435 100 -99419
rect -100 -99493 100 -99477
rect -100 -99527 -84 -99493
rect 84 -99527 100 -99493
rect -100 -99574 100 -99527
rect -100 -100421 100 -100374
rect -100 -100455 -84 -100421
rect 84 -100455 100 -100421
rect -100 -100471 100 -100455
rect -100 -100529 100 -100513
rect -100 -100563 -84 -100529
rect 84 -100563 100 -100529
rect -100 -100610 100 -100563
rect -100 -101457 100 -101410
rect -100 -101491 -84 -101457
rect 84 -101491 100 -101457
rect -100 -101507 100 -101491
rect -100 -101565 100 -101549
rect -100 -101599 -84 -101565
rect 84 -101599 100 -101565
rect -100 -101646 100 -101599
rect -100 -102493 100 -102446
rect -100 -102527 -84 -102493
rect 84 -102527 100 -102493
rect -100 -102543 100 -102527
rect -100 -102601 100 -102585
rect -100 -102635 -84 -102601
rect 84 -102635 100 -102601
rect -100 -102682 100 -102635
rect -100 -103529 100 -103482
rect -100 -103563 -84 -103529
rect 84 -103563 100 -103529
rect -100 -103579 100 -103563
rect -100 -103637 100 -103621
rect -100 -103671 -84 -103637
rect 84 -103671 100 -103637
rect -100 -103718 100 -103671
rect -100 -104565 100 -104518
rect -100 -104599 -84 -104565
rect 84 -104599 100 -104565
rect -100 -104615 100 -104599
rect -100 -104673 100 -104657
rect -100 -104707 -84 -104673
rect 84 -104707 100 -104673
rect -100 -104754 100 -104707
rect -100 -105601 100 -105554
rect -100 -105635 -84 -105601
rect 84 -105635 100 -105601
rect -100 -105651 100 -105635
rect -100 -105709 100 -105693
rect -100 -105743 -84 -105709
rect 84 -105743 100 -105709
rect -100 -105790 100 -105743
rect -100 -106637 100 -106590
rect -100 -106671 -84 -106637
rect 84 -106671 100 -106637
rect -100 -106687 100 -106671
rect -100 -106745 100 -106729
rect -100 -106779 -84 -106745
rect 84 -106779 100 -106745
rect -100 -106826 100 -106779
rect -100 -107673 100 -107626
rect -100 -107707 -84 -107673
rect 84 -107707 100 -107673
rect -100 -107723 100 -107707
rect -100 -107781 100 -107765
rect -100 -107815 -84 -107781
rect 84 -107815 100 -107781
rect -100 -107862 100 -107815
rect -100 -108709 100 -108662
rect -100 -108743 -84 -108709
rect 84 -108743 100 -108709
rect -100 -108759 100 -108743
rect -100 -108817 100 -108801
rect -100 -108851 -84 -108817
rect 84 -108851 100 -108817
rect -100 -108898 100 -108851
rect -100 -109745 100 -109698
rect -100 -109779 -84 -109745
rect 84 -109779 100 -109745
rect -100 -109795 100 -109779
rect -100 -109853 100 -109837
rect -100 -109887 -84 -109853
rect 84 -109887 100 -109853
rect -100 -109934 100 -109887
rect -100 -110781 100 -110734
rect -100 -110815 -84 -110781
rect 84 -110815 100 -110781
rect -100 -110831 100 -110815
rect -100 -110889 100 -110873
rect -100 -110923 -84 -110889
rect 84 -110923 100 -110889
rect -100 -110970 100 -110923
rect -100 -111817 100 -111770
rect -100 -111851 -84 -111817
rect 84 -111851 100 -111817
rect -100 -111867 100 -111851
rect -100 -111925 100 -111909
rect -100 -111959 -84 -111925
rect 84 -111959 100 -111925
rect -100 -112006 100 -111959
rect -100 -112853 100 -112806
rect -100 -112887 -84 -112853
rect 84 -112887 100 -112853
rect -100 -112903 100 -112887
rect -100 -112961 100 -112945
rect -100 -112995 -84 -112961
rect 84 -112995 100 -112961
rect -100 -113042 100 -112995
rect -100 -113889 100 -113842
rect -100 -113923 -84 -113889
rect 84 -113923 100 -113889
rect -100 -113939 100 -113923
rect -100 -113997 100 -113981
rect -100 -114031 -84 -113997
rect 84 -114031 100 -113997
rect -100 -114078 100 -114031
rect -100 -114925 100 -114878
rect -100 -114959 -84 -114925
rect 84 -114959 100 -114925
rect -100 -114975 100 -114959
rect -100 -115033 100 -115017
rect -100 -115067 -84 -115033
rect 84 -115067 100 -115033
rect -100 -115114 100 -115067
rect -100 -115961 100 -115914
rect -100 -115995 -84 -115961
rect 84 -115995 100 -115961
rect -100 -116011 100 -115995
rect -100 -116069 100 -116053
rect -100 -116103 -84 -116069
rect 84 -116103 100 -116069
rect -100 -116150 100 -116103
rect -100 -116997 100 -116950
rect -100 -117031 -84 -116997
rect 84 -117031 100 -116997
rect -100 -117047 100 -117031
rect -100 -117105 100 -117089
rect -100 -117139 -84 -117105
rect 84 -117139 100 -117105
rect -100 -117186 100 -117139
rect -100 -118033 100 -117986
rect -100 -118067 -84 -118033
rect 84 -118067 100 -118033
rect -100 -118083 100 -118067
rect -100 -118141 100 -118125
rect -100 -118175 -84 -118141
rect 84 -118175 100 -118141
rect -100 -118222 100 -118175
rect -100 -119069 100 -119022
rect -100 -119103 -84 -119069
rect 84 -119103 100 -119069
rect -100 -119119 100 -119103
rect -100 -119177 100 -119161
rect -100 -119211 -84 -119177
rect 84 -119211 100 -119177
rect -100 -119258 100 -119211
rect -100 -120105 100 -120058
rect -100 -120139 -84 -120105
rect 84 -120139 100 -120105
rect -100 -120155 100 -120139
rect -100 -120213 100 -120197
rect -100 -120247 -84 -120213
rect 84 -120247 100 -120213
rect -100 -120294 100 -120247
rect -100 -121141 100 -121094
rect -100 -121175 -84 -121141
rect 84 -121175 100 -121141
rect -100 -121191 100 -121175
rect -100 -121249 100 -121233
rect -100 -121283 -84 -121249
rect 84 -121283 100 -121249
rect -100 -121330 100 -121283
rect -100 -122177 100 -122130
rect -100 -122211 -84 -122177
rect 84 -122211 100 -122177
rect -100 -122227 100 -122211
rect -100 -122285 100 -122269
rect -100 -122319 -84 -122285
rect 84 -122319 100 -122285
rect -100 -122366 100 -122319
rect -100 -123213 100 -123166
rect -100 -123247 -84 -123213
rect 84 -123247 100 -123213
rect -100 -123263 100 -123247
rect -100 -123321 100 -123305
rect -100 -123355 -84 -123321
rect 84 -123355 100 -123321
rect -100 -123402 100 -123355
rect -100 -124249 100 -124202
rect -100 -124283 -84 -124249
rect 84 -124283 100 -124249
rect -100 -124299 100 -124283
rect -100 -124357 100 -124341
rect -100 -124391 -84 -124357
rect 84 -124391 100 -124357
rect -100 -124438 100 -124391
rect -100 -125285 100 -125238
rect -100 -125319 -84 -125285
rect 84 -125319 100 -125285
rect -100 -125335 100 -125319
rect -100 -125393 100 -125377
rect -100 -125427 -84 -125393
rect 84 -125427 100 -125393
rect -100 -125474 100 -125427
rect -100 -126321 100 -126274
rect -100 -126355 -84 -126321
rect 84 -126355 100 -126321
rect -100 -126371 100 -126355
rect -100 -126429 100 -126413
rect -100 -126463 -84 -126429
rect 84 -126463 100 -126429
rect -100 -126510 100 -126463
rect -100 -127357 100 -127310
rect -100 -127391 -84 -127357
rect 84 -127391 100 -127357
rect -100 -127407 100 -127391
rect -100 -127465 100 -127449
rect -100 -127499 -84 -127465
rect 84 -127499 100 -127465
rect -100 -127546 100 -127499
rect -100 -128393 100 -128346
rect -100 -128427 -84 -128393
rect 84 -128427 100 -128393
rect -100 -128443 100 -128427
rect -100 -128501 100 -128485
rect -100 -128535 -84 -128501
rect 84 -128535 100 -128501
rect -100 -128582 100 -128535
rect -100 -129429 100 -129382
rect -100 -129463 -84 -129429
rect 84 -129463 100 -129429
rect -100 -129479 100 -129463
rect -100 -129537 100 -129521
rect -100 -129571 -84 -129537
rect 84 -129571 100 -129537
rect -100 -129618 100 -129571
rect -100 -130465 100 -130418
rect -100 -130499 -84 -130465
rect 84 -130499 100 -130465
rect -100 -130515 100 -130499
rect -100 -130573 100 -130557
rect -100 -130607 -84 -130573
rect 84 -130607 100 -130573
rect -100 -130654 100 -130607
rect -100 -131501 100 -131454
rect -100 -131535 -84 -131501
rect 84 -131535 100 -131501
rect -100 -131551 100 -131535
rect -100 -131609 100 -131593
rect -100 -131643 -84 -131609
rect 84 -131643 100 -131609
rect -100 -131690 100 -131643
rect -100 -132537 100 -132490
rect -100 -132571 -84 -132537
rect 84 -132571 100 -132537
rect -100 -132587 100 -132571
<< polycont >>
rect -84 132537 84 132571
rect -84 131609 84 131643
rect -84 131501 84 131535
rect -84 130573 84 130607
rect -84 130465 84 130499
rect -84 129537 84 129571
rect -84 129429 84 129463
rect -84 128501 84 128535
rect -84 128393 84 128427
rect -84 127465 84 127499
rect -84 127357 84 127391
rect -84 126429 84 126463
rect -84 126321 84 126355
rect -84 125393 84 125427
rect -84 125285 84 125319
rect -84 124357 84 124391
rect -84 124249 84 124283
rect -84 123321 84 123355
rect -84 123213 84 123247
rect -84 122285 84 122319
rect -84 122177 84 122211
rect -84 121249 84 121283
rect -84 121141 84 121175
rect -84 120213 84 120247
rect -84 120105 84 120139
rect -84 119177 84 119211
rect -84 119069 84 119103
rect -84 118141 84 118175
rect -84 118033 84 118067
rect -84 117105 84 117139
rect -84 116997 84 117031
rect -84 116069 84 116103
rect -84 115961 84 115995
rect -84 115033 84 115067
rect -84 114925 84 114959
rect -84 113997 84 114031
rect -84 113889 84 113923
rect -84 112961 84 112995
rect -84 112853 84 112887
rect -84 111925 84 111959
rect -84 111817 84 111851
rect -84 110889 84 110923
rect -84 110781 84 110815
rect -84 109853 84 109887
rect -84 109745 84 109779
rect -84 108817 84 108851
rect -84 108709 84 108743
rect -84 107781 84 107815
rect -84 107673 84 107707
rect -84 106745 84 106779
rect -84 106637 84 106671
rect -84 105709 84 105743
rect -84 105601 84 105635
rect -84 104673 84 104707
rect -84 104565 84 104599
rect -84 103637 84 103671
rect -84 103529 84 103563
rect -84 102601 84 102635
rect -84 102493 84 102527
rect -84 101565 84 101599
rect -84 101457 84 101491
rect -84 100529 84 100563
rect -84 100421 84 100455
rect -84 99493 84 99527
rect -84 99385 84 99419
rect -84 98457 84 98491
rect -84 98349 84 98383
rect -84 97421 84 97455
rect -84 97313 84 97347
rect -84 96385 84 96419
rect -84 96277 84 96311
rect -84 95349 84 95383
rect -84 95241 84 95275
rect -84 94313 84 94347
rect -84 94205 84 94239
rect -84 93277 84 93311
rect -84 93169 84 93203
rect -84 92241 84 92275
rect -84 92133 84 92167
rect -84 91205 84 91239
rect -84 91097 84 91131
rect -84 90169 84 90203
rect -84 90061 84 90095
rect -84 89133 84 89167
rect -84 89025 84 89059
rect -84 88097 84 88131
rect -84 87989 84 88023
rect -84 87061 84 87095
rect -84 86953 84 86987
rect -84 86025 84 86059
rect -84 85917 84 85951
rect -84 84989 84 85023
rect -84 84881 84 84915
rect -84 83953 84 83987
rect -84 83845 84 83879
rect -84 82917 84 82951
rect -84 82809 84 82843
rect -84 81881 84 81915
rect -84 81773 84 81807
rect -84 80845 84 80879
rect -84 80737 84 80771
rect -84 79809 84 79843
rect -84 79701 84 79735
rect -84 78773 84 78807
rect -84 78665 84 78699
rect -84 77737 84 77771
rect -84 77629 84 77663
rect -84 76701 84 76735
rect -84 76593 84 76627
rect -84 75665 84 75699
rect -84 75557 84 75591
rect -84 74629 84 74663
rect -84 74521 84 74555
rect -84 73593 84 73627
rect -84 73485 84 73519
rect -84 72557 84 72591
rect -84 72449 84 72483
rect -84 71521 84 71555
rect -84 71413 84 71447
rect -84 70485 84 70519
rect -84 70377 84 70411
rect -84 69449 84 69483
rect -84 69341 84 69375
rect -84 68413 84 68447
rect -84 68305 84 68339
rect -84 67377 84 67411
rect -84 67269 84 67303
rect -84 66341 84 66375
rect -84 66233 84 66267
rect -84 65305 84 65339
rect -84 65197 84 65231
rect -84 64269 84 64303
rect -84 64161 84 64195
rect -84 63233 84 63267
rect -84 63125 84 63159
rect -84 62197 84 62231
rect -84 62089 84 62123
rect -84 61161 84 61195
rect -84 61053 84 61087
rect -84 60125 84 60159
rect -84 60017 84 60051
rect -84 59089 84 59123
rect -84 58981 84 59015
rect -84 58053 84 58087
rect -84 57945 84 57979
rect -84 57017 84 57051
rect -84 56909 84 56943
rect -84 55981 84 56015
rect -84 55873 84 55907
rect -84 54945 84 54979
rect -84 54837 84 54871
rect -84 53909 84 53943
rect -84 53801 84 53835
rect -84 52873 84 52907
rect -84 52765 84 52799
rect -84 51837 84 51871
rect -84 51729 84 51763
rect -84 50801 84 50835
rect -84 50693 84 50727
rect -84 49765 84 49799
rect -84 49657 84 49691
rect -84 48729 84 48763
rect -84 48621 84 48655
rect -84 47693 84 47727
rect -84 47585 84 47619
rect -84 46657 84 46691
rect -84 46549 84 46583
rect -84 45621 84 45655
rect -84 45513 84 45547
rect -84 44585 84 44619
rect -84 44477 84 44511
rect -84 43549 84 43583
rect -84 43441 84 43475
rect -84 42513 84 42547
rect -84 42405 84 42439
rect -84 41477 84 41511
rect -84 41369 84 41403
rect -84 40441 84 40475
rect -84 40333 84 40367
rect -84 39405 84 39439
rect -84 39297 84 39331
rect -84 38369 84 38403
rect -84 38261 84 38295
rect -84 37333 84 37367
rect -84 37225 84 37259
rect -84 36297 84 36331
rect -84 36189 84 36223
rect -84 35261 84 35295
rect -84 35153 84 35187
rect -84 34225 84 34259
rect -84 34117 84 34151
rect -84 33189 84 33223
rect -84 33081 84 33115
rect -84 32153 84 32187
rect -84 32045 84 32079
rect -84 31117 84 31151
rect -84 31009 84 31043
rect -84 30081 84 30115
rect -84 29973 84 30007
rect -84 29045 84 29079
rect -84 28937 84 28971
rect -84 28009 84 28043
rect -84 27901 84 27935
rect -84 26973 84 27007
rect -84 26865 84 26899
rect -84 25937 84 25971
rect -84 25829 84 25863
rect -84 24901 84 24935
rect -84 24793 84 24827
rect -84 23865 84 23899
rect -84 23757 84 23791
rect -84 22829 84 22863
rect -84 22721 84 22755
rect -84 21793 84 21827
rect -84 21685 84 21719
rect -84 20757 84 20791
rect -84 20649 84 20683
rect -84 19721 84 19755
rect -84 19613 84 19647
rect -84 18685 84 18719
rect -84 18577 84 18611
rect -84 17649 84 17683
rect -84 17541 84 17575
rect -84 16613 84 16647
rect -84 16505 84 16539
rect -84 15577 84 15611
rect -84 15469 84 15503
rect -84 14541 84 14575
rect -84 14433 84 14467
rect -84 13505 84 13539
rect -84 13397 84 13431
rect -84 12469 84 12503
rect -84 12361 84 12395
rect -84 11433 84 11467
rect -84 11325 84 11359
rect -84 10397 84 10431
rect -84 10289 84 10323
rect -84 9361 84 9395
rect -84 9253 84 9287
rect -84 8325 84 8359
rect -84 8217 84 8251
rect -84 7289 84 7323
rect -84 7181 84 7215
rect -84 6253 84 6287
rect -84 6145 84 6179
rect -84 5217 84 5251
rect -84 5109 84 5143
rect -84 4181 84 4215
rect -84 4073 84 4107
rect -84 3145 84 3179
rect -84 3037 84 3071
rect -84 2109 84 2143
rect -84 2001 84 2035
rect -84 1073 84 1107
rect -84 965 84 999
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -999 84 -965
rect -84 -1107 84 -1073
rect -84 -2035 84 -2001
rect -84 -2143 84 -2109
rect -84 -3071 84 -3037
rect -84 -3179 84 -3145
rect -84 -4107 84 -4073
rect -84 -4215 84 -4181
rect -84 -5143 84 -5109
rect -84 -5251 84 -5217
rect -84 -6179 84 -6145
rect -84 -6287 84 -6253
rect -84 -7215 84 -7181
rect -84 -7323 84 -7289
rect -84 -8251 84 -8217
rect -84 -8359 84 -8325
rect -84 -9287 84 -9253
rect -84 -9395 84 -9361
rect -84 -10323 84 -10289
rect -84 -10431 84 -10397
rect -84 -11359 84 -11325
rect -84 -11467 84 -11433
rect -84 -12395 84 -12361
rect -84 -12503 84 -12469
rect -84 -13431 84 -13397
rect -84 -13539 84 -13505
rect -84 -14467 84 -14433
rect -84 -14575 84 -14541
rect -84 -15503 84 -15469
rect -84 -15611 84 -15577
rect -84 -16539 84 -16505
rect -84 -16647 84 -16613
rect -84 -17575 84 -17541
rect -84 -17683 84 -17649
rect -84 -18611 84 -18577
rect -84 -18719 84 -18685
rect -84 -19647 84 -19613
rect -84 -19755 84 -19721
rect -84 -20683 84 -20649
rect -84 -20791 84 -20757
rect -84 -21719 84 -21685
rect -84 -21827 84 -21793
rect -84 -22755 84 -22721
rect -84 -22863 84 -22829
rect -84 -23791 84 -23757
rect -84 -23899 84 -23865
rect -84 -24827 84 -24793
rect -84 -24935 84 -24901
rect -84 -25863 84 -25829
rect -84 -25971 84 -25937
rect -84 -26899 84 -26865
rect -84 -27007 84 -26973
rect -84 -27935 84 -27901
rect -84 -28043 84 -28009
rect -84 -28971 84 -28937
rect -84 -29079 84 -29045
rect -84 -30007 84 -29973
rect -84 -30115 84 -30081
rect -84 -31043 84 -31009
rect -84 -31151 84 -31117
rect -84 -32079 84 -32045
rect -84 -32187 84 -32153
rect -84 -33115 84 -33081
rect -84 -33223 84 -33189
rect -84 -34151 84 -34117
rect -84 -34259 84 -34225
rect -84 -35187 84 -35153
rect -84 -35295 84 -35261
rect -84 -36223 84 -36189
rect -84 -36331 84 -36297
rect -84 -37259 84 -37225
rect -84 -37367 84 -37333
rect -84 -38295 84 -38261
rect -84 -38403 84 -38369
rect -84 -39331 84 -39297
rect -84 -39439 84 -39405
rect -84 -40367 84 -40333
rect -84 -40475 84 -40441
rect -84 -41403 84 -41369
rect -84 -41511 84 -41477
rect -84 -42439 84 -42405
rect -84 -42547 84 -42513
rect -84 -43475 84 -43441
rect -84 -43583 84 -43549
rect -84 -44511 84 -44477
rect -84 -44619 84 -44585
rect -84 -45547 84 -45513
rect -84 -45655 84 -45621
rect -84 -46583 84 -46549
rect -84 -46691 84 -46657
rect -84 -47619 84 -47585
rect -84 -47727 84 -47693
rect -84 -48655 84 -48621
rect -84 -48763 84 -48729
rect -84 -49691 84 -49657
rect -84 -49799 84 -49765
rect -84 -50727 84 -50693
rect -84 -50835 84 -50801
rect -84 -51763 84 -51729
rect -84 -51871 84 -51837
rect -84 -52799 84 -52765
rect -84 -52907 84 -52873
rect -84 -53835 84 -53801
rect -84 -53943 84 -53909
rect -84 -54871 84 -54837
rect -84 -54979 84 -54945
rect -84 -55907 84 -55873
rect -84 -56015 84 -55981
rect -84 -56943 84 -56909
rect -84 -57051 84 -57017
rect -84 -57979 84 -57945
rect -84 -58087 84 -58053
rect -84 -59015 84 -58981
rect -84 -59123 84 -59089
rect -84 -60051 84 -60017
rect -84 -60159 84 -60125
rect -84 -61087 84 -61053
rect -84 -61195 84 -61161
rect -84 -62123 84 -62089
rect -84 -62231 84 -62197
rect -84 -63159 84 -63125
rect -84 -63267 84 -63233
rect -84 -64195 84 -64161
rect -84 -64303 84 -64269
rect -84 -65231 84 -65197
rect -84 -65339 84 -65305
rect -84 -66267 84 -66233
rect -84 -66375 84 -66341
rect -84 -67303 84 -67269
rect -84 -67411 84 -67377
rect -84 -68339 84 -68305
rect -84 -68447 84 -68413
rect -84 -69375 84 -69341
rect -84 -69483 84 -69449
rect -84 -70411 84 -70377
rect -84 -70519 84 -70485
rect -84 -71447 84 -71413
rect -84 -71555 84 -71521
rect -84 -72483 84 -72449
rect -84 -72591 84 -72557
rect -84 -73519 84 -73485
rect -84 -73627 84 -73593
rect -84 -74555 84 -74521
rect -84 -74663 84 -74629
rect -84 -75591 84 -75557
rect -84 -75699 84 -75665
rect -84 -76627 84 -76593
rect -84 -76735 84 -76701
rect -84 -77663 84 -77629
rect -84 -77771 84 -77737
rect -84 -78699 84 -78665
rect -84 -78807 84 -78773
rect -84 -79735 84 -79701
rect -84 -79843 84 -79809
rect -84 -80771 84 -80737
rect -84 -80879 84 -80845
rect -84 -81807 84 -81773
rect -84 -81915 84 -81881
rect -84 -82843 84 -82809
rect -84 -82951 84 -82917
rect -84 -83879 84 -83845
rect -84 -83987 84 -83953
rect -84 -84915 84 -84881
rect -84 -85023 84 -84989
rect -84 -85951 84 -85917
rect -84 -86059 84 -86025
rect -84 -86987 84 -86953
rect -84 -87095 84 -87061
rect -84 -88023 84 -87989
rect -84 -88131 84 -88097
rect -84 -89059 84 -89025
rect -84 -89167 84 -89133
rect -84 -90095 84 -90061
rect -84 -90203 84 -90169
rect -84 -91131 84 -91097
rect -84 -91239 84 -91205
rect -84 -92167 84 -92133
rect -84 -92275 84 -92241
rect -84 -93203 84 -93169
rect -84 -93311 84 -93277
rect -84 -94239 84 -94205
rect -84 -94347 84 -94313
rect -84 -95275 84 -95241
rect -84 -95383 84 -95349
rect -84 -96311 84 -96277
rect -84 -96419 84 -96385
rect -84 -97347 84 -97313
rect -84 -97455 84 -97421
rect -84 -98383 84 -98349
rect -84 -98491 84 -98457
rect -84 -99419 84 -99385
rect -84 -99527 84 -99493
rect -84 -100455 84 -100421
rect -84 -100563 84 -100529
rect -84 -101491 84 -101457
rect -84 -101599 84 -101565
rect -84 -102527 84 -102493
rect -84 -102635 84 -102601
rect -84 -103563 84 -103529
rect -84 -103671 84 -103637
rect -84 -104599 84 -104565
rect -84 -104707 84 -104673
rect -84 -105635 84 -105601
rect -84 -105743 84 -105709
rect -84 -106671 84 -106637
rect -84 -106779 84 -106745
rect -84 -107707 84 -107673
rect -84 -107815 84 -107781
rect -84 -108743 84 -108709
rect -84 -108851 84 -108817
rect -84 -109779 84 -109745
rect -84 -109887 84 -109853
rect -84 -110815 84 -110781
rect -84 -110923 84 -110889
rect -84 -111851 84 -111817
rect -84 -111959 84 -111925
rect -84 -112887 84 -112853
rect -84 -112995 84 -112961
rect -84 -113923 84 -113889
rect -84 -114031 84 -113997
rect -84 -114959 84 -114925
rect -84 -115067 84 -115033
rect -84 -115995 84 -115961
rect -84 -116103 84 -116069
rect -84 -117031 84 -116997
rect -84 -117139 84 -117105
rect -84 -118067 84 -118033
rect -84 -118175 84 -118141
rect -84 -119103 84 -119069
rect -84 -119211 84 -119177
rect -84 -120139 84 -120105
rect -84 -120247 84 -120213
rect -84 -121175 84 -121141
rect -84 -121283 84 -121249
rect -84 -122211 84 -122177
rect -84 -122319 84 -122285
rect -84 -123247 84 -123213
rect -84 -123355 84 -123321
rect -84 -124283 84 -124249
rect -84 -124391 84 -124357
rect -84 -125319 84 -125285
rect -84 -125427 84 -125393
rect -84 -126355 84 -126321
rect -84 -126463 84 -126429
rect -84 -127391 84 -127357
rect -84 -127499 84 -127465
rect -84 -128427 84 -128393
rect -84 -128535 84 -128501
rect -84 -129463 84 -129429
rect -84 -129571 84 -129537
rect -84 -130499 84 -130465
rect -84 -130607 84 -130573
rect -84 -131535 84 -131501
rect -84 -131643 84 -131609
rect -84 -132571 84 -132537
<< locali >>
rect -280 132675 -184 132709
rect 184 132675 280 132709
rect -280 132613 -246 132675
rect 246 132613 280 132675
rect -100 132537 -84 132571
rect 84 132537 100 132571
rect -146 132478 -112 132494
rect -146 131686 -112 131702
rect 112 132478 146 132494
rect 112 131686 146 131702
rect -100 131609 -84 131643
rect 84 131609 100 131643
rect -100 131501 -84 131535
rect 84 131501 100 131535
rect -146 131442 -112 131458
rect -146 130650 -112 130666
rect 112 131442 146 131458
rect 112 130650 146 130666
rect -100 130573 -84 130607
rect 84 130573 100 130607
rect -100 130465 -84 130499
rect 84 130465 100 130499
rect -146 130406 -112 130422
rect -146 129614 -112 129630
rect 112 130406 146 130422
rect 112 129614 146 129630
rect -100 129537 -84 129571
rect 84 129537 100 129571
rect -100 129429 -84 129463
rect 84 129429 100 129463
rect -146 129370 -112 129386
rect -146 128578 -112 128594
rect 112 129370 146 129386
rect 112 128578 146 128594
rect -100 128501 -84 128535
rect 84 128501 100 128535
rect -100 128393 -84 128427
rect 84 128393 100 128427
rect -146 128334 -112 128350
rect -146 127542 -112 127558
rect 112 128334 146 128350
rect 112 127542 146 127558
rect -100 127465 -84 127499
rect 84 127465 100 127499
rect -100 127357 -84 127391
rect 84 127357 100 127391
rect -146 127298 -112 127314
rect -146 126506 -112 126522
rect 112 127298 146 127314
rect 112 126506 146 126522
rect -100 126429 -84 126463
rect 84 126429 100 126463
rect -100 126321 -84 126355
rect 84 126321 100 126355
rect -146 126262 -112 126278
rect -146 125470 -112 125486
rect 112 126262 146 126278
rect 112 125470 146 125486
rect -100 125393 -84 125427
rect 84 125393 100 125427
rect -100 125285 -84 125319
rect 84 125285 100 125319
rect -146 125226 -112 125242
rect -146 124434 -112 124450
rect 112 125226 146 125242
rect 112 124434 146 124450
rect -100 124357 -84 124391
rect 84 124357 100 124391
rect -100 124249 -84 124283
rect 84 124249 100 124283
rect -146 124190 -112 124206
rect -146 123398 -112 123414
rect 112 124190 146 124206
rect 112 123398 146 123414
rect -100 123321 -84 123355
rect 84 123321 100 123355
rect -100 123213 -84 123247
rect 84 123213 100 123247
rect -146 123154 -112 123170
rect -146 122362 -112 122378
rect 112 123154 146 123170
rect 112 122362 146 122378
rect -100 122285 -84 122319
rect 84 122285 100 122319
rect -100 122177 -84 122211
rect 84 122177 100 122211
rect -146 122118 -112 122134
rect -146 121326 -112 121342
rect 112 122118 146 122134
rect 112 121326 146 121342
rect -100 121249 -84 121283
rect 84 121249 100 121283
rect -100 121141 -84 121175
rect 84 121141 100 121175
rect -146 121082 -112 121098
rect -146 120290 -112 120306
rect 112 121082 146 121098
rect 112 120290 146 120306
rect -100 120213 -84 120247
rect 84 120213 100 120247
rect -100 120105 -84 120139
rect 84 120105 100 120139
rect -146 120046 -112 120062
rect -146 119254 -112 119270
rect 112 120046 146 120062
rect 112 119254 146 119270
rect -100 119177 -84 119211
rect 84 119177 100 119211
rect -100 119069 -84 119103
rect 84 119069 100 119103
rect -146 119010 -112 119026
rect -146 118218 -112 118234
rect 112 119010 146 119026
rect 112 118218 146 118234
rect -100 118141 -84 118175
rect 84 118141 100 118175
rect -100 118033 -84 118067
rect 84 118033 100 118067
rect -146 117974 -112 117990
rect -146 117182 -112 117198
rect 112 117974 146 117990
rect 112 117182 146 117198
rect -100 117105 -84 117139
rect 84 117105 100 117139
rect -100 116997 -84 117031
rect 84 116997 100 117031
rect -146 116938 -112 116954
rect -146 116146 -112 116162
rect 112 116938 146 116954
rect 112 116146 146 116162
rect -100 116069 -84 116103
rect 84 116069 100 116103
rect -100 115961 -84 115995
rect 84 115961 100 115995
rect -146 115902 -112 115918
rect -146 115110 -112 115126
rect 112 115902 146 115918
rect 112 115110 146 115126
rect -100 115033 -84 115067
rect 84 115033 100 115067
rect -100 114925 -84 114959
rect 84 114925 100 114959
rect -146 114866 -112 114882
rect -146 114074 -112 114090
rect 112 114866 146 114882
rect 112 114074 146 114090
rect -100 113997 -84 114031
rect 84 113997 100 114031
rect -100 113889 -84 113923
rect 84 113889 100 113923
rect -146 113830 -112 113846
rect -146 113038 -112 113054
rect 112 113830 146 113846
rect 112 113038 146 113054
rect -100 112961 -84 112995
rect 84 112961 100 112995
rect -100 112853 -84 112887
rect 84 112853 100 112887
rect -146 112794 -112 112810
rect -146 112002 -112 112018
rect 112 112794 146 112810
rect 112 112002 146 112018
rect -100 111925 -84 111959
rect 84 111925 100 111959
rect -100 111817 -84 111851
rect 84 111817 100 111851
rect -146 111758 -112 111774
rect -146 110966 -112 110982
rect 112 111758 146 111774
rect 112 110966 146 110982
rect -100 110889 -84 110923
rect 84 110889 100 110923
rect -100 110781 -84 110815
rect 84 110781 100 110815
rect -146 110722 -112 110738
rect -146 109930 -112 109946
rect 112 110722 146 110738
rect 112 109930 146 109946
rect -100 109853 -84 109887
rect 84 109853 100 109887
rect -100 109745 -84 109779
rect 84 109745 100 109779
rect -146 109686 -112 109702
rect -146 108894 -112 108910
rect 112 109686 146 109702
rect 112 108894 146 108910
rect -100 108817 -84 108851
rect 84 108817 100 108851
rect -100 108709 -84 108743
rect 84 108709 100 108743
rect -146 108650 -112 108666
rect -146 107858 -112 107874
rect 112 108650 146 108666
rect 112 107858 146 107874
rect -100 107781 -84 107815
rect 84 107781 100 107815
rect -100 107673 -84 107707
rect 84 107673 100 107707
rect -146 107614 -112 107630
rect -146 106822 -112 106838
rect 112 107614 146 107630
rect 112 106822 146 106838
rect -100 106745 -84 106779
rect 84 106745 100 106779
rect -100 106637 -84 106671
rect 84 106637 100 106671
rect -146 106578 -112 106594
rect -146 105786 -112 105802
rect 112 106578 146 106594
rect 112 105786 146 105802
rect -100 105709 -84 105743
rect 84 105709 100 105743
rect -100 105601 -84 105635
rect 84 105601 100 105635
rect -146 105542 -112 105558
rect -146 104750 -112 104766
rect 112 105542 146 105558
rect 112 104750 146 104766
rect -100 104673 -84 104707
rect 84 104673 100 104707
rect -100 104565 -84 104599
rect 84 104565 100 104599
rect -146 104506 -112 104522
rect -146 103714 -112 103730
rect 112 104506 146 104522
rect 112 103714 146 103730
rect -100 103637 -84 103671
rect 84 103637 100 103671
rect -100 103529 -84 103563
rect 84 103529 100 103563
rect -146 103470 -112 103486
rect -146 102678 -112 102694
rect 112 103470 146 103486
rect 112 102678 146 102694
rect -100 102601 -84 102635
rect 84 102601 100 102635
rect -100 102493 -84 102527
rect 84 102493 100 102527
rect -146 102434 -112 102450
rect -146 101642 -112 101658
rect 112 102434 146 102450
rect 112 101642 146 101658
rect -100 101565 -84 101599
rect 84 101565 100 101599
rect -100 101457 -84 101491
rect 84 101457 100 101491
rect -146 101398 -112 101414
rect -146 100606 -112 100622
rect 112 101398 146 101414
rect 112 100606 146 100622
rect -100 100529 -84 100563
rect 84 100529 100 100563
rect -100 100421 -84 100455
rect 84 100421 100 100455
rect -146 100362 -112 100378
rect -146 99570 -112 99586
rect 112 100362 146 100378
rect 112 99570 146 99586
rect -100 99493 -84 99527
rect 84 99493 100 99527
rect -100 99385 -84 99419
rect 84 99385 100 99419
rect -146 99326 -112 99342
rect -146 98534 -112 98550
rect 112 99326 146 99342
rect 112 98534 146 98550
rect -100 98457 -84 98491
rect 84 98457 100 98491
rect -100 98349 -84 98383
rect 84 98349 100 98383
rect -146 98290 -112 98306
rect -146 97498 -112 97514
rect 112 98290 146 98306
rect 112 97498 146 97514
rect -100 97421 -84 97455
rect 84 97421 100 97455
rect -100 97313 -84 97347
rect 84 97313 100 97347
rect -146 97254 -112 97270
rect -146 96462 -112 96478
rect 112 97254 146 97270
rect 112 96462 146 96478
rect -100 96385 -84 96419
rect 84 96385 100 96419
rect -100 96277 -84 96311
rect 84 96277 100 96311
rect -146 96218 -112 96234
rect -146 95426 -112 95442
rect 112 96218 146 96234
rect 112 95426 146 95442
rect -100 95349 -84 95383
rect 84 95349 100 95383
rect -100 95241 -84 95275
rect 84 95241 100 95275
rect -146 95182 -112 95198
rect -146 94390 -112 94406
rect 112 95182 146 95198
rect 112 94390 146 94406
rect -100 94313 -84 94347
rect 84 94313 100 94347
rect -100 94205 -84 94239
rect 84 94205 100 94239
rect -146 94146 -112 94162
rect -146 93354 -112 93370
rect 112 94146 146 94162
rect 112 93354 146 93370
rect -100 93277 -84 93311
rect 84 93277 100 93311
rect -100 93169 -84 93203
rect 84 93169 100 93203
rect -146 93110 -112 93126
rect -146 92318 -112 92334
rect 112 93110 146 93126
rect 112 92318 146 92334
rect -100 92241 -84 92275
rect 84 92241 100 92275
rect -100 92133 -84 92167
rect 84 92133 100 92167
rect -146 92074 -112 92090
rect -146 91282 -112 91298
rect 112 92074 146 92090
rect 112 91282 146 91298
rect -100 91205 -84 91239
rect 84 91205 100 91239
rect -100 91097 -84 91131
rect 84 91097 100 91131
rect -146 91038 -112 91054
rect -146 90246 -112 90262
rect 112 91038 146 91054
rect 112 90246 146 90262
rect -100 90169 -84 90203
rect 84 90169 100 90203
rect -100 90061 -84 90095
rect 84 90061 100 90095
rect -146 90002 -112 90018
rect -146 89210 -112 89226
rect 112 90002 146 90018
rect 112 89210 146 89226
rect -100 89133 -84 89167
rect 84 89133 100 89167
rect -100 89025 -84 89059
rect 84 89025 100 89059
rect -146 88966 -112 88982
rect -146 88174 -112 88190
rect 112 88966 146 88982
rect 112 88174 146 88190
rect -100 88097 -84 88131
rect 84 88097 100 88131
rect -100 87989 -84 88023
rect 84 87989 100 88023
rect -146 87930 -112 87946
rect -146 87138 -112 87154
rect 112 87930 146 87946
rect 112 87138 146 87154
rect -100 87061 -84 87095
rect 84 87061 100 87095
rect -100 86953 -84 86987
rect 84 86953 100 86987
rect -146 86894 -112 86910
rect -146 86102 -112 86118
rect 112 86894 146 86910
rect 112 86102 146 86118
rect -100 86025 -84 86059
rect 84 86025 100 86059
rect -100 85917 -84 85951
rect 84 85917 100 85951
rect -146 85858 -112 85874
rect -146 85066 -112 85082
rect 112 85858 146 85874
rect 112 85066 146 85082
rect -100 84989 -84 85023
rect 84 84989 100 85023
rect -100 84881 -84 84915
rect 84 84881 100 84915
rect -146 84822 -112 84838
rect -146 84030 -112 84046
rect 112 84822 146 84838
rect 112 84030 146 84046
rect -100 83953 -84 83987
rect 84 83953 100 83987
rect -100 83845 -84 83879
rect 84 83845 100 83879
rect -146 83786 -112 83802
rect -146 82994 -112 83010
rect 112 83786 146 83802
rect 112 82994 146 83010
rect -100 82917 -84 82951
rect 84 82917 100 82951
rect -100 82809 -84 82843
rect 84 82809 100 82843
rect -146 82750 -112 82766
rect -146 81958 -112 81974
rect 112 82750 146 82766
rect 112 81958 146 81974
rect -100 81881 -84 81915
rect 84 81881 100 81915
rect -100 81773 -84 81807
rect 84 81773 100 81807
rect -146 81714 -112 81730
rect -146 80922 -112 80938
rect 112 81714 146 81730
rect 112 80922 146 80938
rect -100 80845 -84 80879
rect 84 80845 100 80879
rect -100 80737 -84 80771
rect 84 80737 100 80771
rect -146 80678 -112 80694
rect -146 79886 -112 79902
rect 112 80678 146 80694
rect 112 79886 146 79902
rect -100 79809 -84 79843
rect 84 79809 100 79843
rect -100 79701 -84 79735
rect 84 79701 100 79735
rect -146 79642 -112 79658
rect -146 78850 -112 78866
rect 112 79642 146 79658
rect 112 78850 146 78866
rect -100 78773 -84 78807
rect 84 78773 100 78807
rect -100 78665 -84 78699
rect 84 78665 100 78699
rect -146 78606 -112 78622
rect -146 77814 -112 77830
rect 112 78606 146 78622
rect 112 77814 146 77830
rect -100 77737 -84 77771
rect 84 77737 100 77771
rect -100 77629 -84 77663
rect 84 77629 100 77663
rect -146 77570 -112 77586
rect -146 76778 -112 76794
rect 112 77570 146 77586
rect 112 76778 146 76794
rect -100 76701 -84 76735
rect 84 76701 100 76735
rect -100 76593 -84 76627
rect 84 76593 100 76627
rect -146 76534 -112 76550
rect -146 75742 -112 75758
rect 112 76534 146 76550
rect 112 75742 146 75758
rect -100 75665 -84 75699
rect 84 75665 100 75699
rect -100 75557 -84 75591
rect 84 75557 100 75591
rect -146 75498 -112 75514
rect -146 74706 -112 74722
rect 112 75498 146 75514
rect 112 74706 146 74722
rect -100 74629 -84 74663
rect 84 74629 100 74663
rect -100 74521 -84 74555
rect 84 74521 100 74555
rect -146 74462 -112 74478
rect -146 73670 -112 73686
rect 112 74462 146 74478
rect 112 73670 146 73686
rect -100 73593 -84 73627
rect 84 73593 100 73627
rect -100 73485 -84 73519
rect 84 73485 100 73519
rect -146 73426 -112 73442
rect -146 72634 -112 72650
rect 112 73426 146 73442
rect 112 72634 146 72650
rect -100 72557 -84 72591
rect 84 72557 100 72591
rect -100 72449 -84 72483
rect 84 72449 100 72483
rect -146 72390 -112 72406
rect -146 71598 -112 71614
rect 112 72390 146 72406
rect 112 71598 146 71614
rect -100 71521 -84 71555
rect 84 71521 100 71555
rect -100 71413 -84 71447
rect 84 71413 100 71447
rect -146 71354 -112 71370
rect -146 70562 -112 70578
rect 112 71354 146 71370
rect 112 70562 146 70578
rect -100 70485 -84 70519
rect 84 70485 100 70519
rect -100 70377 -84 70411
rect 84 70377 100 70411
rect -146 70318 -112 70334
rect -146 69526 -112 69542
rect 112 70318 146 70334
rect 112 69526 146 69542
rect -100 69449 -84 69483
rect 84 69449 100 69483
rect -100 69341 -84 69375
rect 84 69341 100 69375
rect -146 69282 -112 69298
rect -146 68490 -112 68506
rect 112 69282 146 69298
rect 112 68490 146 68506
rect -100 68413 -84 68447
rect 84 68413 100 68447
rect -100 68305 -84 68339
rect 84 68305 100 68339
rect -146 68246 -112 68262
rect -146 67454 -112 67470
rect 112 68246 146 68262
rect 112 67454 146 67470
rect -100 67377 -84 67411
rect 84 67377 100 67411
rect -100 67269 -84 67303
rect 84 67269 100 67303
rect -146 67210 -112 67226
rect -146 66418 -112 66434
rect 112 67210 146 67226
rect 112 66418 146 66434
rect -100 66341 -84 66375
rect 84 66341 100 66375
rect -100 66233 -84 66267
rect 84 66233 100 66267
rect -146 66174 -112 66190
rect -146 65382 -112 65398
rect 112 66174 146 66190
rect 112 65382 146 65398
rect -100 65305 -84 65339
rect 84 65305 100 65339
rect -100 65197 -84 65231
rect 84 65197 100 65231
rect -146 65138 -112 65154
rect -146 64346 -112 64362
rect 112 65138 146 65154
rect 112 64346 146 64362
rect -100 64269 -84 64303
rect 84 64269 100 64303
rect -100 64161 -84 64195
rect 84 64161 100 64195
rect -146 64102 -112 64118
rect -146 63310 -112 63326
rect 112 64102 146 64118
rect 112 63310 146 63326
rect -100 63233 -84 63267
rect 84 63233 100 63267
rect -100 63125 -84 63159
rect 84 63125 100 63159
rect -146 63066 -112 63082
rect -146 62274 -112 62290
rect 112 63066 146 63082
rect 112 62274 146 62290
rect -100 62197 -84 62231
rect 84 62197 100 62231
rect -100 62089 -84 62123
rect 84 62089 100 62123
rect -146 62030 -112 62046
rect -146 61238 -112 61254
rect 112 62030 146 62046
rect 112 61238 146 61254
rect -100 61161 -84 61195
rect 84 61161 100 61195
rect -100 61053 -84 61087
rect 84 61053 100 61087
rect -146 60994 -112 61010
rect -146 60202 -112 60218
rect 112 60994 146 61010
rect 112 60202 146 60218
rect -100 60125 -84 60159
rect 84 60125 100 60159
rect -100 60017 -84 60051
rect 84 60017 100 60051
rect -146 59958 -112 59974
rect -146 59166 -112 59182
rect 112 59958 146 59974
rect 112 59166 146 59182
rect -100 59089 -84 59123
rect 84 59089 100 59123
rect -100 58981 -84 59015
rect 84 58981 100 59015
rect -146 58922 -112 58938
rect -146 58130 -112 58146
rect 112 58922 146 58938
rect 112 58130 146 58146
rect -100 58053 -84 58087
rect 84 58053 100 58087
rect -100 57945 -84 57979
rect 84 57945 100 57979
rect -146 57886 -112 57902
rect -146 57094 -112 57110
rect 112 57886 146 57902
rect 112 57094 146 57110
rect -100 57017 -84 57051
rect 84 57017 100 57051
rect -100 56909 -84 56943
rect 84 56909 100 56943
rect -146 56850 -112 56866
rect -146 56058 -112 56074
rect 112 56850 146 56866
rect 112 56058 146 56074
rect -100 55981 -84 56015
rect 84 55981 100 56015
rect -100 55873 -84 55907
rect 84 55873 100 55907
rect -146 55814 -112 55830
rect -146 55022 -112 55038
rect 112 55814 146 55830
rect 112 55022 146 55038
rect -100 54945 -84 54979
rect 84 54945 100 54979
rect -100 54837 -84 54871
rect 84 54837 100 54871
rect -146 54778 -112 54794
rect -146 53986 -112 54002
rect 112 54778 146 54794
rect 112 53986 146 54002
rect -100 53909 -84 53943
rect 84 53909 100 53943
rect -100 53801 -84 53835
rect 84 53801 100 53835
rect -146 53742 -112 53758
rect -146 52950 -112 52966
rect 112 53742 146 53758
rect 112 52950 146 52966
rect -100 52873 -84 52907
rect 84 52873 100 52907
rect -100 52765 -84 52799
rect 84 52765 100 52799
rect -146 52706 -112 52722
rect -146 51914 -112 51930
rect 112 52706 146 52722
rect 112 51914 146 51930
rect -100 51837 -84 51871
rect 84 51837 100 51871
rect -100 51729 -84 51763
rect 84 51729 100 51763
rect -146 51670 -112 51686
rect -146 50878 -112 50894
rect 112 51670 146 51686
rect 112 50878 146 50894
rect -100 50801 -84 50835
rect 84 50801 100 50835
rect -100 50693 -84 50727
rect 84 50693 100 50727
rect -146 50634 -112 50650
rect -146 49842 -112 49858
rect 112 50634 146 50650
rect 112 49842 146 49858
rect -100 49765 -84 49799
rect 84 49765 100 49799
rect -100 49657 -84 49691
rect 84 49657 100 49691
rect -146 49598 -112 49614
rect -146 48806 -112 48822
rect 112 49598 146 49614
rect 112 48806 146 48822
rect -100 48729 -84 48763
rect 84 48729 100 48763
rect -100 48621 -84 48655
rect 84 48621 100 48655
rect -146 48562 -112 48578
rect -146 47770 -112 47786
rect 112 48562 146 48578
rect 112 47770 146 47786
rect -100 47693 -84 47727
rect 84 47693 100 47727
rect -100 47585 -84 47619
rect 84 47585 100 47619
rect -146 47526 -112 47542
rect -146 46734 -112 46750
rect 112 47526 146 47542
rect 112 46734 146 46750
rect -100 46657 -84 46691
rect 84 46657 100 46691
rect -100 46549 -84 46583
rect 84 46549 100 46583
rect -146 46490 -112 46506
rect -146 45698 -112 45714
rect 112 46490 146 46506
rect 112 45698 146 45714
rect -100 45621 -84 45655
rect 84 45621 100 45655
rect -100 45513 -84 45547
rect 84 45513 100 45547
rect -146 45454 -112 45470
rect -146 44662 -112 44678
rect 112 45454 146 45470
rect 112 44662 146 44678
rect -100 44585 -84 44619
rect 84 44585 100 44619
rect -100 44477 -84 44511
rect 84 44477 100 44511
rect -146 44418 -112 44434
rect -146 43626 -112 43642
rect 112 44418 146 44434
rect 112 43626 146 43642
rect -100 43549 -84 43583
rect 84 43549 100 43583
rect -100 43441 -84 43475
rect 84 43441 100 43475
rect -146 43382 -112 43398
rect -146 42590 -112 42606
rect 112 43382 146 43398
rect 112 42590 146 42606
rect -100 42513 -84 42547
rect 84 42513 100 42547
rect -100 42405 -84 42439
rect 84 42405 100 42439
rect -146 42346 -112 42362
rect -146 41554 -112 41570
rect 112 42346 146 42362
rect 112 41554 146 41570
rect -100 41477 -84 41511
rect 84 41477 100 41511
rect -100 41369 -84 41403
rect 84 41369 100 41403
rect -146 41310 -112 41326
rect -146 40518 -112 40534
rect 112 41310 146 41326
rect 112 40518 146 40534
rect -100 40441 -84 40475
rect 84 40441 100 40475
rect -100 40333 -84 40367
rect 84 40333 100 40367
rect -146 40274 -112 40290
rect -146 39482 -112 39498
rect 112 40274 146 40290
rect 112 39482 146 39498
rect -100 39405 -84 39439
rect 84 39405 100 39439
rect -100 39297 -84 39331
rect 84 39297 100 39331
rect -146 39238 -112 39254
rect -146 38446 -112 38462
rect 112 39238 146 39254
rect 112 38446 146 38462
rect -100 38369 -84 38403
rect 84 38369 100 38403
rect -100 38261 -84 38295
rect 84 38261 100 38295
rect -146 38202 -112 38218
rect -146 37410 -112 37426
rect 112 38202 146 38218
rect 112 37410 146 37426
rect -100 37333 -84 37367
rect 84 37333 100 37367
rect -100 37225 -84 37259
rect 84 37225 100 37259
rect -146 37166 -112 37182
rect -146 36374 -112 36390
rect 112 37166 146 37182
rect 112 36374 146 36390
rect -100 36297 -84 36331
rect 84 36297 100 36331
rect -100 36189 -84 36223
rect 84 36189 100 36223
rect -146 36130 -112 36146
rect -146 35338 -112 35354
rect 112 36130 146 36146
rect 112 35338 146 35354
rect -100 35261 -84 35295
rect 84 35261 100 35295
rect -100 35153 -84 35187
rect 84 35153 100 35187
rect -146 35094 -112 35110
rect -146 34302 -112 34318
rect 112 35094 146 35110
rect 112 34302 146 34318
rect -100 34225 -84 34259
rect 84 34225 100 34259
rect -100 34117 -84 34151
rect 84 34117 100 34151
rect -146 34058 -112 34074
rect -146 33266 -112 33282
rect 112 34058 146 34074
rect 112 33266 146 33282
rect -100 33189 -84 33223
rect 84 33189 100 33223
rect -100 33081 -84 33115
rect 84 33081 100 33115
rect -146 33022 -112 33038
rect -146 32230 -112 32246
rect 112 33022 146 33038
rect 112 32230 146 32246
rect -100 32153 -84 32187
rect 84 32153 100 32187
rect -100 32045 -84 32079
rect 84 32045 100 32079
rect -146 31986 -112 32002
rect -146 31194 -112 31210
rect 112 31986 146 32002
rect 112 31194 146 31210
rect -100 31117 -84 31151
rect 84 31117 100 31151
rect -100 31009 -84 31043
rect 84 31009 100 31043
rect -146 30950 -112 30966
rect -146 30158 -112 30174
rect 112 30950 146 30966
rect 112 30158 146 30174
rect -100 30081 -84 30115
rect 84 30081 100 30115
rect -100 29973 -84 30007
rect 84 29973 100 30007
rect -146 29914 -112 29930
rect -146 29122 -112 29138
rect 112 29914 146 29930
rect 112 29122 146 29138
rect -100 29045 -84 29079
rect 84 29045 100 29079
rect -100 28937 -84 28971
rect 84 28937 100 28971
rect -146 28878 -112 28894
rect -146 28086 -112 28102
rect 112 28878 146 28894
rect 112 28086 146 28102
rect -100 28009 -84 28043
rect 84 28009 100 28043
rect -100 27901 -84 27935
rect 84 27901 100 27935
rect -146 27842 -112 27858
rect -146 27050 -112 27066
rect 112 27842 146 27858
rect 112 27050 146 27066
rect -100 26973 -84 27007
rect 84 26973 100 27007
rect -100 26865 -84 26899
rect 84 26865 100 26899
rect -146 26806 -112 26822
rect -146 26014 -112 26030
rect 112 26806 146 26822
rect 112 26014 146 26030
rect -100 25937 -84 25971
rect 84 25937 100 25971
rect -100 25829 -84 25863
rect 84 25829 100 25863
rect -146 25770 -112 25786
rect -146 24978 -112 24994
rect 112 25770 146 25786
rect 112 24978 146 24994
rect -100 24901 -84 24935
rect 84 24901 100 24935
rect -100 24793 -84 24827
rect 84 24793 100 24827
rect -146 24734 -112 24750
rect -146 23942 -112 23958
rect 112 24734 146 24750
rect 112 23942 146 23958
rect -100 23865 -84 23899
rect 84 23865 100 23899
rect -100 23757 -84 23791
rect 84 23757 100 23791
rect -146 23698 -112 23714
rect -146 22906 -112 22922
rect 112 23698 146 23714
rect 112 22906 146 22922
rect -100 22829 -84 22863
rect 84 22829 100 22863
rect -100 22721 -84 22755
rect 84 22721 100 22755
rect -146 22662 -112 22678
rect -146 21870 -112 21886
rect 112 22662 146 22678
rect 112 21870 146 21886
rect -100 21793 -84 21827
rect 84 21793 100 21827
rect -100 21685 -84 21719
rect 84 21685 100 21719
rect -146 21626 -112 21642
rect -146 20834 -112 20850
rect 112 21626 146 21642
rect 112 20834 146 20850
rect -100 20757 -84 20791
rect 84 20757 100 20791
rect -100 20649 -84 20683
rect 84 20649 100 20683
rect -146 20590 -112 20606
rect -146 19798 -112 19814
rect 112 20590 146 20606
rect 112 19798 146 19814
rect -100 19721 -84 19755
rect 84 19721 100 19755
rect -100 19613 -84 19647
rect 84 19613 100 19647
rect -146 19554 -112 19570
rect -146 18762 -112 18778
rect 112 19554 146 19570
rect 112 18762 146 18778
rect -100 18685 -84 18719
rect 84 18685 100 18719
rect -100 18577 -84 18611
rect 84 18577 100 18611
rect -146 18518 -112 18534
rect -146 17726 -112 17742
rect 112 18518 146 18534
rect 112 17726 146 17742
rect -100 17649 -84 17683
rect 84 17649 100 17683
rect -100 17541 -84 17575
rect 84 17541 100 17575
rect -146 17482 -112 17498
rect -146 16690 -112 16706
rect 112 17482 146 17498
rect 112 16690 146 16706
rect -100 16613 -84 16647
rect 84 16613 100 16647
rect -100 16505 -84 16539
rect 84 16505 100 16539
rect -146 16446 -112 16462
rect -146 15654 -112 15670
rect 112 16446 146 16462
rect 112 15654 146 15670
rect -100 15577 -84 15611
rect 84 15577 100 15611
rect -100 15469 -84 15503
rect 84 15469 100 15503
rect -146 15410 -112 15426
rect -146 14618 -112 14634
rect 112 15410 146 15426
rect 112 14618 146 14634
rect -100 14541 -84 14575
rect 84 14541 100 14575
rect -100 14433 -84 14467
rect 84 14433 100 14467
rect -146 14374 -112 14390
rect -146 13582 -112 13598
rect 112 14374 146 14390
rect 112 13582 146 13598
rect -100 13505 -84 13539
rect 84 13505 100 13539
rect -100 13397 -84 13431
rect 84 13397 100 13431
rect -146 13338 -112 13354
rect -146 12546 -112 12562
rect 112 13338 146 13354
rect 112 12546 146 12562
rect -100 12469 -84 12503
rect 84 12469 100 12503
rect -100 12361 -84 12395
rect 84 12361 100 12395
rect -146 12302 -112 12318
rect -146 11510 -112 11526
rect 112 12302 146 12318
rect 112 11510 146 11526
rect -100 11433 -84 11467
rect 84 11433 100 11467
rect -100 11325 -84 11359
rect 84 11325 100 11359
rect -146 11266 -112 11282
rect -146 10474 -112 10490
rect 112 11266 146 11282
rect 112 10474 146 10490
rect -100 10397 -84 10431
rect 84 10397 100 10431
rect -100 10289 -84 10323
rect 84 10289 100 10323
rect -146 10230 -112 10246
rect -146 9438 -112 9454
rect 112 10230 146 10246
rect 112 9438 146 9454
rect -100 9361 -84 9395
rect 84 9361 100 9395
rect -100 9253 -84 9287
rect 84 9253 100 9287
rect -146 9194 -112 9210
rect -146 8402 -112 8418
rect 112 9194 146 9210
rect 112 8402 146 8418
rect -100 8325 -84 8359
rect 84 8325 100 8359
rect -100 8217 -84 8251
rect 84 8217 100 8251
rect -146 8158 -112 8174
rect -146 7366 -112 7382
rect 112 8158 146 8174
rect 112 7366 146 7382
rect -100 7289 -84 7323
rect 84 7289 100 7323
rect -100 7181 -84 7215
rect 84 7181 100 7215
rect -146 7122 -112 7138
rect -146 6330 -112 6346
rect 112 7122 146 7138
rect 112 6330 146 6346
rect -100 6253 -84 6287
rect 84 6253 100 6287
rect -100 6145 -84 6179
rect 84 6145 100 6179
rect -146 6086 -112 6102
rect -146 5294 -112 5310
rect 112 6086 146 6102
rect 112 5294 146 5310
rect -100 5217 -84 5251
rect 84 5217 100 5251
rect -100 5109 -84 5143
rect 84 5109 100 5143
rect -146 5050 -112 5066
rect -146 4258 -112 4274
rect 112 5050 146 5066
rect 112 4258 146 4274
rect -100 4181 -84 4215
rect 84 4181 100 4215
rect -100 4073 -84 4107
rect 84 4073 100 4107
rect -146 4014 -112 4030
rect -146 3222 -112 3238
rect 112 4014 146 4030
rect 112 3222 146 3238
rect -100 3145 -84 3179
rect 84 3145 100 3179
rect -100 3037 -84 3071
rect 84 3037 100 3071
rect -146 2978 -112 2994
rect -146 2186 -112 2202
rect 112 2978 146 2994
rect 112 2186 146 2202
rect -100 2109 -84 2143
rect 84 2109 100 2143
rect -100 2001 -84 2035
rect 84 2001 100 2035
rect -146 1942 -112 1958
rect -146 1150 -112 1166
rect 112 1942 146 1958
rect 112 1150 146 1166
rect -100 1073 -84 1107
rect 84 1073 100 1107
rect -100 965 -84 999
rect 84 965 100 999
rect -146 906 -112 922
rect -146 114 -112 130
rect 112 906 146 922
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -922 -112 -906
rect 112 -130 146 -114
rect 112 -922 146 -906
rect -100 -999 -84 -965
rect 84 -999 100 -965
rect -100 -1107 -84 -1073
rect 84 -1107 100 -1073
rect -146 -1166 -112 -1150
rect -146 -1958 -112 -1942
rect 112 -1166 146 -1150
rect 112 -1958 146 -1942
rect -100 -2035 -84 -2001
rect 84 -2035 100 -2001
rect -100 -2143 -84 -2109
rect 84 -2143 100 -2109
rect -146 -2202 -112 -2186
rect -146 -2994 -112 -2978
rect 112 -2202 146 -2186
rect 112 -2994 146 -2978
rect -100 -3071 -84 -3037
rect 84 -3071 100 -3037
rect -100 -3179 -84 -3145
rect 84 -3179 100 -3145
rect -146 -3238 -112 -3222
rect -146 -4030 -112 -4014
rect 112 -3238 146 -3222
rect 112 -4030 146 -4014
rect -100 -4107 -84 -4073
rect 84 -4107 100 -4073
rect -100 -4215 -84 -4181
rect 84 -4215 100 -4181
rect -146 -4274 -112 -4258
rect -146 -5066 -112 -5050
rect 112 -4274 146 -4258
rect 112 -5066 146 -5050
rect -100 -5143 -84 -5109
rect 84 -5143 100 -5109
rect -100 -5251 -84 -5217
rect 84 -5251 100 -5217
rect -146 -5310 -112 -5294
rect -146 -6102 -112 -6086
rect 112 -5310 146 -5294
rect 112 -6102 146 -6086
rect -100 -6179 -84 -6145
rect 84 -6179 100 -6145
rect -100 -6287 -84 -6253
rect 84 -6287 100 -6253
rect -146 -6346 -112 -6330
rect -146 -7138 -112 -7122
rect 112 -6346 146 -6330
rect 112 -7138 146 -7122
rect -100 -7215 -84 -7181
rect 84 -7215 100 -7181
rect -100 -7323 -84 -7289
rect 84 -7323 100 -7289
rect -146 -7382 -112 -7366
rect -146 -8174 -112 -8158
rect 112 -7382 146 -7366
rect 112 -8174 146 -8158
rect -100 -8251 -84 -8217
rect 84 -8251 100 -8217
rect -100 -8359 -84 -8325
rect 84 -8359 100 -8325
rect -146 -8418 -112 -8402
rect -146 -9210 -112 -9194
rect 112 -8418 146 -8402
rect 112 -9210 146 -9194
rect -100 -9287 -84 -9253
rect 84 -9287 100 -9253
rect -100 -9395 -84 -9361
rect 84 -9395 100 -9361
rect -146 -9454 -112 -9438
rect -146 -10246 -112 -10230
rect 112 -9454 146 -9438
rect 112 -10246 146 -10230
rect -100 -10323 -84 -10289
rect 84 -10323 100 -10289
rect -100 -10431 -84 -10397
rect 84 -10431 100 -10397
rect -146 -10490 -112 -10474
rect -146 -11282 -112 -11266
rect 112 -10490 146 -10474
rect 112 -11282 146 -11266
rect -100 -11359 -84 -11325
rect 84 -11359 100 -11325
rect -100 -11467 -84 -11433
rect 84 -11467 100 -11433
rect -146 -11526 -112 -11510
rect -146 -12318 -112 -12302
rect 112 -11526 146 -11510
rect 112 -12318 146 -12302
rect -100 -12395 -84 -12361
rect 84 -12395 100 -12361
rect -100 -12503 -84 -12469
rect 84 -12503 100 -12469
rect -146 -12562 -112 -12546
rect -146 -13354 -112 -13338
rect 112 -12562 146 -12546
rect 112 -13354 146 -13338
rect -100 -13431 -84 -13397
rect 84 -13431 100 -13397
rect -100 -13539 -84 -13505
rect 84 -13539 100 -13505
rect -146 -13598 -112 -13582
rect -146 -14390 -112 -14374
rect 112 -13598 146 -13582
rect 112 -14390 146 -14374
rect -100 -14467 -84 -14433
rect 84 -14467 100 -14433
rect -100 -14575 -84 -14541
rect 84 -14575 100 -14541
rect -146 -14634 -112 -14618
rect -146 -15426 -112 -15410
rect 112 -14634 146 -14618
rect 112 -15426 146 -15410
rect -100 -15503 -84 -15469
rect 84 -15503 100 -15469
rect -100 -15611 -84 -15577
rect 84 -15611 100 -15577
rect -146 -15670 -112 -15654
rect -146 -16462 -112 -16446
rect 112 -15670 146 -15654
rect 112 -16462 146 -16446
rect -100 -16539 -84 -16505
rect 84 -16539 100 -16505
rect -100 -16647 -84 -16613
rect 84 -16647 100 -16613
rect -146 -16706 -112 -16690
rect -146 -17498 -112 -17482
rect 112 -16706 146 -16690
rect 112 -17498 146 -17482
rect -100 -17575 -84 -17541
rect 84 -17575 100 -17541
rect -100 -17683 -84 -17649
rect 84 -17683 100 -17649
rect -146 -17742 -112 -17726
rect -146 -18534 -112 -18518
rect 112 -17742 146 -17726
rect 112 -18534 146 -18518
rect -100 -18611 -84 -18577
rect 84 -18611 100 -18577
rect -100 -18719 -84 -18685
rect 84 -18719 100 -18685
rect -146 -18778 -112 -18762
rect -146 -19570 -112 -19554
rect 112 -18778 146 -18762
rect 112 -19570 146 -19554
rect -100 -19647 -84 -19613
rect 84 -19647 100 -19613
rect -100 -19755 -84 -19721
rect 84 -19755 100 -19721
rect -146 -19814 -112 -19798
rect -146 -20606 -112 -20590
rect 112 -19814 146 -19798
rect 112 -20606 146 -20590
rect -100 -20683 -84 -20649
rect 84 -20683 100 -20649
rect -100 -20791 -84 -20757
rect 84 -20791 100 -20757
rect -146 -20850 -112 -20834
rect -146 -21642 -112 -21626
rect 112 -20850 146 -20834
rect 112 -21642 146 -21626
rect -100 -21719 -84 -21685
rect 84 -21719 100 -21685
rect -100 -21827 -84 -21793
rect 84 -21827 100 -21793
rect -146 -21886 -112 -21870
rect -146 -22678 -112 -22662
rect 112 -21886 146 -21870
rect 112 -22678 146 -22662
rect -100 -22755 -84 -22721
rect 84 -22755 100 -22721
rect -100 -22863 -84 -22829
rect 84 -22863 100 -22829
rect -146 -22922 -112 -22906
rect -146 -23714 -112 -23698
rect 112 -22922 146 -22906
rect 112 -23714 146 -23698
rect -100 -23791 -84 -23757
rect 84 -23791 100 -23757
rect -100 -23899 -84 -23865
rect 84 -23899 100 -23865
rect -146 -23958 -112 -23942
rect -146 -24750 -112 -24734
rect 112 -23958 146 -23942
rect 112 -24750 146 -24734
rect -100 -24827 -84 -24793
rect 84 -24827 100 -24793
rect -100 -24935 -84 -24901
rect 84 -24935 100 -24901
rect -146 -24994 -112 -24978
rect -146 -25786 -112 -25770
rect 112 -24994 146 -24978
rect 112 -25786 146 -25770
rect -100 -25863 -84 -25829
rect 84 -25863 100 -25829
rect -100 -25971 -84 -25937
rect 84 -25971 100 -25937
rect -146 -26030 -112 -26014
rect -146 -26822 -112 -26806
rect 112 -26030 146 -26014
rect 112 -26822 146 -26806
rect -100 -26899 -84 -26865
rect 84 -26899 100 -26865
rect -100 -27007 -84 -26973
rect 84 -27007 100 -26973
rect -146 -27066 -112 -27050
rect -146 -27858 -112 -27842
rect 112 -27066 146 -27050
rect 112 -27858 146 -27842
rect -100 -27935 -84 -27901
rect 84 -27935 100 -27901
rect -100 -28043 -84 -28009
rect 84 -28043 100 -28009
rect -146 -28102 -112 -28086
rect -146 -28894 -112 -28878
rect 112 -28102 146 -28086
rect 112 -28894 146 -28878
rect -100 -28971 -84 -28937
rect 84 -28971 100 -28937
rect -100 -29079 -84 -29045
rect 84 -29079 100 -29045
rect -146 -29138 -112 -29122
rect -146 -29930 -112 -29914
rect 112 -29138 146 -29122
rect 112 -29930 146 -29914
rect -100 -30007 -84 -29973
rect 84 -30007 100 -29973
rect -100 -30115 -84 -30081
rect 84 -30115 100 -30081
rect -146 -30174 -112 -30158
rect -146 -30966 -112 -30950
rect 112 -30174 146 -30158
rect 112 -30966 146 -30950
rect -100 -31043 -84 -31009
rect 84 -31043 100 -31009
rect -100 -31151 -84 -31117
rect 84 -31151 100 -31117
rect -146 -31210 -112 -31194
rect -146 -32002 -112 -31986
rect 112 -31210 146 -31194
rect 112 -32002 146 -31986
rect -100 -32079 -84 -32045
rect 84 -32079 100 -32045
rect -100 -32187 -84 -32153
rect 84 -32187 100 -32153
rect -146 -32246 -112 -32230
rect -146 -33038 -112 -33022
rect 112 -32246 146 -32230
rect 112 -33038 146 -33022
rect -100 -33115 -84 -33081
rect 84 -33115 100 -33081
rect -100 -33223 -84 -33189
rect 84 -33223 100 -33189
rect -146 -33282 -112 -33266
rect -146 -34074 -112 -34058
rect 112 -33282 146 -33266
rect 112 -34074 146 -34058
rect -100 -34151 -84 -34117
rect 84 -34151 100 -34117
rect -100 -34259 -84 -34225
rect 84 -34259 100 -34225
rect -146 -34318 -112 -34302
rect -146 -35110 -112 -35094
rect 112 -34318 146 -34302
rect 112 -35110 146 -35094
rect -100 -35187 -84 -35153
rect 84 -35187 100 -35153
rect -100 -35295 -84 -35261
rect 84 -35295 100 -35261
rect -146 -35354 -112 -35338
rect -146 -36146 -112 -36130
rect 112 -35354 146 -35338
rect 112 -36146 146 -36130
rect -100 -36223 -84 -36189
rect 84 -36223 100 -36189
rect -100 -36331 -84 -36297
rect 84 -36331 100 -36297
rect -146 -36390 -112 -36374
rect -146 -37182 -112 -37166
rect 112 -36390 146 -36374
rect 112 -37182 146 -37166
rect -100 -37259 -84 -37225
rect 84 -37259 100 -37225
rect -100 -37367 -84 -37333
rect 84 -37367 100 -37333
rect -146 -37426 -112 -37410
rect -146 -38218 -112 -38202
rect 112 -37426 146 -37410
rect 112 -38218 146 -38202
rect -100 -38295 -84 -38261
rect 84 -38295 100 -38261
rect -100 -38403 -84 -38369
rect 84 -38403 100 -38369
rect -146 -38462 -112 -38446
rect -146 -39254 -112 -39238
rect 112 -38462 146 -38446
rect 112 -39254 146 -39238
rect -100 -39331 -84 -39297
rect 84 -39331 100 -39297
rect -100 -39439 -84 -39405
rect 84 -39439 100 -39405
rect -146 -39498 -112 -39482
rect -146 -40290 -112 -40274
rect 112 -39498 146 -39482
rect 112 -40290 146 -40274
rect -100 -40367 -84 -40333
rect 84 -40367 100 -40333
rect -100 -40475 -84 -40441
rect 84 -40475 100 -40441
rect -146 -40534 -112 -40518
rect -146 -41326 -112 -41310
rect 112 -40534 146 -40518
rect 112 -41326 146 -41310
rect -100 -41403 -84 -41369
rect 84 -41403 100 -41369
rect -100 -41511 -84 -41477
rect 84 -41511 100 -41477
rect -146 -41570 -112 -41554
rect -146 -42362 -112 -42346
rect 112 -41570 146 -41554
rect 112 -42362 146 -42346
rect -100 -42439 -84 -42405
rect 84 -42439 100 -42405
rect -100 -42547 -84 -42513
rect 84 -42547 100 -42513
rect -146 -42606 -112 -42590
rect -146 -43398 -112 -43382
rect 112 -42606 146 -42590
rect 112 -43398 146 -43382
rect -100 -43475 -84 -43441
rect 84 -43475 100 -43441
rect -100 -43583 -84 -43549
rect 84 -43583 100 -43549
rect -146 -43642 -112 -43626
rect -146 -44434 -112 -44418
rect 112 -43642 146 -43626
rect 112 -44434 146 -44418
rect -100 -44511 -84 -44477
rect 84 -44511 100 -44477
rect -100 -44619 -84 -44585
rect 84 -44619 100 -44585
rect -146 -44678 -112 -44662
rect -146 -45470 -112 -45454
rect 112 -44678 146 -44662
rect 112 -45470 146 -45454
rect -100 -45547 -84 -45513
rect 84 -45547 100 -45513
rect -100 -45655 -84 -45621
rect 84 -45655 100 -45621
rect -146 -45714 -112 -45698
rect -146 -46506 -112 -46490
rect 112 -45714 146 -45698
rect 112 -46506 146 -46490
rect -100 -46583 -84 -46549
rect 84 -46583 100 -46549
rect -100 -46691 -84 -46657
rect 84 -46691 100 -46657
rect -146 -46750 -112 -46734
rect -146 -47542 -112 -47526
rect 112 -46750 146 -46734
rect 112 -47542 146 -47526
rect -100 -47619 -84 -47585
rect 84 -47619 100 -47585
rect -100 -47727 -84 -47693
rect 84 -47727 100 -47693
rect -146 -47786 -112 -47770
rect -146 -48578 -112 -48562
rect 112 -47786 146 -47770
rect 112 -48578 146 -48562
rect -100 -48655 -84 -48621
rect 84 -48655 100 -48621
rect -100 -48763 -84 -48729
rect 84 -48763 100 -48729
rect -146 -48822 -112 -48806
rect -146 -49614 -112 -49598
rect 112 -48822 146 -48806
rect 112 -49614 146 -49598
rect -100 -49691 -84 -49657
rect 84 -49691 100 -49657
rect -100 -49799 -84 -49765
rect 84 -49799 100 -49765
rect -146 -49858 -112 -49842
rect -146 -50650 -112 -50634
rect 112 -49858 146 -49842
rect 112 -50650 146 -50634
rect -100 -50727 -84 -50693
rect 84 -50727 100 -50693
rect -100 -50835 -84 -50801
rect 84 -50835 100 -50801
rect -146 -50894 -112 -50878
rect -146 -51686 -112 -51670
rect 112 -50894 146 -50878
rect 112 -51686 146 -51670
rect -100 -51763 -84 -51729
rect 84 -51763 100 -51729
rect -100 -51871 -84 -51837
rect 84 -51871 100 -51837
rect -146 -51930 -112 -51914
rect -146 -52722 -112 -52706
rect 112 -51930 146 -51914
rect 112 -52722 146 -52706
rect -100 -52799 -84 -52765
rect 84 -52799 100 -52765
rect -100 -52907 -84 -52873
rect 84 -52907 100 -52873
rect -146 -52966 -112 -52950
rect -146 -53758 -112 -53742
rect 112 -52966 146 -52950
rect 112 -53758 146 -53742
rect -100 -53835 -84 -53801
rect 84 -53835 100 -53801
rect -100 -53943 -84 -53909
rect 84 -53943 100 -53909
rect -146 -54002 -112 -53986
rect -146 -54794 -112 -54778
rect 112 -54002 146 -53986
rect 112 -54794 146 -54778
rect -100 -54871 -84 -54837
rect 84 -54871 100 -54837
rect -100 -54979 -84 -54945
rect 84 -54979 100 -54945
rect -146 -55038 -112 -55022
rect -146 -55830 -112 -55814
rect 112 -55038 146 -55022
rect 112 -55830 146 -55814
rect -100 -55907 -84 -55873
rect 84 -55907 100 -55873
rect -100 -56015 -84 -55981
rect 84 -56015 100 -55981
rect -146 -56074 -112 -56058
rect -146 -56866 -112 -56850
rect 112 -56074 146 -56058
rect 112 -56866 146 -56850
rect -100 -56943 -84 -56909
rect 84 -56943 100 -56909
rect -100 -57051 -84 -57017
rect 84 -57051 100 -57017
rect -146 -57110 -112 -57094
rect -146 -57902 -112 -57886
rect 112 -57110 146 -57094
rect 112 -57902 146 -57886
rect -100 -57979 -84 -57945
rect 84 -57979 100 -57945
rect -100 -58087 -84 -58053
rect 84 -58087 100 -58053
rect -146 -58146 -112 -58130
rect -146 -58938 -112 -58922
rect 112 -58146 146 -58130
rect 112 -58938 146 -58922
rect -100 -59015 -84 -58981
rect 84 -59015 100 -58981
rect -100 -59123 -84 -59089
rect 84 -59123 100 -59089
rect -146 -59182 -112 -59166
rect -146 -59974 -112 -59958
rect 112 -59182 146 -59166
rect 112 -59974 146 -59958
rect -100 -60051 -84 -60017
rect 84 -60051 100 -60017
rect -100 -60159 -84 -60125
rect 84 -60159 100 -60125
rect -146 -60218 -112 -60202
rect -146 -61010 -112 -60994
rect 112 -60218 146 -60202
rect 112 -61010 146 -60994
rect -100 -61087 -84 -61053
rect 84 -61087 100 -61053
rect -100 -61195 -84 -61161
rect 84 -61195 100 -61161
rect -146 -61254 -112 -61238
rect -146 -62046 -112 -62030
rect 112 -61254 146 -61238
rect 112 -62046 146 -62030
rect -100 -62123 -84 -62089
rect 84 -62123 100 -62089
rect -100 -62231 -84 -62197
rect 84 -62231 100 -62197
rect -146 -62290 -112 -62274
rect -146 -63082 -112 -63066
rect 112 -62290 146 -62274
rect 112 -63082 146 -63066
rect -100 -63159 -84 -63125
rect 84 -63159 100 -63125
rect -100 -63267 -84 -63233
rect 84 -63267 100 -63233
rect -146 -63326 -112 -63310
rect -146 -64118 -112 -64102
rect 112 -63326 146 -63310
rect 112 -64118 146 -64102
rect -100 -64195 -84 -64161
rect 84 -64195 100 -64161
rect -100 -64303 -84 -64269
rect 84 -64303 100 -64269
rect -146 -64362 -112 -64346
rect -146 -65154 -112 -65138
rect 112 -64362 146 -64346
rect 112 -65154 146 -65138
rect -100 -65231 -84 -65197
rect 84 -65231 100 -65197
rect -100 -65339 -84 -65305
rect 84 -65339 100 -65305
rect -146 -65398 -112 -65382
rect -146 -66190 -112 -66174
rect 112 -65398 146 -65382
rect 112 -66190 146 -66174
rect -100 -66267 -84 -66233
rect 84 -66267 100 -66233
rect -100 -66375 -84 -66341
rect 84 -66375 100 -66341
rect -146 -66434 -112 -66418
rect -146 -67226 -112 -67210
rect 112 -66434 146 -66418
rect 112 -67226 146 -67210
rect -100 -67303 -84 -67269
rect 84 -67303 100 -67269
rect -100 -67411 -84 -67377
rect 84 -67411 100 -67377
rect -146 -67470 -112 -67454
rect -146 -68262 -112 -68246
rect 112 -67470 146 -67454
rect 112 -68262 146 -68246
rect -100 -68339 -84 -68305
rect 84 -68339 100 -68305
rect -100 -68447 -84 -68413
rect 84 -68447 100 -68413
rect -146 -68506 -112 -68490
rect -146 -69298 -112 -69282
rect 112 -68506 146 -68490
rect 112 -69298 146 -69282
rect -100 -69375 -84 -69341
rect 84 -69375 100 -69341
rect -100 -69483 -84 -69449
rect 84 -69483 100 -69449
rect -146 -69542 -112 -69526
rect -146 -70334 -112 -70318
rect 112 -69542 146 -69526
rect 112 -70334 146 -70318
rect -100 -70411 -84 -70377
rect 84 -70411 100 -70377
rect -100 -70519 -84 -70485
rect 84 -70519 100 -70485
rect -146 -70578 -112 -70562
rect -146 -71370 -112 -71354
rect 112 -70578 146 -70562
rect 112 -71370 146 -71354
rect -100 -71447 -84 -71413
rect 84 -71447 100 -71413
rect -100 -71555 -84 -71521
rect 84 -71555 100 -71521
rect -146 -71614 -112 -71598
rect -146 -72406 -112 -72390
rect 112 -71614 146 -71598
rect 112 -72406 146 -72390
rect -100 -72483 -84 -72449
rect 84 -72483 100 -72449
rect -100 -72591 -84 -72557
rect 84 -72591 100 -72557
rect -146 -72650 -112 -72634
rect -146 -73442 -112 -73426
rect 112 -72650 146 -72634
rect 112 -73442 146 -73426
rect -100 -73519 -84 -73485
rect 84 -73519 100 -73485
rect -100 -73627 -84 -73593
rect 84 -73627 100 -73593
rect -146 -73686 -112 -73670
rect -146 -74478 -112 -74462
rect 112 -73686 146 -73670
rect 112 -74478 146 -74462
rect -100 -74555 -84 -74521
rect 84 -74555 100 -74521
rect -100 -74663 -84 -74629
rect 84 -74663 100 -74629
rect -146 -74722 -112 -74706
rect -146 -75514 -112 -75498
rect 112 -74722 146 -74706
rect 112 -75514 146 -75498
rect -100 -75591 -84 -75557
rect 84 -75591 100 -75557
rect -100 -75699 -84 -75665
rect 84 -75699 100 -75665
rect -146 -75758 -112 -75742
rect -146 -76550 -112 -76534
rect 112 -75758 146 -75742
rect 112 -76550 146 -76534
rect -100 -76627 -84 -76593
rect 84 -76627 100 -76593
rect -100 -76735 -84 -76701
rect 84 -76735 100 -76701
rect -146 -76794 -112 -76778
rect -146 -77586 -112 -77570
rect 112 -76794 146 -76778
rect 112 -77586 146 -77570
rect -100 -77663 -84 -77629
rect 84 -77663 100 -77629
rect -100 -77771 -84 -77737
rect 84 -77771 100 -77737
rect -146 -77830 -112 -77814
rect -146 -78622 -112 -78606
rect 112 -77830 146 -77814
rect 112 -78622 146 -78606
rect -100 -78699 -84 -78665
rect 84 -78699 100 -78665
rect -100 -78807 -84 -78773
rect 84 -78807 100 -78773
rect -146 -78866 -112 -78850
rect -146 -79658 -112 -79642
rect 112 -78866 146 -78850
rect 112 -79658 146 -79642
rect -100 -79735 -84 -79701
rect 84 -79735 100 -79701
rect -100 -79843 -84 -79809
rect 84 -79843 100 -79809
rect -146 -79902 -112 -79886
rect -146 -80694 -112 -80678
rect 112 -79902 146 -79886
rect 112 -80694 146 -80678
rect -100 -80771 -84 -80737
rect 84 -80771 100 -80737
rect -100 -80879 -84 -80845
rect 84 -80879 100 -80845
rect -146 -80938 -112 -80922
rect -146 -81730 -112 -81714
rect 112 -80938 146 -80922
rect 112 -81730 146 -81714
rect -100 -81807 -84 -81773
rect 84 -81807 100 -81773
rect -100 -81915 -84 -81881
rect 84 -81915 100 -81881
rect -146 -81974 -112 -81958
rect -146 -82766 -112 -82750
rect 112 -81974 146 -81958
rect 112 -82766 146 -82750
rect -100 -82843 -84 -82809
rect 84 -82843 100 -82809
rect -100 -82951 -84 -82917
rect 84 -82951 100 -82917
rect -146 -83010 -112 -82994
rect -146 -83802 -112 -83786
rect 112 -83010 146 -82994
rect 112 -83802 146 -83786
rect -100 -83879 -84 -83845
rect 84 -83879 100 -83845
rect -100 -83987 -84 -83953
rect 84 -83987 100 -83953
rect -146 -84046 -112 -84030
rect -146 -84838 -112 -84822
rect 112 -84046 146 -84030
rect 112 -84838 146 -84822
rect -100 -84915 -84 -84881
rect 84 -84915 100 -84881
rect -100 -85023 -84 -84989
rect 84 -85023 100 -84989
rect -146 -85082 -112 -85066
rect -146 -85874 -112 -85858
rect 112 -85082 146 -85066
rect 112 -85874 146 -85858
rect -100 -85951 -84 -85917
rect 84 -85951 100 -85917
rect -100 -86059 -84 -86025
rect 84 -86059 100 -86025
rect -146 -86118 -112 -86102
rect -146 -86910 -112 -86894
rect 112 -86118 146 -86102
rect 112 -86910 146 -86894
rect -100 -86987 -84 -86953
rect 84 -86987 100 -86953
rect -100 -87095 -84 -87061
rect 84 -87095 100 -87061
rect -146 -87154 -112 -87138
rect -146 -87946 -112 -87930
rect 112 -87154 146 -87138
rect 112 -87946 146 -87930
rect -100 -88023 -84 -87989
rect 84 -88023 100 -87989
rect -100 -88131 -84 -88097
rect 84 -88131 100 -88097
rect -146 -88190 -112 -88174
rect -146 -88982 -112 -88966
rect 112 -88190 146 -88174
rect 112 -88982 146 -88966
rect -100 -89059 -84 -89025
rect 84 -89059 100 -89025
rect -100 -89167 -84 -89133
rect 84 -89167 100 -89133
rect -146 -89226 -112 -89210
rect -146 -90018 -112 -90002
rect 112 -89226 146 -89210
rect 112 -90018 146 -90002
rect -100 -90095 -84 -90061
rect 84 -90095 100 -90061
rect -100 -90203 -84 -90169
rect 84 -90203 100 -90169
rect -146 -90262 -112 -90246
rect -146 -91054 -112 -91038
rect 112 -90262 146 -90246
rect 112 -91054 146 -91038
rect -100 -91131 -84 -91097
rect 84 -91131 100 -91097
rect -100 -91239 -84 -91205
rect 84 -91239 100 -91205
rect -146 -91298 -112 -91282
rect -146 -92090 -112 -92074
rect 112 -91298 146 -91282
rect 112 -92090 146 -92074
rect -100 -92167 -84 -92133
rect 84 -92167 100 -92133
rect -100 -92275 -84 -92241
rect 84 -92275 100 -92241
rect -146 -92334 -112 -92318
rect -146 -93126 -112 -93110
rect 112 -92334 146 -92318
rect 112 -93126 146 -93110
rect -100 -93203 -84 -93169
rect 84 -93203 100 -93169
rect -100 -93311 -84 -93277
rect 84 -93311 100 -93277
rect -146 -93370 -112 -93354
rect -146 -94162 -112 -94146
rect 112 -93370 146 -93354
rect 112 -94162 146 -94146
rect -100 -94239 -84 -94205
rect 84 -94239 100 -94205
rect -100 -94347 -84 -94313
rect 84 -94347 100 -94313
rect -146 -94406 -112 -94390
rect -146 -95198 -112 -95182
rect 112 -94406 146 -94390
rect 112 -95198 146 -95182
rect -100 -95275 -84 -95241
rect 84 -95275 100 -95241
rect -100 -95383 -84 -95349
rect 84 -95383 100 -95349
rect -146 -95442 -112 -95426
rect -146 -96234 -112 -96218
rect 112 -95442 146 -95426
rect 112 -96234 146 -96218
rect -100 -96311 -84 -96277
rect 84 -96311 100 -96277
rect -100 -96419 -84 -96385
rect 84 -96419 100 -96385
rect -146 -96478 -112 -96462
rect -146 -97270 -112 -97254
rect 112 -96478 146 -96462
rect 112 -97270 146 -97254
rect -100 -97347 -84 -97313
rect 84 -97347 100 -97313
rect -100 -97455 -84 -97421
rect 84 -97455 100 -97421
rect -146 -97514 -112 -97498
rect -146 -98306 -112 -98290
rect 112 -97514 146 -97498
rect 112 -98306 146 -98290
rect -100 -98383 -84 -98349
rect 84 -98383 100 -98349
rect -100 -98491 -84 -98457
rect 84 -98491 100 -98457
rect -146 -98550 -112 -98534
rect -146 -99342 -112 -99326
rect 112 -98550 146 -98534
rect 112 -99342 146 -99326
rect -100 -99419 -84 -99385
rect 84 -99419 100 -99385
rect -100 -99527 -84 -99493
rect 84 -99527 100 -99493
rect -146 -99586 -112 -99570
rect -146 -100378 -112 -100362
rect 112 -99586 146 -99570
rect 112 -100378 146 -100362
rect -100 -100455 -84 -100421
rect 84 -100455 100 -100421
rect -100 -100563 -84 -100529
rect 84 -100563 100 -100529
rect -146 -100622 -112 -100606
rect -146 -101414 -112 -101398
rect 112 -100622 146 -100606
rect 112 -101414 146 -101398
rect -100 -101491 -84 -101457
rect 84 -101491 100 -101457
rect -100 -101599 -84 -101565
rect 84 -101599 100 -101565
rect -146 -101658 -112 -101642
rect -146 -102450 -112 -102434
rect 112 -101658 146 -101642
rect 112 -102450 146 -102434
rect -100 -102527 -84 -102493
rect 84 -102527 100 -102493
rect -100 -102635 -84 -102601
rect 84 -102635 100 -102601
rect -146 -102694 -112 -102678
rect -146 -103486 -112 -103470
rect 112 -102694 146 -102678
rect 112 -103486 146 -103470
rect -100 -103563 -84 -103529
rect 84 -103563 100 -103529
rect -100 -103671 -84 -103637
rect 84 -103671 100 -103637
rect -146 -103730 -112 -103714
rect -146 -104522 -112 -104506
rect 112 -103730 146 -103714
rect 112 -104522 146 -104506
rect -100 -104599 -84 -104565
rect 84 -104599 100 -104565
rect -100 -104707 -84 -104673
rect 84 -104707 100 -104673
rect -146 -104766 -112 -104750
rect -146 -105558 -112 -105542
rect 112 -104766 146 -104750
rect 112 -105558 146 -105542
rect -100 -105635 -84 -105601
rect 84 -105635 100 -105601
rect -100 -105743 -84 -105709
rect 84 -105743 100 -105709
rect -146 -105802 -112 -105786
rect -146 -106594 -112 -106578
rect 112 -105802 146 -105786
rect 112 -106594 146 -106578
rect -100 -106671 -84 -106637
rect 84 -106671 100 -106637
rect -100 -106779 -84 -106745
rect 84 -106779 100 -106745
rect -146 -106838 -112 -106822
rect -146 -107630 -112 -107614
rect 112 -106838 146 -106822
rect 112 -107630 146 -107614
rect -100 -107707 -84 -107673
rect 84 -107707 100 -107673
rect -100 -107815 -84 -107781
rect 84 -107815 100 -107781
rect -146 -107874 -112 -107858
rect -146 -108666 -112 -108650
rect 112 -107874 146 -107858
rect 112 -108666 146 -108650
rect -100 -108743 -84 -108709
rect 84 -108743 100 -108709
rect -100 -108851 -84 -108817
rect 84 -108851 100 -108817
rect -146 -108910 -112 -108894
rect -146 -109702 -112 -109686
rect 112 -108910 146 -108894
rect 112 -109702 146 -109686
rect -100 -109779 -84 -109745
rect 84 -109779 100 -109745
rect -100 -109887 -84 -109853
rect 84 -109887 100 -109853
rect -146 -109946 -112 -109930
rect -146 -110738 -112 -110722
rect 112 -109946 146 -109930
rect 112 -110738 146 -110722
rect -100 -110815 -84 -110781
rect 84 -110815 100 -110781
rect -100 -110923 -84 -110889
rect 84 -110923 100 -110889
rect -146 -110982 -112 -110966
rect -146 -111774 -112 -111758
rect 112 -110982 146 -110966
rect 112 -111774 146 -111758
rect -100 -111851 -84 -111817
rect 84 -111851 100 -111817
rect -100 -111959 -84 -111925
rect 84 -111959 100 -111925
rect -146 -112018 -112 -112002
rect -146 -112810 -112 -112794
rect 112 -112018 146 -112002
rect 112 -112810 146 -112794
rect -100 -112887 -84 -112853
rect 84 -112887 100 -112853
rect -100 -112995 -84 -112961
rect 84 -112995 100 -112961
rect -146 -113054 -112 -113038
rect -146 -113846 -112 -113830
rect 112 -113054 146 -113038
rect 112 -113846 146 -113830
rect -100 -113923 -84 -113889
rect 84 -113923 100 -113889
rect -100 -114031 -84 -113997
rect 84 -114031 100 -113997
rect -146 -114090 -112 -114074
rect -146 -114882 -112 -114866
rect 112 -114090 146 -114074
rect 112 -114882 146 -114866
rect -100 -114959 -84 -114925
rect 84 -114959 100 -114925
rect -100 -115067 -84 -115033
rect 84 -115067 100 -115033
rect -146 -115126 -112 -115110
rect -146 -115918 -112 -115902
rect 112 -115126 146 -115110
rect 112 -115918 146 -115902
rect -100 -115995 -84 -115961
rect 84 -115995 100 -115961
rect -100 -116103 -84 -116069
rect 84 -116103 100 -116069
rect -146 -116162 -112 -116146
rect -146 -116954 -112 -116938
rect 112 -116162 146 -116146
rect 112 -116954 146 -116938
rect -100 -117031 -84 -116997
rect 84 -117031 100 -116997
rect -100 -117139 -84 -117105
rect 84 -117139 100 -117105
rect -146 -117198 -112 -117182
rect -146 -117990 -112 -117974
rect 112 -117198 146 -117182
rect 112 -117990 146 -117974
rect -100 -118067 -84 -118033
rect 84 -118067 100 -118033
rect -100 -118175 -84 -118141
rect 84 -118175 100 -118141
rect -146 -118234 -112 -118218
rect -146 -119026 -112 -119010
rect 112 -118234 146 -118218
rect 112 -119026 146 -119010
rect -100 -119103 -84 -119069
rect 84 -119103 100 -119069
rect -100 -119211 -84 -119177
rect 84 -119211 100 -119177
rect -146 -119270 -112 -119254
rect -146 -120062 -112 -120046
rect 112 -119270 146 -119254
rect 112 -120062 146 -120046
rect -100 -120139 -84 -120105
rect 84 -120139 100 -120105
rect -100 -120247 -84 -120213
rect 84 -120247 100 -120213
rect -146 -120306 -112 -120290
rect -146 -121098 -112 -121082
rect 112 -120306 146 -120290
rect 112 -121098 146 -121082
rect -100 -121175 -84 -121141
rect 84 -121175 100 -121141
rect -100 -121283 -84 -121249
rect 84 -121283 100 -121249
rect -146 -121342 -112 -121326
rect -146 -122134 -112 -122118
rect 112 -121342 146 -121326
rect 112 -122134 146 -122118
rect -100 -122211 -84 -122177
rect 84 -122211 100 -122177
rect -100 -122319 -84 -122285
rect 84 -122319 100 -122285
rect -146 -122378 -112 -122362
rect -146 -123170 -112 -123154
rect 112 -122378 146 -122362
rect 112 -123170 146 -123154
rect -100 -123247 -84 -123213
rect 84 -123247 100 -123213
rect -100 -123355 -84 -123321
rect 84 -123355 100 -123321
rect -146 -123414 -112 -123398
rect -146 -124206 -112 -124190
rect 112 -123414 146 -123398
rect 112 -124206 146 -124190
rect -100 -124283 -84 -124249
rect 84 -124283 100 -124249
rect -100 -124391 -84 -124357
rect 84 -124391 100 -124357
rect -146 -124450 -112 -124434
rect -146 -125242 -112 -125226
rect 112 -124450 146 -124434
rect 112 -125242 146 -125226
rect -100 -125319 -84 -125285
rect 84 -125319 100 -125285
rect -100 -125427 -84 -125393
rect 84 -125427 100 -125393
rect -146 -125486 -112 -125470
rect -146 -126278 -112 -126262
rect 112 -125486 146 -125470
rect 112 -126278 146 -126262
rect -100 -126355 -84 -126321
rect 84 -126355 100 -126321
rect -100 -126463 -84 -126429
rect 84 -126463 100 -126429
rect -146 -126522 -112 -126506
rect -146 -127314 -112 -127298
rect 112 -126522 146 -126506
rect 112 -127314 146 -127298
rect -100 -127391 -84 -127357
rect 84 -127391 100 -127357
rect -100 -127499 -84 -127465
rect 84 -127499 100 -127465
rect -146 -127558 -112 -127542
rect -146 -128350 -112 -128334
rect 112 -127558 146 -127542
rect 112 -128350 146 -128334
rect -100 -128427 -84 -128393
rect 84 -128427 100 -128393
rect -100 -128535 -84 -128501
rect 84 -128535 100 -128501
rect -146 -128594 -112 -128578
rect -146 -129386 -112 -129370
rect 112 -128594 146 -128578
rect 112 -129386 146 -129370
rect -100 -129463 -84 -129429
rect 84 -129463 100 -129429
rect -100 -129571 -84 -129537
rect 84 -129571 100 -129537
rect -146 -129630 -112 -129614
rect -146 -130422 -112 -130406
rect 112 -129630 146 -129614
rect 112 -130422 146 -130406
rect -100 -130499 -84 -130465
rect 84 -130499 100 -130465
rect -100 -130607 -84 -130573
rect 84 -130607 100 -130573
rect -146 -130666 -112 -130650
rect -146 -131458 -112 -131442
rect 112 -130666 146 -130650
rect 112 -131458 146 -131442
rect -100 -131535 -84 -131501
rect 84 -131535 100 -131501
rect -100 -131643 -84 -131609
rect 84 -131643 100 -131609
rect -146 -131702 -112 -131686
rect -146 -132494 -112 -132478
rect 112 -131702 146 -131686
rect 112 -132494 146 -132478
rect -100 -132571 -84 -132537
rect 84 -132571 100 -132537
rect -280 -132675 -246 -132613
rect 246 -132675 280 -132613
rect -280 -132709 -184 -132675
rect 184 -132709 280 -132675
<< viali >>
rect -84 132537 84 132571
rect -146 131702 -112 132478
rect 112 131702 146 132478
rect -84 131609 84 131643
rect -84 131501 84 131535
rect -146 130666 -112 131442
rect 112 130666 146 131442
rect -84 130573 84 130607
rect -84 130465 84 130499
rect -146 129630 -112 130406
rect 112 129630 146 130406
rect -84 129537 84 129571
rect -84 129429 84 129463
rect -146 128594 -112 129370
rect 112 128594 146 129370
rect -84 128501 84 128535
rect -84 128393 84 128427
rect -146 127558 -112 128334
rect 112 127558 146 128334
rect -84 127465 84 127499
rect -84 127357 84 127391
rect -146 126522 -112 127298
rect 112 126522 146 127298
rect -84 126429 84 126463
rect -84 126321 84 126355
rect -146 125486 -112 126262
rect 112 125486 146 126262
rect -84 125393 84 125427
rect -84 125285 84 125319
rect -146 124450 -112 125226
rect 112 124450 146 125226
rect -84 124357 84 124391
rect -84 124249 84 124283
rect -146 123414 -112 124190
rect 112 123414 146 124190
rect -84 123321 84 123355
rect -84 123213 84 123247
rect -146 122378 -112 123154
rect 112 122378 146 123154
rect -84 122285 84 122319
rect -84 122177 84 122211
rect -146 121342 -112 122118
rect 112 121342 146 122118
rect -84 121249 84 121283
rect -84 121141 84 121175
rect -146 120306 -112 121082
rect 112 120306 146 121082
rect -84 120213 84 120247
rect -84 120105 84 120139
rect -146 119270 -112 120046
rect 112 119270 146 120046
rect -84 119177 84 119211
rect -84 119069 84 119103
rect -146 118234 -112 119010
rect 112 118234 146 119010
rect -84 118141 84 118175
rect -84 118033 84 118067
rect -146 117198 -112 117974
rect 112 117198 146 117974
rect -84 117105 84 117139
rect -84 116997 84 117031
rect -146 116162 -112 116938
rect 112 116162 146 116938
rect -84 116069 84 116103
rect -84 115961 84 115995
rect -146 115126 -112 115902
rect 112 115126 146 115902
rect -84 115033 84 115067
rect -84 114925 84 114959
rect -146 114090 -112 114866
rect 112 114090 146 114866
rect -84 113997 84 114031
rect -84 113889 84 113923
rect -146 113054 -112 113830
rect 112 113054 146 113830
rect -84 112961 84 112995
rect -84 112853 84 112887
rect -146 112018 -112 112794
rect 112 112018 146 112794
rect -84 111925 84 111959
rect -84 111817 84 111851
rect -146 110982 -112 111758
rect 112 110982 146 111758
rect -84 110889 84 110923
rect -84 110781 84 110815
rect -146 109946 -112 110722
rect 112 109946 146 110722
rect -84 109853 84 109887
rect -84 109745 84 109779
rect -146 108910 -112 109686
rect 112 108910 146 109686
rect -84 108817 84 108851
rect -84 108709 84 108743
rect -146 107874 -112 108650
rect 112 107874 146 108650
rect -84 107781 84 107815
rect -84 107673 84 107707
rect -146 106838 -112 107614
rect 112 106838 146 107614
rect -84 106745 84 106779
rect -84 106637 84 106671
rect -146 105802 -112 106578
rect 112 105802 146 106578
rect -84 105709 84 105743
rect -84 105601 84 105635
rect -146 104766 -112 105542
rect 112 104766 146 105542
rect -84 104673 84 104707
rect -84 104565 84 104599
rect -146 103730 -112 104506
rect 112 103730 146 104506
rect -84 103637 84 103671
rect -84 103529 84 103563
rect -146 102694 -112 103470
rect 112 102694 146 103470
rect -84 102601 84 102635
rect -84 102493 84 102527
rect -146 101658 -112 102434
rect 112 101658 146 102434
rect -84 101565 84 101599
rect -84 101457 84 101491
rect -146 100622 -112 101398
rect 112 100622 146 101398
rect -84 100529 84 100563
rect -84 100421 84 100455
rect -146 99586 -112 100362
rect 112 99586 146 100362
rect -84 99493 84 99527
rect -84 99385 84 99419
rect -146 98550 -112 99326
rect 112 98550 146 99326
rect -84 98457 84 98491
rect -84 98349 84 98383
rect -146 97514 -112 98290
rect 112 97514 146 98290
rect -84 97421 84 97455
rect -84 97313 84 97347
rect -146 96478 -112 97254
rect 112 96478 146 97254
rect -84 96385 84 96419
rect -84 96277 84 96311
rect -146 95442 -112 96218
rect 112 95442 146 96218
rect -84 95349 84 95383
rect -84 95241 84 95275
rect -146 94406 -112 95182
rect 112 94406 146 95182
rect -84 94313 84 94347
rect -84 94205 84 94239
rect -146 93370 -112 94146
rect 112 93370 146 94146
rect -84 93277 84 93311
rect -84 93169 84 93203
rect -146 92334 -112 93110
rect 112 92334 146 93110
rect -84 92241 84 92275
rect -84 92133 84 92167
rect -146 91298 -112 92074
rect 112 91298 146 92074
rect -84 91205 84 91239
rect -84 91097 84 91131
rect -146 90262 -112 91038
rect 112 90262 146 91038
rect -84 90169 84 90203
rect -84 90061 84 90095
rect -146 89226 -112 90002
rect 112 89226 146 90002
rect -84 89133 84 89167
rect -84 89025 84 89059
rect -146 88190 -112 88966
rect 112 88190 146 88966
rect -84 88097 84 88131
rect -84 87989 84 88023
rect -146 87154 -112 87930
rect 112 87154 146 87930
rect -84 87061 84 87095
rect -84 86953 84 86987
rect -146 86118 -112 86894
rect 112 86118 146 86894
rect -84 86025 84 86059
rect -84 85917 84 85951
rect -146 85082 -112 85858
rect 112 85082 146 85858
rect -84 84989 84 85023
rect -84 84881 84 84915
rect -146 84046 -112 84822
rect 112 84046 146 84822
rect -84 83953 84 83987
rect -84 83845 84 83879
rect -146 83010 -112 83786
rect 112 83010 146 83786
rect -84 82917 84 82951
rect -84 82809 84 82843
rect -146 81974 -112 82750
rect 112 81974 146 82750
rect -84 81881 84 81915
rect -84 81773 84 81807
rect -146 80938 -112 81714
rect 112 80938 146 81714
rect -84 80845 84 80879
rect -84 80737 84 80771
rect -146 79902 -112 80678
rect 112 79902 146 80678
rect -84 79809 84 79843
rect -84 79701 84 79735
rect -146 78866 -112 79642
rect 112 78866 146 79642
rect -84 78773 84 78807
rect -84 78665 84 78699
rect -146 77830 -112 78606
rect 112 77830 146 78606
rect -84 77737 84 77771
rect -84 77629 84 77663
rect -146 76794 -112 77570
rect 112 76794 146 77570
rect -84 76701 84 76735
rect -84 76593 84 76627
rect -146 75758 -112 76534
rect 112 75758 146 76534
rect -84 75665 84 75699
rect -84 75557 84 75591
rect -146 74722 -112 75498
rect 112 74722 146 75498
rect -84 74629 84 74663
rect -84 74521 84 74555
rect -146 73686 -112 74462
rect 112 73686 146 74462
rect -84 73593 84 73627
rect -84 73485 84 73519
rect -146 72650 -112 73426
rect 112 72650 146 73426
rect -84 72557 84 72591
rect -84 72449 84 72483
rect -146 71614 -112 72390
rect 112 71614 146 72390
rect -84 71521 84 71555
rect -84 71413 84 71447
rect -146 70578 -112 71354
rect 112 70578 146 71354
rect -84 70485 84 70519
rect -84 70377 84 70411
rect -146 69542 -112 70318
rect 112 69542 146 70318
rect -84 69449 84 69483
rect -84 69341 84 69375
rect -146 68506 -112 69282
rect 112 68506 146 69282
rect -84 68413 84 68447
rect -84 68305 84 68339
rect -146 67470 -112 68246
rect 112 67470 146 68246
rect -84 67377 84 67411
rect -84 67269 84 67303
rect -146 66434 -112 67210
rect 112 66434 146 67210
rect -84 66341 84 66375
rect -84 66233 84 66267
rect -146 65398 -112 66174
rect 112 65398 146 66174
rect -84 65305 84 65339
rect -84 65197 84 65231
rect -146 64362 -112 65138
rect 112 64362 146 65138
rect -84 64269 84 64303
rect -84 64161 84 64195
rect -146 63326 -112 64102
rect 112 63326 146 64102
rect -84 63233 84 63267
rect -84 63125 84 63159
rect -146 62290 -112 63066
rect 112 62290 146 63066
rect -84 62197 84 62231
rect -84 62089 84 62123
rect -146 61254 -112 62030
rect 112 61254 146 62030
rect -84 61161 84 61195
rect -84 61053 84 61087
rect -146 60218 -112 60994
rect 112 60218 146 60994
rect -84 60125 84 60159
rect -84 60017 84 60051
rect -146 59182 -112 59958
rect 112 59182 146 59958
rect -84 59089 84 59123
rect -84 58981 84 59015
rect -146 58146 -112 58922
rect 112 58146 146 58922
rect -84 58053 84 58087
rect -84 57945 84 57979
rect -146 57110 -112 57886
rect 112 57110 146 57886
rect -84 57017 84 57051
rect -84 56909 84 56943
rect -146 56074 -112 56850
rect 112 56074 146 56850
rect -84 55981 84 56015
rect -84 55873 84 55907
rect -146 55038 -112 55814
rect 112 55038 146 55814
rect -84 54945 84 54979
rect -84 54837 84 54871
rect -146 54002 -112 54778
rect 112 54002 146 54778
rect -84 53909 84 53943
rect -84 53801 84 53835
rect -146 52966 -112 53742
rect 112 52966 146 53742
rect -84 52873 84 52907
rect -84 52765 84 52799
rect -146 51930 -112 52706
rect 112 51930 146 52706
rect -84 51837 84 51871
rect -84 51729 84 51763
rect -146 50894 -112 51670
rect 112 50894 146 51670
rect -84 50801 84 50835
rect -84 50693 84 50727
rect -146 49858 -112 50634
rect 112 49858 146 50634
rect -84 49765 84 49799
rect -84 49657 84 49691
rect -146 48822 -112 49598
rect 112 48822 146 49598
rect -84 48729 84 48763
rect -84 48621 84 48655
rect -146 47786 -112 48562
rect 112 47786 146 48562
rect -84 47693 84 47727
rect -84 47585 84 47619
rect -146 46750 -112 47526
rect 112 46750 146 47526
rect -84 46657 84 46691
rect -84 46549 84 46583
rect -146 45714 -112 46490
rect 112 45714 146 46490
rect -84 45621 84 45655
rect -84 45513 84 45547
rect -146 44678 -112 45454
rect 112 44678 146 45454
rect -84 44585 84 44619
rect -84 44477 84 44511
rect -146 43642 -112 44418
rect 112 43642 146 44418
rect -84 43549 84 43583
rect -84 43441 84 43475
rect -146 42606 -112 43382
rect 112 42606 146 43382
rect -84 42513 84 42547
rect -84 42405 84 42439
rect -146 41570 -112 42346
rect 112 41570 146 42346
rect -84 41477 84 41511
rect -84 41369 84 41403
rect -146 40534 -112 41310
rect 112 40534 146 41310
rect -84 40441 84 40475
rect -84 40333 84 40367
rect -146 39498 -112 40274
rect 112 39498 146 40274
rect -84 39405 84 39439
rect -84 39297 84 39331
rect -146 38462 -112 39238
rect 112 38462 146 39238
rect -84 38369 84 38403
rect -84 38261 84 38295
rect -146 37426 -112 38202
rect 112 37426 146 38202
rect -84 37333 84 37367
rect -84 37225 84 37259
rect -146 36390 -112 37166
rect 112 36390 146 37166
rect -84 36297 84 36331
rect -84 36189 84 36223
rect -146 35354 -112 36130
rect 112 35354 146 36130
rect -84 35261 84 35295
rect -84 35153 84 35187
rect -146 34318 -112 35094
rect 112 34318 146 35094
rect -84 34225 84 34259
rect -84 34117 84 34151
rect -146 33282 -112 34058
rect 112 33282 146 34058
rect -84 33189 84 33223
rect -84 33081 84 33115
rect -146 32246 -112 33022
rect 112 32246 146 33022
rect -84 32153 84 32187
rect -84 32045 84 32079
rect -146 31210 -112 31986
rect 112 31210 146 31986
rect -84 31117 84 31151
rect -84 31009 84 31043
rect -146 30174 -112 30950
rect 112 30174 146 30950
rect -84 30081 84 30115
rect -84 29973 84 30007
rect -146 29138 -112 29914
rect 112 29138 146 29914
rect -84 29045 84 29079
rect -84 28937 84 28971
rect -146 28102 -112 28878
rect 112 28102 146 28878
rect -84 28009 84 28043
rect -84 27901 84 27935
rect -146 27066 -112 27842
rect 112 27066 146 27842
rect -84 26973 84 27007
rect -84 26865 84 26899
rect -146 26030 -112 26806
rect 112 26030 146 26806
rect -84 25937 84 25971
rect -84 25829 84 25863
rect -146 24994 -112 25770
rect 112 24994 146 25770
rect -84 24901 84 24935
rect -84 24793 84 24827
rect -146 23958 -112 24734
rect 112 23958 146 24734
rect -84 23865 84 23899
rect -84 23757 84 23791
rect -146 22922 -112 23698
rect 112 22922 146 23698
rect -84 22829 84 22863
rect -84 22721 84 22755
rect -146 21886 -112 22662
rect 112 21886 146 22662
rect -84 21793 84 21827
rect -84 21685 84 21719
rect -146 20850 -112 21626
rect 112 20850 146 21626
rect -84 20757 84 20791
rect -84 20649 84 20683
rect -146 19814 -112 20590
rect 112 19814 146 20590
rect -84 19721 84 19755
rect -84 19613 84 19647
rect -146 18778 -112 19554
rect 112 18778 146 19554
rect -84 18685 84 18719
rect -84 18577 84 18611
rect -146 17742 -112 18518
rect 112 17742 146 18518
rect -84 17649 84 17683
rect -84 17541 84 17575
rect -146 16706 -112 17482
rect 112 16706 146 17482
rect -84 16613 84 16647
rect -84 16505 84 16539
rect -146 15670 -112 16446
rect 112 15670 146 16446
rect -84 15577 84 15611
rect -84 15469 84 15503
rect -146 14634 -112 15410
rect 112 14634 146 15410
rect -84 14541 84 14575
rect -84 14433 84 14467
rect -146 13598 -112 14374
rect 112 13598 146 14374
rect -84 13505 84 13539
rect -84 13397 84 13431
rect -146 12562 -112 13338
rect 112 12562 146 13338
rect -84 12469 84 12503
rect -84 12361 84 12395
rect -146 11526 -112 12302
rect 112 11526 146 12302
rect -84 11433 84 11467
rect -84 11325 84 11359
rect -146 10490 -112 11266
rect 112 10490 146 11266
rect -84 10397 84 10431
rect -84 10289 84 10323
rect -146 9454 -112 10230
rect 112 9454 146 10230
rect -84 9361 84 9395
rect -84 9253 84 9287
rect -146 8418 -112 9194
rect 112 8418 146 9194
rect -84 8325 84 8359
rect -84 8217 84 8251
rect -146 7382 -112 8158
rect 112 7382 146 8158
rect -84 7289 84 7323
rect -84 7181 84 7215
rect -146 6346 -112 7122
rect 112 6346 146 7122
rect -84 6253 84 6287
rect -84 6145 84 6179
rect -146 5310 -112 6086
rect 112 5310 146 6086
rect -84 5217 84 5251
rect -84 5109 84 5143
rect -146 4274 -112 5050
rect 112 4274 146 5050
rect -84 4181 84 4215
rect -84 4073 84 4107
rect -146 3238 -112 4014
rect 112 3238 146 4014
rect -84 3145 84 3179
rect -84 3037 84 3071
rect -146 2202 -112 2978
rect 112 2202 146 2978
rect -84 2109 84 2143
rect -84 2001 84 2035
rect -146 1166 -112 1942
rect 112 1166 146 1942
rect -84 1073 84 1107
rect -84 965 84 999
rect -146 130 -112 906
rect 112 130 146 906
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -906 -112 -130
rect 112 -906 146 -130
rect -84 -999 84 -965
rect -84 -1107 84 -1073
rect -146 -1942 -112 -1166
rect 112 -1942 146 -1166
rect -84 -2035 84 -2001
rect -84 -2143 84 -2109
rect -146 -2978 -112 -2202
rect 112 -2978 146 -2202
rect -84 -3071 84 -3037
rect -84 -3179 84 -3145
rect -146 -4014 -112 -3238
rect 112 -4014 146 -3238
rect -84 -4107 84 -4073
rect -84 -4215 84 -4181
rect -146 -5050 -112 -4274
rect 112 -5050 146 -4274
rect -84 -5143 84 -5109
rect -84 -5251 84 -5217
rect -146 -6086 -112 -5310
rect 112 -6086 146 -5310
rect -84 -6179 84 -6145
rect -84 -6287 84 -6253
rect -146 -7122 -112 -6346
rect 112 -7122 146 -6346
rect -84 -7215 84 -7181
rect -84 -7323 84 -7289
rect -146 -8158 -112 -7382
rect 112 -8158 146 -7382
rect -84 -8251 84 -8217
rect -84 -8359 84 -8325
rect -146 -9194 -112 -8418
rect 112 -9194 146 -8418
rect -84 -9287 84 -9253
rect -84 -9395 84 -9361
rect -146 -10230 -112 -9454
rect 112 -10230 146 -9454
rect -84 -10323 84 -10289
rect -84 -10431 84 -10397
rect -146 -11266 -112 -10490
rect 112 -11266 146 -10490
rect -84 -11359 84 -11325
rect -84 -11467 84 -11433
rect -146 -12302 -112 -11526
rect 112 -12302 146 -11526
rect -84 -12395 84 -12361
rect -84 -12503 84 -12469
rect -146 -13338 -112 -12562
rect 112 -13338 146 -12562
rect -84 -13431 84 -13397
rect -84 -13539 84 -13505
rect -146 -14374 -112 -13598
rect 112 -14374 146 -13598
rect -84 -14467 84 -14433
rect -84 -14575 84 -14541
rect -146 -15410 -112 -14634
rect 112 -15410 146 -14634
rect -84 -15503 84 -15469
rect -84 -15611 84 -15577
rect -146 -16446 -112 -15670
rect 112 -16446 146 -15670
rect -84 -16539 84 -16505
rect -84 -16647 84 -16613
rect -146 -17482 -112 -16706
rect 112 -17482 146 -16706
rect -84 -17575 84 -17541
rect -84 -17683 84 -17649
rect -146 -18518 -112 -17742
rect 112 -18518 146 -17742
rect -84 -18611 84 -18577
rect -84 -18719 84 -18685
rect -146 -19554 -112 -18778
rect 112 -19554 146 -18778
rect -84 -19647 84 -19613
rect -84 -19755 84 -19721
rect -146 -20590 -112 -19814
rect 112 -20590 146 -19814
rect -84 -20683 84 -20649
rect -84 -20791 84 -20757
rect -146 -21626 -112 -20850
rect 112 -21626 146 -20850
rect -84 -21719 84 -21685
rect -84 -21827 84 -21793
rect -146 -22662 -112 -21886
rect 112 -22662 146 -21886
rect -84 -22755 84 -22721
rect -84 -22863 84 -22829
rect -146 -23698 -112 -22922
rect 112 -23698 146 -22922
rect -84 -23791 84 -23757
rect -84 -23899 84 -23865
rect -146 -24734 -112 -23958
rect 112 -24734 146 -23958
rect -84 -24827 84 -24793
rect -84 -24935 84 -24901
rect -146 -25770 -112 -24994
rect 112 -25770 146 -24994
rect -84 -25863 84 -25829
rect -84 -25971 84 -25937
rect -146 -26806 -112 -26030
rect 112 -26806 146 -26030
rect -84 -26899 84 -26865
rect -84 -27007 84 -26973
rect -146 -27842 -112 -27066
rect 112 -27842 146 -27066
rect -84 -27935 84 -27901
rect -84 -28043 84 -28009
rect -146 -28878 -112 -28102
rect 112 -28878 146 -28102
rect -84 -28971 84 -28937
rect -84 -29079 84 -29045
rect -146 -29914 -112 -29138
rect 112 -29914 146 -29138
rect -84 -30007 84 -29973
rect -84 -30115 84 -30081
rect -146 -30950 -112 -30174
rect 112 -30950 146 -30174
rect -84 -31043 84 -31009
rect -84 -31151 84 -31117
rect -146 -31986 -112 -31210
rect 112 -31986 146 -31210
rect -84 -32079 84 -32045
rect -84 -32187 84 -32153
rect -146 -33022 -112 -32246
rect 112 -33022 146 -32246
rect -84 -33115 84 -33081
rect -84 -33223 84 -33189
rect -146 -34058 -112 -33282
rect 112 -34058 146 -33282
rect -84 -34151 84 -34117
rect -84 -34259 84 -34225
rect -146 -35094 -112 -34318
rect 112 -35094 146 -34318
rect -84 -35187 84 -35153
rect -84 -35295 84 -35261
rect -146 -36130 -112 -35354
rect 112 -36130 146 -35354
rect -84 -36223 84 -36189
rect -84 -36331 84 -36297
rect -146 -37166 -112 -36390
rect 112 -37166 146 -36390
rect -84 -37259 84 -37225
rect -84 -37367 84 -37333
rect -146 -38202 -112 -37426
rect 112 -38202 146 -37426
rect -84 -38295 84 -38261
rect -84 -38403 84 -38369
rect -146 -39238 -112 -38462
rect 112 -39238 146 -38462
rect -84 -39331 84 -39297
rect -84 -39439 84 -39405
rect -146 -40274 -112 -39498
rect 112 -40274 146 -39498
rect -84 -40367 84 -40333
rect -84 -40475 84 -40441
rect -146 -41310 -112 -40534
rect 112 -41310 146 -40534
rect -84 -41403 84 -41369
rect -84 -41511 84 -41477
rect -146 -42346 -112 -41570
rect 112 -42346 146 -41570
rect -84 -42439 84 -42405
rect -84 -42547 84 -42513
rect -146 -43382 -112 -42606
rect 112 -43382 146 -42606
rect -84 -43475 84 -43441
rect -84 -43583 84 -43549
rect -146 -44418 -112 -43642
rect 112 -44418 146 -43642
rect -84 -44511 84 -44477
rect -84 -44619 84 -44585
rect -146 -45454 -112 -44678
rect 112 -45454 146 -44678
rect -84 -45547 84 -45513
rect -84 -45655 84 -45621
rect -146 -46490 -112 -45714
rect 112 -46490 146 -45714
rect -84 -46583 84 -46549
rect -84 -46691 84 -46657
rect -146 -47526 -112 -46750
rect 112 -47526 146 -46750
rect -84 -47619 84 -47585
rect -84 -47727 84 -47693
rect -146 -48562 -112 -47786
rect 112 -48562 146 -47786
rect -84 -48655 84 -48621
rect -84 -48763 84 -48729
rect -146 -49598 -112 -48822
rect 112 -49598 146 -48822
rect -84 -49691 84 -49657
rect -84 -49799 84 -49765
rect -146 -50634 -112 -49858
rect 112 -50634 146 -49858
rect -84 -50727 84 -50693
rect -84 -50835 84 -50801
rect -146 -51670 -112 -50894
rect 112 -51670 146 -50894
rect -84 -51763 84 -51729
rect -84 -51871 84 -51837
rect -146 -52706 -112 -51930
rect 112 -52706 146 -51930
rect -84 -52799 84 -52765
rect -84 -52907 84 -52873
rect -146 -53742 -112 -52966
rect 112 -53742 146 -52966
rect -84 -53835 84 -53801
rect -84 -53943 84 -53909
rect -146 -54778 -112 -54002
rect 112 -54778 146 -54002
rect -84 -54871 84 -54837
rect -84 -54979 84 -54945
rect -146 -55814 -112 -55038
rect 112 -55814 146 -55038
rect -84 -55907 84 -55873
rect -84 -56015 84 -55981
rect -146 -56850 -112 -56074
rect 112 -56850 146 -56074
rect -84 -56943 84 -56909
rect -84 -57051 84 -57017
rect -146 -57886 -112 -57110
rect 112 -57886 146 -57110
rect -84 -57979 84 -57945
rect -84 -58087 84 -58053
rect -146 -58922 -112 -58146
rect 112 -58922 146 -58146
rect -84 -59015 84 -58981
rect -84 -59123 84 -59089
rect -146 -59958 -112 -59182
rect 112 -59958 146 -59182
rect -84 -60051 84 -60017
rect -84 -60159 84 -60125
rect -146 -60994 -112 -60218
rect 112 -60994 146 -60218
rect -84 -61087 84 -61053
rect -84 -61195 84 -61161
rect -146 -62030 -112 -61254
rect 112 -62030 146 -61254
rect -84 -62123 84 -62089
rect -84 -62231 84 -62197
rect -146 -63066 -112 -62290
rect 112 -63066 146 -62290
rect -84 -63159 84 -63125
rect -84 -63267 84 -63233
rect -146 -64102 -112 -63326
rect 112 -64102 146 -63326
rect -84 -64195 84 -64161
rect -84 -64303 84 -64269
rect -146 -65138 -112 -64362
rect 112 -65138 146 -64362
rect -84 -65231 84 -65197
rect -84 -65339 84 -65305
rect -146 -66174 -112 -65398
rect 112 -66174 146 -65398
rect -84 -66267 84 -66233
rect -84 -66375 84 -66341
rect -146 -67210 -112 -66434
rect 112 -67210 146 -66434
rect -84 -67303 84 -67269
rect -84 -67411 84 -67377
rect -146 -68246 -112 -67470
rect 112 -68246 146 -67470
rect -84 -68339 84 -68305
rect -84 -68447 84 -68413
rect -146 -69282 -112 -68506
rect 112 -69282 146 -68506
rect -84 -69375 84 -69341
rect -84 -69483 84 -69449
rect -146 -70318 -112 -69542
rect 112 -70318 146 -69542
rect -84 -70411 84 -70377
rect -84 -70519 84 -70485
rect -146 -71354 -112 -70578
rect 112 -71354 146 -70578
rect -84 -71447 84 -71413
rect -84 -71555 84 -71521
rect -146 -72390 -112 -71614
rect 112 -72390 146 -71614
rect -84 -72483 84 -72449
rect -84 -72591 84 -72557
rect -146 -73426 -112 -72650
rect 112 -73426 146 -72650
rect -84 -73519 84 -73485
rect -84 -73627 84 -73593
rect -146 -74462 -112 -73686
rect 112 -74462 146 -73686
rect -84 -74555 84 -74521
rect -84 -74663 84 -74629
rect -146 -75498 -112 -74722
rect 112 -75498 146 -74722
rect -84 -75591 84 -75557
rect -84 -75699 84 -75665
rect -146 -76534 -112 -75758
rect 112 -76534 146 -75758
rect -84 -76627 84 -76593
rect -84 -76735 84 -76701
rect -146 -77570 -112 -76794
rect 112 -77570 146 -76794
rect -84 -77663 84 -77629
rect -84 -77771 84 -77737
rect -146 -78606 -112 -77830
rect 112 -78606 146 -77830
rect -84 -78699 84 -78665
rect -84 -78807 84 -78773
rect -146 -79642 -112 -78866
rect 112 -79642 146 -78866
rect -84 -79735 84 -79701
rect -84 -79843 84 -79809
rect -146 -80678 -112 -79902
rect 112 -80678 146 -79902
rect -84 -80771 84 -80737
rect -84 -80879 84 -80845
rect -146 -81714 -112 -80938
rect 112 -81714 146 -80938
rect -84 -81807 84 -81773
rect -84 -81915 84 -81881
rect -146 -82750 -112 -81974
rect 112 -82750 146 -81974
rect -84 -82843 84 -82809
rect -84 -82951 84 -82917
rect -146 -83786 -112 -83010
rect 112 -83786 146 -83010
rect -84 -83879 84 -83845
rect -84 -83987 84 -83953
rect -146 -84822 -112 -84046
rect 112 -84822 146 -84046
rect -84 -84915 84 -84881
rect -84 -85023 84 -84989
rect -146 -85858 -112 -85082
rect 112 -85858 146 -85082
rect -84 -85951 84 -85917
rect -84 -86059 84 -86025
rect -146 -86894 -112 -86118
rect 112 -86894 146 -86118
rect -84 -86987 84 -86953
rect -84 -87095 84 -87061
rect -146 -87930 -112 -87154
rect 112 -87930 146 -87154
rect -84 -88023 84 -87989
rect -84 -88131 84 -88097
rect -146 -88966 -112 -88190
rect 112 -88966 146 -88190
rect -84 -89059 84 -89025
rect -84 -89167 84 -89133
rect -146 -90002 -112 -89226
rect 112 -90002 146 -89226
rect -84 -90095 84 -90061
rect -84 -90203 84 -90169
rect -146 -91038 -112 -90262
rect 112 -91038 146 -90262
rect -84 -91131 84 -91097
rect -84 -91239 84 -91205
rect -146 -92074 -112 -91298
rect 112 -92074 146 -91298
rect -84 -92167 84 -92133
rect -84 -92275 84 -92241
rect -146 -93110 -112 -92334
rect 112 -93110 146 -92334
rect -84 -93203 84 -93169
rect -84 -93311 84 -93277
rect -146 -94146 -112 -93370
rect 112 -94146 146 -93370
rect -84 -94239 84 -94205
rect -84 -94347 84 -94313
rect -146 -95182 -112 -94406
rect 112 -95182 146 -94406
rect -84 -95275 84 -95241
rect -84 -95383 84 -95349
rect -146 -96218 -112 -95442
rect 112 -96218 146 -95442
rect -84 -96311 84 -96277
rect -84 -96419 84 -96385
rect -146 -97254 -112 -96478
rect 112 -97254 146 -96478
rect -84 -97347 84 -97313
rect -84 -97455 84 -97421
rect -146 -98290 -112 -97514
rect 112 -98290 146 -97514
rect -84 -98383 84 -98349
rect -84 -98491 84 -98457
rect -146 -99326 -112 -98550
rect 112 -99326 146 -98550
rect -84 -99419 84 -99385
rect -84 -99527 84 -99493
rect -146 -100362 -112 -99586
rect 112 -100362 146 -99586
rect -84 -100455 84 -100421
rect -84 -100563 84 -100529
rect -146 -101398 -112 -100622
rect 112 -101398 146 -100622
rect -84 -101491 84 -101457
rect -84 -101599 84 -101565
rect -146 -102434 -112 -101658
rect 112 -102434 146 -101658
rect -84 -102527 84 -102493
rect -84 -102635 84 -102601
rect -146 -103470 -112 -102694
rect 112 -103470 146 -102694
rect -84 -103563 84 -103529
rect -84 -103671 84 -103637
rect -146 -104506 -112 -103730
rect 112 -104506 146 -103730
rect -84 -104599 84 -104565
rect -84 -104707 84 -104673
rect -146 -105542 -112 -104766
rect 112 -105542 146 -104766
rect -84 -105635 84 -105601
rect -84 -105743 84 -105709
rect -146 -106578 -112 -105802
rect 112 -106578 146 -105802
rect -84 -106671 84 -106637
rect -84 -106779 84 -106745
rect -146 -107614 -112 -106838
rect 112 -107614 146 -106838
rect -84 -107707 84 -107673
rect -84 -107815 84 -107781
rect -146 -108650 -112 -107874
rect 112 -108650 146 -107874
rect -84 -108743 84 -108709
rect -84 -108851 84 -108817
rect -146 -109686 -112 -108910
rect 112 -109686 146 -108910
rect -84 -109779 84 -109745
rect -84 -109887 84 -109853
rect -146 -110722 -112 -109946
rect 112 -110722 146 -109946
rect -84 -110815 84 -110781
rect -84 -110923 84 -110889
rect -146 -111758 -112 -110982
rect 112 -111758 146 -110982
rect -84 -111851 84 -111817
rect -84 -111959 84 -111925
rect -146 -112794 -112 -112018
rect 112 -112794 146 -112018
rect -84 -112887 84 -112853
rect -84 -112995 84 -112961
rect -146 -113830 -112 -113054
rect 112 -113830 146 -113054
rect -84 -113923 84 -113889
rect -84 -114031 84 -113997
rect -146 -114866 -112 -114090
rect 112 -114866 146 -114090
rect -84 -114959 84 -114925
rect -84 -115067 84 -115033
rect -146 -115902 -112 -115126
rect 112 -115902 146 -115126
rect -84 -115995 84 -115961
rect -84 -116103 84 -116069
rect -146 -116938 -112 -116162
rect 112 -116938 146 -116162
rect -84 -117031 84 -116997
rect -84 -117139 84 -117105
rect -146 -117974 -112 -117198
rect 112 -117974 146 -117198
rect -84 -118067 84 -118033
rect -84 -118175 84 -118141
rect -146 -119010 -112 -118234
rect 112 -119010 146 -118234
rect -84 -119103 84 -119069
rect -84 -119211 84 -119177
rect -146 -120046 -112 -119270
rect 112 -120046 146 -119270
rect -84 -120139 84 -120105
rect -84 -120247 84 -120213
rect -146 -121082 -112 -120306
rect 112 -121082 146 -120306
rect -84 -121175 84 -121141
rect -84 -121283 84 -121249
rect -146 -122118 -112 -121342
rect 112 -122118 146 -121342
rect -84 -122211 84 -122177
rect -84 -122319 84 -122285
rect -146 -123154 -112 -122378
rect 112 -123154 146 -122378
rect -84 -123247 84 -123213
rect -84 -123355 84 -123321
rect -146 -124190 -112 -123414
rect 112 -124190 146 -123414
rect -84 -124283 84 -124249
rect -84 -124391 84 -124357
rect -146 -125226 -112 -124450
rect 112 -125226 146 -124450
rect -84 -125319 84 -125285
rect -84 -125427 84 -125393
rect -146 -126262 -112 -125486
rect 112 -126262 146 -125486
rect -84 -126355 84 -126321
rect -84 -126463 84 -126429
rect -146 -127298 -112 -126522
rect 112 -127298 146 -126522
rect -84 -127391 84 -127357
rect -84 -127499 84 -127465
rect -146 -128334 -112 -127558
rect 112 -128334 146 -127558
rect -84 -128427 84 -128393
rect -84 -128535 84 -128501
rect -146 -129370 -112 -128594
rect 112 -129370 146 -128594
rect -84 -129463 84 -129429
rect -84 -129571 84 -129537
rect -146 -130406 -112 -129630
rect 112 -130406 146 -129630
rect -84 -130499 84 -130465
rect -84 -130607 84 -130573
rect -146 -131442 -112 -130666
rect 112 -131442 146 -130666
rect -84 -131535 84 -131501
rect -84 -131643 84 -131609
rect -146 -132478 -112 -131702
rect 112 -132478 146 -131702
rect -84 -132571 84 -132537
<< metal1 >>
rect -96 132571 96 132577
rect -96 132537 -84 132571
rect 84 132537 96 132571
rect -96 132531 96 132537
rect -152 132478 -106 132490
rect -152 131702 -146 132478
rect -112 131702 -106 132478
rect -152 131690 -106 131702
rect 106 132478 152 132490
rect 106 131702 112 132478
rect 146 131702 152 132478
rect 106 131690 152 131702
rect -96 131643 96 131649
rect -96 131609 -84 131643
rect 84 131609 96 131643
rect -96 131603 96 131609
rect -96 131535 96 131541
rect -96 131501 -84 131535
rect 84 131501 96 131535
rect -96 131495 96 131501
rect -152 131442 -106 131454
rect -152 130666 -146 131442
rect -112 130666 -106 131442
rect -152 130654 -106 130666
rect 106 131442 152 131454
rect 106 130666 112 131442
rect 146 130666 152 131442
rect 106 130654 152 130666
rect -96 130607 96 130613
rect -96 130573 -84 130607
rect 84 130573 96 130607
rect -96 130567 96 130573
rect -96 130499 96 130505
rect -96 130465 -84 130499
rect 84 130465 96 130499
rect -96 130459 96 130465
rect -152 130406 -106 130418
rect -152 129630 -146 130406
rect -112 129630 -106 130406
rect -152 129618 -106 129630
rect 106 130406 152 130418
rect 106 129630 112 130406
rect 146 129630 152 130406
rect 106 129618 152 129630
rect -96 129571 96 129577
rect -96 129537 -84 129571
rect 84 129537 96 129571
rect -96 129531 96 129537
rect -96 129463 96 129469
rect -96 129429 -84 129463
rect 84 129429 96 129463
rect -96 129423 96 129429
rect -152 129370 -106 129382
rect -152 128594 -146 129370
rect -112 128594 -106 129370
rect -152 128582 -106 128594
rect 106 129370 152 129382
rect 106 128594 112 129370
rect 146 128594 152 129370
rect 106 128582 152 128594
rect -96 128535 96 128541
rect -96 128501 -84 128535
rect 84 128501 96 128535
rect -96 128495 96 128501
rect -96 128427 96 128433
rect -96 128393 -84 128427
rect 84 128393 96 128427
rect -96 128387 96 128393
rect -152 128334 -106 128346
rect -152 127558 -146 128334
rect -112 127558 -106 128334
rect -152 127546 -106 127558
rect 106 128334 152 128346
rect 106 127558 112 128334
rect 146 127558 152 128334
rect 106 127546 152 127558
rect -96 127499 96 127505
rect -96 127465 -84 127499
rect 84 127465 96 127499
rect -96 127459 96 127465
rect -96 127391 96 127397
rect -96 127357 -84 127391
rect 84 127357 96 127391
rect -96 127351 96 127357
rect -152 127298 -106 127310
rect -152 126522 -146 127298
rect -112 126522 -106 127298
rect -152 126510 -106 126522
rect 106 127298 152 127310
rect 106 126522 112 127298
rect 146 126522 152 127298
rect 106 126510 152 126522
rect -96 126463 96 126469
rect -96 126429 -84 126463
rect 84 126429 96 126463
rect -96 126423 96 126429
rect -96 126355 96 126361
rect -96 126321 -84 126355
rect 84 126321 96 126355
rect -96 126315 96 126321
rect -152 126262 -106 126274
rect -152 125486 -146 126262
rect -112 125486 -106 126262
rect -152 125474 -106 125486
rect 106 126262 152 126274
rect 106 125486 112 126262
rect 146 125486 152 126262
rect 106 125474 152 125486
rect -96 125427 96 125433
rect -96 125393 -84 125427
rect 84 125393 96 125427
rect -96 125387 96 125393
rect -96 125319 96 125325
rect -96 125285 -84 125319
rect 84 125285 96 125319
rect -96 125279 96 125285
rect -152 125226 -106 125238
rect -152 124450 -146 125226
rect -112 124450 -106 125226
rect -152 124438 -106 124450
rect 106 125226 152 125238
rect 106 124450 112 125226
rect 146 124450 152 125226
rect 106 124438 152 124450
rect -96 124391 96 124397
rect -96 124357 -84 124391
rect 84 124357 96 124391
rect -96 124351 96 124357
rect -96 124283 96 124289
rect -96 124249 -84 124283
rect 84 124249 96 124283
rect -96 124243 96 124249
rect -152 124190 -106 124202
rect -152 123414 -146 124190
rect -112 123414 -106 124190
rect -152 123402 -106 123414
rect 106 124190 152 124202
rect 106 123414 112 124190
rect 146 123414 152 124190
rect 106 123402 152 123414
rect -96 123355 96 123361
rect -96 123321 -84 123355
rect 84 123321 96 123355
rect -96 123315 96 123321
rect -96 123247 96 123253
rect -96 123213 -84 123247
rect 84 123213 96 123247
rect -96 123207 96 123213
rect -152 123154 -106 123166
rect -152 122378 -146 123154
rect -112 122378 -106 123154
rect -152 122366 -106 122378
rect 106 123154 152 123166
rect 106 122378 112 123154
rect 146 122378 152 123154
rect 106 122366 152 122378
rect -96 122319 96 122325
rect -96 122285 -84 122319
rect 84 122285 96 122319
rect -96 122279 96 122285
rect -96 122211 96 122217
rect -96 122177 -84 122211
rect 84 122177 96 122211
rect -96 122171 96 122177
rect -152 122118 -106 122130
rect -152 121342 -146 122118
rect -112 121342 -106 122118
rect -152 121330 -106 121342
rect 106 122118 152 122130
rect 106 121342 112 122118
rect 146 121342 152 122118
rect 106 121330 152 121342
rect -96 121283 96 121289
rect -96 121249 -84 121283
rect 84 121249 96 121283
rect -96 121243 96 121249
rect -96 121175 96 121181
rect -96 121141 -84 121175
rect 84 121141 96 121175
rect -96 121135 96 121141
rect -152 121082 -106 121094
rect -152 120306 -146 121082
rect -112 120306 -106 121082
rect -152 120294 -106 120306
rect 106 121082 152 121094
rect 106 120306 112 121082
rect 146 120306 152 121082
rect 106 120294 152 120306
rect -96 120247 96 120253
rect -96 120213 -84 120247
rect 84 120213 96 120247
rect -96 120207 96 120213
rect -96 120139 96 120145
rect -96 120105 -84 120139
rect 84 120105 96 120139
rect -96 120099 96 120105
rect -152 120046 -106 120058
rect -152 119270 -146 120046
rect -112 119270 -106 120046
rect -152 119258 -106 119270
rect 106 120046 152 120058
rect 106 119270 112 120046
rect 146 119270 152 120046
rect 106 119258 152 119270
rect -96 119211 96 119217
rect -96 119177 -84 119211
rect 84 119177 96 119211
rect -96 119171 96 119177
rect -96 119103 96 119109
rect -96 119069 -84 119103
rect 84 119069 96 119103
rect -96 119063 96 119069
rect -152 119010 -106 119022
rect -152 118234 -146 119010
rect -112 118234 -106 119010
rect -152 118222 -106 118234
rect 106 119010 152 119022
rect 106 118234 112 119010
rect 146 118234 152 119010
rect 106 118222 152 118234
rect -96 118175 96 118181
rect -96 118141 -84 118175
rect 84 118141 96 118175
rect -96 118135 96 118141
rect -96 118067 96 118073
rect -96 118033 -84 118067
rect 84 118033 96 118067
rect -96 118027 96 118033
rect -152 117974 -106 117986
rect -152 117198 -146 117974
rect -112 117198 -106 117974
rect -152 117186 -106 117198
rect 106 117974 152 117986
rect 106 117198 112 117974
rect 146 117198 152 117974
rect 106 117186 152 117198
rect -96 117139 96 117145
rect -96 117105 -84 117139
rect 84 117105 96 117139
rect -96 117099 96 117105
rect -96 117031 96 117037
rect -96 116997 -84 117031
rect 84 116997 96 117031
rect -96 116991 96 116997
rect -152 116938 -106 116950
rect -152 116162 -146 116938
rect -112 116162 -106 116938
rect -152 116150 -106 116162
rect 106 116938 152 116950
rect 106 116162 112 116938
rect 146 116162 152 116938
rect 106 116150 152 116162
rect -96 116103 96 116109
rect -96 116069 -84 116103
rect 84 116069 96 116103
rect -96 116063 96 116069
rect -96 115995 96 116001
rect -96 115961 -84 115995
rect 84 115961 96 115995
rect -96 115955 96 115961
rect -152 115902 -106 115914
rect -152 115126 -146 115902
rect -112 115126 -106 115902
rect -152 115114 -106 115126
rect 106 115902 152 115914
rect 106 115126 112 115902
rect 146 115126 152 115902
rect 106 115114 152 115126
rect -96 115067 96 115073
rect -96 115033 -84 115067
rect 84 115033 96 115067
rect -96 115027 96 115033
rect -96 114959 96 114965
rect -96 114925 -84 114959
rect 84 114925 96 114959
rect -96 114919 96 114925
rect -152 114866 -106 114878
rect -152 114090 -146 114866
rect -112 114090 -106 114866
rect -152 114078 -106 114090
rect 106 114866 152 114878
rect 106 114090 112 114866
rect 146 114090 152 114866
rect 106 114078 152 114090
rect -96 114031 96 114037
rect -96 113997 -84 114031
rect 84 113997 96 114031
rect -96 113991 96 113997
rect -96 113923 96 113929
rect -96 113889 -84 113923
rect 84 113889 96 113923
rect -96 113883 96 113889
rect -152 113830 -106 113842
rect -152 113054 -146 113830
rect -112 113054 -106 113830
rect -152 113042 -106 113054
rect 106 113830 152 113842
rect 106 113054 112 113830
rect 146 113054 152 113830
rect 106 113042 152 113054
rect -96 112995 96 113001
rect -96 112961 -84 112995
rect 84 112961 96 112995
rect -96 112955 96 112961
rect -96 112887 96 112893
rect -96 112853 -84 112887
rect 84 112853 96 112887
rect -96 112847 96 112853
rect -152 112794 -106 112806
rect -152 112018 -146 112794
rect -112 112018 -106 112794
rect -152 112006 -106 112018
rect 106 112794 152 112806
rect 106 112018 112 112794
rect 146 112018 152 112794
rect 106 112006 152 112018
rect -96 111959 96 111965
rect -96 111925 -84 111959
rect 84 111925 96 111959
rect -96 111919 96 111925
rect -96 111851 96 111857
rect -96 111817 -84 111851
rect 84 111817 96 111851
rect -96 111811 96 111817
rect -152 111758 -106 111770
rect -152 110982 -146 111758
rect -112 110982 -106 111758
rect -152 110970 -106 110982
rect 106 111758 152 111770
rect 106 110982 112 111758
rect 146 110982 152 111758
rect 106 110970 152 110982
rect -96 110923 96 110929
rect -96 110889 -84 110923
rect 84 110889 96 110923
rect -96 110883 96 110889
rect -96 110815 96 110821
rect -96 110781 -84 110815
rect 84 110781 96 110815
rect -96 110775 96 110781
rect -152 110722 -106 110734
rect -152 109946 -146 110722
rect -112 109946 -106 110722
rect -152 109934 -106 109946
rect 106 110722 152 110734
rect 106 109946 112 110722
rect 146 109946 152 110722
rect 106 109934 152 109946
rect -96 109887 96 109893
rect -96 109853 -84 109887
rect 84 109853 96 109887
rect -96 109847 96 109853
rect -96 109779 96 109785
rect -96 109745 -84 109779
rect 84 109745 96 109779
rect -96 109739 96 109745
rect -152 109686 -106 109698
rect -152 108910 -146 109686
rect -112 108910 -106 109686
rect -152 108898 -106 108910
rect 106 109686 152 109698
rect 106 108910 112 109686
rect 146 108910 152 109686
rect 106 108898 152 108910
rect -96 108851 96 108857
rect -96 108817 -84 108851
rect 84 108817 96 108851
rect -96 108811 96 108817
rect -96 108743 96 108749
rect -96 108709 -84 108743
rect 84 108709 96 108743
rect -96 108703 96 108709
rect -152 108650 -106 108662
rect -152 107874 -146 108650
rect -112 107874 -106 108650
rect -152 107862 -106 107874
rect 106 108650 152 108662
rect 106 107874 112 108650
rect 146 107874 152 108650
rect 106 107862 152 107874
rect -96 107815 96 107821
rect -96 107781 -84 107815
rect 84 107781 96 107815
rect -96 107775 96 107781
rect -96 107707 96 107713
rect -96 107673 -84 107707
rect 84 107673 96 107707
rect -96 107667 96 107673
rect -152 107614 -106 107626
rect -152 106838 -146 107614
rect -112 106838 -106 107614
rect -152 106826 -106 106838
rect 106 107614 152 107626
rect 106 106838 112 107614
rect 146 106838 152 107614
rect 106 106826 152 106838
rect -96 106779 96 106785
rect -96 106745 -84 106779
rect 84 106745 96 106779
rect -96 106739 96 106745
rect -96 106671 96 106677
rect -96 106637 -84 106671
rect 84 106637 96 106671
rect -96 106631 96 106637
rect -152 106578 -106 106590
rect -152 105802 -146 106578
rect -112 105802 -106 106578
rect -152 105790 -106 105802
rect 106 106578 152 106590
rect 106 105802 112 106578
rect 146 105802 152 106578
rect 106 105790 152 105802
rect -96 105743 96 105749
rect -96 105709 -84 105743
rect 84 105709 96 105743
rect -96 105703 96 105709
rect -96 105635 96 105641
rect -96 105601 -84 105635
rect 84 105601 96 105635
rect -96 105595 96 105601
rect -152 105542 -106 105554
rect -152 104766 -146 105542
rect -112 104766 -106 105542
rect -152 104754 -106 104766
rect 106 105542 152 105554
rect 106 104766 112 105542
rect 146 104766 152 105542
rect 106 104754 152 104766
rect -96 104707 96 104713
rect -96 104673 -84 104707
rect 84 104673 96 104707
rect -96 104667 96 104673
rect -96 104599 96 104605
rect -96 104565 -84 104599
rect 84 104565 96 104599
rect -96 104559 96 104565
rect -152 104506 -106 104518
rect -152 103730 -146 104506
rect -112 103730 -106 104506
rect -152 103718 -106 103730
rect 106 104506 152 104518
rect 106 103730 112 104506
rect 146 103730 152 104506
rect 106 103718 152 103730
rect -96 103671 96 103677
rect -96 103637 -84 103671
rect 84 103637 96 103671
rect -96 103631 96 103637
rect -96 103563 96 103569
rect -96 103529 -84 103563
rect 84 103529 96 103563
rect -96 103523 96 103529
rect -152 103470 -106 103482
rect -152 102694 -146 103470
rect -112 102694 -106 103470
rect -152 102682 -106 102694
rect 106 103470 152 103482
rect 106 102694 112 103470
rect 146 102694 152 103470
rect 106 102682 152 102694
rect -96 102635 96 102641
rect -96 102601 -84 102635
rect 84 102601 96 102635
rect -96 102595 96 102601
rect -96 102527 96 102533
rect -96 102493 -84 102527
rect 84 102493 96 102527
rect -96 102487 96 102493
rect -152 102434 -106 102446
rect -152 101658 -146 102434
rect -112 101658 -106 102434
rect -152 101646 -106 101658
rect 106 102434 152 102446
rect 106 101658 112 102434
rect 146 101658 152 102434
rect 106 101646 152 101658
rect -96 101599 96 101605
rect -96 101565 -84 101599
rect 84 101565 96 101599
rect -96 101559 96 101565
rect -96 101491 96 101497
rect -96 101457 -84 101491
rect 84 101457 96 101491
rect -96 101451 96 101457
rect -152 101398 -106 101410
rect -152 100622 -146 101398
rect -112 100622 -106 101398
rect -152 100610 -106 100622
rect 106 101398 152 101410
rect 106 100622 112 101398
rect 146 100622 152 101398
rect 106 100610 152 100622
rect -96 100563 96 100569
rect -96 100529 -84 100563
rect 84 100529 96 100563
rect -96 100523 96 100529
rect -96 100455 96 100461
rect -96 100421 -84 100455
rect 84 100421 96 100455
rect -96 100415 96 100421
rect -152 100362 -106 100374
rect -152 99586 -146 100362
rect -112 99586 -106 100362
rect -152 99574 -106 99586
rect 106 100362 152 100374
rect 106 99586 112 100362
rect 146 99586 152 100362
rect 106 99574 152 99586
rect -96 99527 96 99533
rect -96 99493 -84 99527
rect 84 99493 96 99527
rect -96 99487 96 99493
rect -96 99419 96 99425
rect -96 99385 -84 99419
rect 84 99385 96 99419
rect -96 99379 96 99385
rect -152 99326 -106 99338
rect -152 98550 -146 99326
rect -112 98550 -106 99326
rect -152 98538 -106 98550
rect 106 99326 152 99338
rect 106 98550 112 99326
rect 146 98550 152 99326
rect 106 98538 152 98550
rect -96 98491 96 98497
rect -96 98457 -84 98491
rect 84 98457 96 98491
rect -96 98451 96 98457
rect -96 98383 96 98389
rect -96 98349 -84 98383
rect 84 98349 96 98383
rect -96 98343 96 98349
rect -152 98290 -106 98302
rect -152 97514 -146 98290
rect -112 97514 -106 98290
rect -152 97502 -106 97514
rect 106 98290 152 98302
rect 106 97514 112 98290
rect 146 97514 152 98290
rect 106 97502 152 97514
rect -96 97455 96 97461
rect -96 97421 -84 97455
rect 84 97421 96 97455
rect -96 97415 96 97421
rect -96 97347 96 97353
rect -96 97313 -84 97347
rect 84 97313 96 97347
rect -96 97307 96 97313
rect -152 97254 -106 97266
rect -152 96478 -146 97254
rect -112 96478 -106 97254
rect -152 96466 -106 96478
rect 106 97254 152 97266
rect 106 96478 112 97254
rect 146 96478 152 97254
rect 106 96466 152 96478
rect -96 96419 96 96425
rect -96 96385 -84 96419
rect 84 96385 96 96419
rect -96 96379 96 96385
rect -96 96311 96 96317
rect -96 96277 -84 96311
rect 84 96277 96 96311
rect -96 96271 96 96277
rect -152 96218 -106 96230
rect -152 95442 -146 96218
rect -112 95442 -106 96218
rect -152 95430 -106 95442
rect 106 96218 152 96230
rect 106 95442 112 96218
rect 146 95442 152 96218
rect 106 95430 152 95442
rect -96 95383 96 95389
rect -96 95349 -84 95383
rect 84 95349 96 95383
rect -96 95343 96 95349
rect -96 95275 96 95281
rect -96 95241 -84 95275
rect 84 95241 96 95275
rect -96 95235 96 95241
rect -152 95182 -106 95194
rect -152 94406 -146 95182
rect -112 94406 -106 95182
rect -152 94394 -106 94406
rect 106 95182 152 95194
rect 106 94406 112 95182
rect 146 94406 152 95182
rect 106 94394 152 94406
rect -96 94347 96 94353
rect -96 94313 -84 94347
rect 84 94313 96 94347
rect -96 94307 96 94313
rect -96 94239 96 94245
rect -96 94205 -84 94239
rect 84 94205 96 94239
rect -96 94199 96 94205
rect -152 94146 -106 94158
rect -152 93370 -146 94146
rect -112 93370 -106 94146
rect -152 93358 -106 93370
rect 106 94146 152 94158
rect 106 93370 112 94146
rect 146 93370 152 94146
rect 106 93358 152 93370
rect -96 93311 96 93317
rect -96 93277 -84 93311
rect 84 93277 96 93311
rect -96 93271 96 93277
rect -96 93203 96 93209
rect -96 93169 -84 93203
rect 84 93169 96 93203
rect -96 93163 96 93169
rect -152 93110 -106 93122
rect -152 92334 -146 93110
rect -112 92334 -106 93110
rect -152 92322 -106 92334
rect 106 93110 152 93122
rect 106 92334 112 93110
rect 146 92334 152 93110
rect 106 92322 152 92334
rect -96 92275 96 92281
rect -96 92241 -84 92275
rect 84 92241 96 92275
rect -96 92235 96 92241
rect -96 92167 96 92173
rect -96 92133 -84 92167
rect 84 92133 96 92167
rect -96 92127 96 92133
rect -152 92074 -106 92086
rect -152 91298 -146 92074
rect -112 91298 -106 92074
rect -152 91286 -106 91298
rect 106 92074 152 92086
rect 106 91298 112 92074
rect 146 91298 152 92074
rect 106 91286 152 91298
rect -96 91239 96 91245
rect -96 91205 -84 91239
rect 84 91205 96 91239
rect -96 91199 96 91205
rect -96 91131 96 91137
rect -96 91097 -84 91131
rect 84 91097 96 91131
rect -96 91091 96 91097
rect -152 91038 -106 91050
rect -152 90262 -146 91038
rect -112 90262 -106 91038
rect -152 90250 -106 90262
rect 106 91038 152 91050
rect 106 90262 112 91038
rect 146 90262 152 91038
rect 106 90250 152 90262
rect -96 90203 96 90209
rect -96 90169 -84 90203
rect 84 90169 96 90203
rect -96 90163 96 90169
rect -96 90095 96 90101
rect -96 90061 -84 90095
rect 84 90061 96 90095
rect -96 90055 96 90061
rect -152 90002 -106 90014
rect -152 89226 -146 90002
rect -112 89226 -106 90002
rect -152 89214 -106 89226
rect 106 90002 152 90014
rect 106 89226 112 90002
rect 146 89226 152 90002
rect 106 89214 152 89226
rect -96 89167 96 89173
rect -96 89133 -84 89167
rect 84 89133 96 89167
rect -96 89127 96 89133
rect -96 89059 96 89065
rect -96 89025 -84 89059
rect 84 89025 96 89059
rect -96 89019 96 89025
rect -152 88966 -106 88978
rect -152 88190 -146 88966
rect -112 88190 -106 88966
rect -152 88178 -106 88190
rect 106 88966 152 88978
rect 106 88190 112 88966
rect 146 88190 152 88966
rect 106 88178 152 88190
rect -96 88131 96 88137
rect -96 88097 -84 88131
rect 84 88097 96 88131
rect -96 88091 96 88097
rect -96 88023 96 88029
rect -96 87989 -84 88023
rect 84 87989 96 88023
rect -96 87983 96 87989
rect -152 87930 -106 87942
rect -152 87154 -146 87930
rect -112 87154 -106 87930
rect -152 87142 -106 87154
rect 106 87930 152 87942
rect 106 87154 112 87930
rect 146 87154 152 87930
rect 106 87142 152 87154
rect -96 87095 96 87101
rect -96 87061 -84 87095
rect 84 87061 96 87095
rect -96 87055 96 87061
rect -96 86987 96 86993
rect -96 86953 -84 86987
rect 84 86953 96 86987
rect -96 86947 96 86953
rect -152 86894 -106 86906
rect -152 86118 -146 86894
rect -112 86118 -106 86894
rect -152 86106 -106 86118
rect 106 86894 152 86906
rect 106 86118 112 86894
rect 146 86118 152 86894
rect 106 86106 152 86118
rect -96 86059 96 86065
rect -96 86025 -84 86059
rect 84 86025 96 86059
rect -96 86019 96 86025
rect -96 85951 96 85957
rect -96 85917 -84 85951
rect 84 85917 96 85951
rect -96 85911 96 85917
rect -152 85858 -106 85870
rect -152 85082 -146 85858
rect -112 85082 -106 85858
rect -152 85070 -106 85082
rect 106 85858 152 85870
rect 106 85082 112 85858
rect 146 85082 152 85858
rect 106 85070 152 85082
rect -96 85023 96 85029
rect -96 84989 -84 85023
rect 84 84989 96 85023
rect -96 84983 96 84989
rect -96 84915 96 84921
rect -96 84881 -84 84915
rect 84 84881 96 84915
rect -96 84875 96 84881
rect -152 84822 -106 84834
rect -152 84046 -146 84822
rect -112 84046 -106 84822
rect -152 84034 -106 84046
rect 106 84822 152 84834
rect 106 84046 112 84822
rect 146 84046 152 84822
rect 106 84034 152 84046
rect -96 83987 96 83993
rect -96 83953 -84 83987
rect 84 83953 96 83987
rect -96 83947 96 83953
rect -96 83879 96 83885
rect -96 83845 -84 83879
rect 84 83845 96 83879
rect -96 83839 96 83845
rect -152 83786 -106 83798
rect -152 83010 -146 83786
rect -112 83010 -106 83786
rect -152 82998 -106 83010
rect 106 83786 152 83798
rect 106 83010 112 83786
rect 146 83010 152 83786
rect 106 82998 152 83010
rect -96 82951 96 82957
rect -96 82917 -84 82951
rect 84 82917 96 82951
rect -96 82911 96 82917
rect -96 82843 96 82849
rect -96 82809 -84 82843
rect 84 82809 96 82843
rect -96 82803 96 82809
rect -152 82750 -106 82762
rect -152 81974 -146 82750
rect -112 81974 -106 82750
rect -152 81962 -106 81974
rect 106 82750 152 82762
rect 106 81974 112 82750
rect 146 81974 152 82750
rect 106 81962 152 81974
rect -96 81915 96 81921
rect -96 81881 -84 81915
rect 84 81881 96 81915
rect -96 81875 96 81881
rect -96 81807 96 81813
rect -96 81773 -84 81807
rect 84 81773 96 81807
rect -96 81767 96 81773
rect -152 81714 -106 81726
rect -152 80938 -146 81714
rect -112 80938 -106 81714
rect -152 80926 -106 80938
rect 106 81714 152 81726
rect 106 80938 112 81714
rect 146 80938 152 81714
rect 106 80926 152 80938
rect -96 80879 96 80885
rect -96 80845 -84 80879
rect 84 80845 96 80879
rect -96 80839 96 80845
rect -96 80771 96 80777
rect -96 80737 -84 80771
rect 84 80737 96 80771
rect -96 80731 96 80737
rect -152 80678 -106 80690
rect -152 79902 -146 80678
rect -112 79902 -106 80678
rect -152 79890 -106 79902
rect 106 80678 152 80690
rect 106 79902 112 80678
rect 146 79902 152 80678
rect 106 79890 152 79902
rect -96 79843 96 79849
rect -96 79809 -84 79843
rect 84 79809 96 79843
rect -96 79803 96 79809
rect -96 79735 96 79741
rect -96 79701 -84 79735
rect 84 79701 96 79735
rect -96 79695 96 79701
rect -152 79642 -106 79654
rect -152 78866 -146 79642
rect -112 78866 -106 79642
rect -152 78854 -106 78866
rect 106 79642 152 79654
rect 106 78866 112 79642
rect 146 78866 152 79642
rect 106 78854 152 78866
rect -96 78807 96 78813
rect -96 78773 -84 78807
rect 84 78773 96 78807
rect -96 78767 96 78773
rect -96 78699 96 78705
rect -96 78665 -84 78699
rect 84 78665 96 78699
rect -96 78659 96 78665
rect -152 78606 -106 78618
rect -152 77830 -146 78606
rect -112 77830 -106 78606
rect -152 77818 -106 77830
rect 106 78606 152 78618
rect 106 77830 112 78606
rect 146 77830 152 78606
rect 106 77818 152 77830
rect -96 77771 96 77777
rect -96 77737 -84 77771
rect 84 77737 96 77771
rect -96 77731 96 77737
rect -96 77663 96 77669
rect -96 77629 -84 77663
rect 84 77629 96 77663
rect -96 77623 96 77629
rect -152 77570 -106 77582
rect -152 76794 -146 77570
rect -112 76794 -106 77570
rect -152 76782 -106 76794
rect 106 77570 152 77582
rect 106 76794 112 77570
rect 146 76794 152 77570
rect 106 76782 152 76794
rect -96 76735 96 76741
rect -96 76701 -84 76735
rect 84 76701 96 76735
rect -96 76695 96 76701
rect -96 76627 96 76633
rect -96 76593 -84 76627
rect 84 76593 96 76627
rect -96 76587 96 76593
rect -152 76534 -106 76546
rect -152 75758 -146 76534
rect -112 75758 -106 76534
rect -152 75746 -106 75758
rect 106 76534 152 76546
rect 106 75758 112 76534
rect 146 75758 152 76534
rect 106 75746 152 75758
rect -96 75699 96 75705
rect -96 75665 -84 75699
rect 84 75665 96 75699
rect -96 75659 96 75665
rect -96 75591 96 75597
rect -96 75557 -84 75591
rect 84 75557 96 75591
rect -96 75551 96 75557
rect -152 75498 -106 75510
rect -152 74722 -146 75498
rect -112 74722 -106 75498
rect -152 74710 -106 74722
rect 106 75498 152 75510
rect 106 74722 112 75498
rect 146 74722 152 75498
rect 106 74710 152 74722
rect -96 74663 96 74669
rect -96 74629 -84 74663
rect 84 74629 96 74663
rect -96 74623 96 74629
rect -96 74555 96 74561
rect -96 74521 -84 74555
rect 84 74521 96 74555
rect -96 74515 96 74521
rect -152 74462 -106 74474
rect -152 73686 -146 74462
rect -112 73686 -106 74462
rect -152 73674 -106 73686
rect 106 74462 152 74474
rect 106 73686 112 74462
rect 146 73686 152 74462
rect 106 73674 152 73686
rect -96 73627 96 73633
rect -96 73593 -84 73627
rect 84 73593 96 73627
rect -96 73587 96 73593
rect -96 73519 96 73525
rect -96 73485 -84 73519
rect 84 73485 96 73519
rect -96 73479 96 73485
rect -152 73426 -106 73438
rect -152 72650 -146 73426
rect -112 72650 -106 73426
rect -152 72638 -106 72650
rect 106 73426 152 73438
rect 106 72650 112 73426
rect 146 72650 152 73426
rect 106 72638 152 72650
rect -96 72591 96 72597
rect -96 72557 -84 72591
rect 84 72557 96 72591
rect -96 72551 96 72557
rect -96 72483 96 72489
rect -96 72449 -84 72483
rect 84 72449 96 72483
rect -96 72443 96 72449
rect -152 72390 -106 72402
rect -152 71614 -146 72390
rect -112 71614 -106 72390
rect -152 71602 -106 71614
rect 106 72390 152 72402
rect 106 71614 112 72390
rect 146 71614 152 72390
rect 106 71602 152 71614
rect -96 71555 96 71561
rect -96 71521 -84 71555
rect 84 71521 96 71555
rect -96 71515 96 71521
rect -96 71447 96 71453
rect -96 71413 -84 71447
rect 84 71413 96 71447
rect -96 71407 96 71413
rect -152 71354 -106 71366
rect -152 70578 -146 71354
rect -112 70578 -106 71354
rect -152 70566 -106 70578
rect 106 71354 152 71366
rect 106 70578 112 71354
rect 146 70578 152 71354
rect 106 70566 152 70578
rect -96 70519 96 70525
rect -96 70485 -84 70519
rect 84 70485 96 70519
rect -96 70479 96 70485
rect -96 70411 96 70417
rect -96 70377 -84 70411
rect 84 70377 96 70411
rect -96 70371 96 70377
rect -152 70318 -106 70330
rect -152 69542 -146 70318
rect -112 69542 -106 70318
rect -152 69530 -106 69542
rect 106 70318 152 70330
rect 106 69542 112 70318
rect 146 69542 152 70318
rect 106 69530 152 69542
rect -96 69483 96 69489
rect -96 69449 -84 69483
rect 84 69449 96 69483
rect -96 69443 96 69449
rect -96 69375 96 69381
rect -96 69341 -84 69375
rect 84 69341 96 69375
rect -96 69335 96 69341
rect -152 69282 -106 69294
rect -152 68506 -146 69282
rect -112 68506 -106 69282
rect -152 68494 -106 68506
rect 106 69282 152 69294
rect 106 68506 112 69282
rect 146 68506 152 69282
rect 106 68494 152 68506
rect -96 68447 96 68453
rect -96 68413 -84 68447
rect 84 68413 96 68447
rect -96 68407 96 68413
rect -96 68339 96 68345
rect -96 68305 -84 68339
rect 84 68305 96 68339
rect -96 68299 96 68305
rect -152 68246 -106 68258
rect -152 67470 -146 68246
rect -112 67470 -106 68246
rect -152 67458 -106 67470
rect 106 68246 152 68258
rect 106 67470 112 68246
rect 146 67470 152 68246
rect 106 67458 152 67470
rect -96 67411 96 67417
rect -96 67377 -84 67411
rect 84 67377 96 67411
rect -96 67371 96 67377
rect -96 67303 96 67309
rect -96 67269 -84 67303
rect 84 67269 96 67303
rect -96 67263 96 67269
rect -152 67210 -106 67222
rect -152 66434 -146 67210
rect -112 66434 -106 67210
rect -152 66422 -106 66434
rect 106 67210 152 67222
rect 106 66434 112 67210
rect 146 66434 152 67210
rect 106 66422 152 66434
rect -96 66375 96 66381
rect -96 66341 -84 66375
rect 84 66341 96 66375
rect -96 66335 96 66341
rect -96 66267 96 66273
rect -96 66233 -84 66267
rect 84 66233 96 66267
rect -96 66227 96 66233
rect -152 66174 -106 66186
rect -152 65398 -146 66174
rect -112 65398 -106 66174
rect -152 65386 -106 65398
rect 106 66174 152 66186
rect 106 65398 112 66174
rect 146 65398 152 66174
rect 106 65386 152 65398
rect -96 65339 96 65345
rect -96 65305 -84 65339
rect 84 65305 96 65339
rect -96 65299 96 65305
rect -96 65231 96 65237
rect -96 65197 -84 65231
rect 84 65197 96 65231
rect -96 65191 96 65197
rect -152 65138 -106 65150
rect -152 64362 -146 65138
rect -112 64362 -106 65138
rect -152 64350 -106 64362
rect 106 65138 152 65150
rect 106 64362 112 65138
rect 146 64362 152 65138
rect 106 64350 152 64362
rect -96 64303 96 64309
rect -96 64269 -84 64303
rect 84 64269 96 64303
rect -96 64263 96 64269
rect -96 64195 96 64201
rect -96 64161 -84 64195
rect 84 64161 96 64195
rect -96 64155 96 64161
rect -152 64102 -106 64114
rect -152 63326 -146 64102
rect -112 63326 -106 64102
rect -152 63314 -106 63326
rect 106 64102 152 64114
rect 106 63326 112 64102
rect 146 63326 152 64102
rect 106 63314 152 63326
rect -96 63267 96 63273
rect -96 63233 -84 63267
rect 84 63233 96 63267
rect -96 63227 96 63233
rect -96 63159 96 63165
rect -96 63125 -84 63159
rect 84 63125 96 63159
rect -96 63119 96 63125
rect -152 63066 -106 63078
rect -152 62290 -146 63066
rect -112 62290 -106 63066
rect -152 62278 -106 62290
rect 106 63066 152 63078
rect 106 62290 112 63066
rect 146 62290 152 63066
rect 106 62278 152 62290
rect -96 62231 96 62237
rect -96 62197 -84 62231
rect 84 62197 96 62231
rect -96 62191 96 62197
rect -96 62123 96 62129
rect -96 62089 -84 62123
rect 84 62089 96 62123
rect -96 62083 96 62089
rect -152 62030 -106 62042
rect -152 61254 -146 62030
rect -112 61254 -106 62030
rect -152 61242 -106 61254
rect 106 62030 152 62042
rect 106 61254 112 62030
rect 146 61254 152 62030
rect 106 61242 152 61254
rect -96 61195 96 61201
rect -96 61161 -84 61195
rect 84 61161 96 61195
rect -96 61155 96 61161
rect -96 61087 96 61093
rect -96 61053 -84 61087
rect 84 61053 96 61087
rect -96 61047 96 61053
rect -152 60994 -106 61006
rect -152 60218 -146 60994
rect -112 60218 -106 60994
rect -152 60206 -106 60218
rect 106 60994 152 61006
rect 106 60218 112 60994
rect 146 60218 152 60994
rect 106 60206 152 60218
rect -96 60159 96 60165
rect -96 60125 -84 60159
rect 84 60125 96 60159
rect -96 60119 96 60125
rect -96 60051 96 60057
rect -96 60017 -84 60051
rect 84 60017 96 60051
rect -96 60011 96 60017
rect -152 59958 -106 59970
rect -152 59182 -146 59958
rect -112 59182 -106 59958
rect -152 59170 -106 59182
rect 106 59958 152 59970
rect 106 59182 112 59958
rect 146 59182 152 59958
rect 106 59170 152 59182
rect -96 59123 96 59129
rect -96 59089 -84 59123
rect 84 59089 96 59123
rect -96 59083 96 59089
rect -96 59015 96 59021
rect -96 58981 -84 59015
rect 84 58981 96 59015
rect -96 58975 96 58981
rect -152 58922 -106 58934
rect -152 58146 -146 58922
rect -112 58146 -106 58922
rect -152 58134 -106 58146
rect 106 58922 152 58934
rect 106 58146 112 58922
rect 146 58146 152 58922
rect 106 58134 152 58146
rect -96 58087 96 58093
rect -96 58053 -84 58087
rect 84 58053 96 58087
rect -96 58047 96 58053
rect -96 57979 96 57985
rect -96 57945 -84 57979
rect 84 57945 96 57979
rect -96 57939 96 57945
rect -152 57886 -106 57898
rect -152 57110 -146 57886
rect -112 57110 -106 57886
rect -152 57098 -106 57110
rect 106 57886 152 57898
rect 106 57110 112 57886
rect 146 57110 152 57886
rect 106 57098 152 57110
rect -96 57051 96 57057
rect -96 57017 -84 57051
rect 84 57017 96 57051
rect -96 57011 96 57017
rect -96 56943 96 56949
rect -96 56909 -84 56943
rect 84 56909 96 56943
rect -96 56903 96 56909
rect -152 56850 -106 56862
rect -152 56074 -146 56850
rect -112 56074 -106 56850
rect -152 56062 -106 56074
rect 106 56850 152 56862
rect 106 56074 112 56850
rect 146 56074 152 56850
rect 106 56062 152 56074
rect -96 56015 96 56021
rect -96 55981 -84 56015
rect 84 55981 96 56015
rect -96 55975 96 55981
rect -96 55907 96 55913
rect -96 55873 -84 55907
rect 84 55873 96 55907
rect -96 55867 96 55873
rect -152 55814 -106 55826
rect -152 55038 -146 55814
rect -112 55038 -106 55814
rect -152 55026 -106 55038
rect 106 55814 152 55826
rect 106 55038 112 55814
rect 146 55038 152 55814
rect 106 55026 152 55038
rect -96 54979 96 54985
rect -96 54945 -84 54979
rect 84 54945 96 54979
rect -96 54939 96 54945
rect -96 54871 96 54877
rect -96 54837 -84 54871
rect 84 54837 96 54871
rect -96 54831 96 54837
rect -152 54778 -106 54790
rect -152 54002 -146 54778
rect -112 54002 -106 54778
rect -152 53990 -106 54002
rect 106 54778 152 54790
rect 106 54002 112 54778
rect 146 54002 152 54778
rect 106 53990 152 54002
rect -96 53943 96 53949
rect -96 53909 -84 53943
rect 84 53909 96 53943
rect -96 53903 96 53909
rect -96 53835 96 53841
rect -96 53801 -84 53835
rect 84 53801 96 53835
rect -96 53795 96 53801
rect -152 53742 -106 53754
rect -152 52966 -146 53742
rect -112 52966 -106 53742
rect -152 52954 -106 52966
rect 106 53742 152 53754
rect 106 52966 112 53742
rect 146 52966 152 53742
rect 106 52954 152 52966
rect -96 52907 96 52913
rect -96 52873 -84 52907
rect 84 52873 96 52907
rect -96 52867 96 52873
rect -96 52799 96 52805
rect -96 52765 -84 52799
rect 84 52765 96 52799
rect -96 52759 96 52765
rect -152 52706 -106 52718
rect -152 51930 -146 52706
rect -112 51930 -106 52706
rect -152 51918 -106 51930
rect 106 52706 152 52718
rect 106 51930 112 52706
rect 146 51930 152 52706
rect 106 51918 152 51930
rect -96 51871 96 51877
rect -96 51837 -84 51871
rect 84 51837 96 51871
rect -96 51831 96 51837
rect -96 51763 96 51769
rect -96 51729 -84 51763
rect 84 51729 96 51763
rect -96 51723 96 51729
rect -152 51670 -106 51682
rect -152 50894 -146 51670
rect -112 50894 -106 51670
rect -152 50882 -106 50894
rect 106 51670 152 51682
rect 106 50894 112 51670
rect 146 50894 152 51670
rect 106 50882 152 50894
rect -96 50835 96 50841
rect -96 50801 -84 50835
rect 84 50801 96 50835
rect -96 50795 96 50801
rect -96 50727 96 50733
rect -96 50693 -84 50727
rect 84 50693 96 50727
rect -96 50687 96 50693
rect -152 50634 -106 50646
rect -152 49858 -146 50634
rect -112 49858 -106 50634
rect -152 49846 -106 49858
rect 106 50634 152 50646
rect 106 49858 112 50634
rect 146 49858 152 50634
rect 106 49846 152 49858
rect -96 49799 96 49805
rect -96 49765 -84 49799
rect 84 49765 96 49799
rect -96 49759 96 49765
rect -96 49691 96 49697
rect -96 49657 -84 49691
rect 84 49657 96 49691
rect -96 49651 96 49657
rect -152 49598 -106 49610
rect -152 48822 -146 49598
rect -112 48822 -106 49598
rect -152 48810 -106 48822
rect 106 49598 152 49610
rect 106 48822 112 49598
rect 146 48822 152 49598
rect 106 48810 152 48822
rect -96 48763 96 48769
rect -96 48729 -84 48763
rect 84 48729 96 48763
rect -96 48723 96 48729
rect -96 48655 96 48661
rect -96 48621 -84 48655
rect 84 48621 96 48655
rect -96 48615 96 48621
rect -152 48562 -106 48574
rect -152 47786 -146 48562
rect -112 47786 -106 48562
rect -152 47774 -106 47786
rect 106 48562 152 48574
rect 106 47786 112 48562
rect 146 47786 152 48562
rect 106 47774 152 47786
rect -96 47727 96 47733
rect -96 47693 -84 47727
rect 84 47693 96 47727
rect -96 47687 96 47693
rect -96 47619 96 47625
rect -96 47585 -84 47619
rect 84 47585 96 47619
rect -96 47579 96 47585
rect -152 47526 -106 47538
rect -152 46750 -146 47526
rect -112 46750 -106 47526
rect -152 46738 -106 46750
rect 106 47526 152 47538
rect 106 46750 112 47526
rect 146 46750 152 47526
rect 106 46738 152 46750
rect -96 46691 96 46697
rect -96 46657 -84 46691
rect 84 46657 96 46691
rect -96 46651 96 46657
rect -96 46583 96 46589
rect -96 46549 -84 46583
rect 84 46549 96 46583
rect -96 46543 96 46549
rect -152 46490 -106 46502
rect -152 45714 -146 46490
rect -112 45714 -106 46490
rect -152 45702 -106 45714
rect 106 46490 152 46502
rect 106 45714 112 46490
rect 146 45714 152 46490
rect 106 45702 152 45714
rect -96 45655 96 45661
rect -96 45621 -84 45655
rect 84 45621 96 45655
rect -96 45615 96 45621
rect -96 45547 96 45553
rect -96 45513 -84 45547
rect 84 45513 96 45547
rect -96 45507 96 45513
rect -152 45454 -106 45466
rect -152 44678 -146 45454
rect -112 44678 -106 45454
rect -152 44666 -106 44678
rect 106 45454 152 45466
rect 106 44678 112 45454
rect 146 44678 152 45454
rect 106 44666 152 44678
rect -96 44619 96 44625
rect -96 44585 -84 44619
rect 84 44585 96 44619
rect -96 44579 96 44585
rect -96 44511 96 44517
rect -96 44477 -84 44511
rect 84 44477 96 44511
rect -96 44471 96 44477
rect -152 44418 -106 44430
rect -152 43642 -146 44418
rect -112 43642 -106 44418
rect -152 43630 -106 43642
rect 106 44418 152 44430
rect 106 43642 112 44418
rect 146 43642 152 44418
rect 106 43630 152 43642
rect -96 43583 96 43589
rect -96 43549 -84 43583
rect 84 43549 96 43583
rect -96 43543 96 43549
rect -96 43475 96 43481
rect -96 43441 -84 43475
rect 84 43441 96 43475
rect -96 43435 96 43441
rect -152 43382 -106 43394
rect -152 42606 -146 43382
rect -112 42606 -106 43382
rect -152 42594 -106 42606
rect 106 43382 152 43394
rect 106 42606 112 43382
rect 146 42606 152 43382
rect 106 42594 152 42606
rect -96 42547 96 42553
rect -96 42513 -84 42547
rect 84 42513 96 42547
rect -96 42507 96 42513
rect -96 42439 96 42445
rect -96 42405 -84 42439
rect 84 42405 96 42439
rect -96 42399 96 42405
rect -152 42346 -106 42358
rect -152 41570 -146 42346
rect -112 41570 -106 42346
rect -152 41558 -106 41570
rect 106 42346 152 42358
rect 106 41570 112 42346
rect 146 41570 152 42346
rect 106 41558 152 41570
rect -96 41511 96 41517
rect -96 41477 -84 41511
rect 84 41477 96 41511
rect -96 41471 96 41477
rect -96 41403 96 41409
rect -96 41369 -84 41403
rect 84 41369 96 41403
rect -96 41363 96 41369
rect -152 41310 -106 41322
rect -152 40534 -146 41310
rect -112 40534 -106 41310
rect -152 40522 -106 40534
rect 106 41310 152 41322
rect 106 40534 112 41310
rect 146 40534 152 41310
rect 106 40522 152 40534
rect -96 40475 96 40481
rect -96 40441 -84 40475
rect 84 40441 96 40475
rect -96 40435 96 40441
rect -96 40367 96 40373
rect -96 40333 -84 40367
rect 84 40333 96 40367
rect -96 40327 96 40333
rect -152 40274 -106 40286
rect -152 39498 -146 40274
rect -112 39498 -106 40274
rect -152 39486 -106 39498
rect 106 40274 152 40286
rect 106 39498 112 40274
rect 146 39498 152 40274
rect 106 39486 152 39498
rect -96 39439 96 39445
rect -96 39405 -84 39439
rect 84 39405 96 39439
rect -96 39399 96 39405
rect -96 39331 96 39337
rect -96 39297 -84 39331
rect 84 39297 96 39331
rect -96 39291 96 39297
rect -152 39238 -106 39250
rect -152 38462 -146 39238
rect -112 38462 -106 39238
rect -152 38450 -106 38462
rect 106 39238 152 39250
rect 106 38462 112 39238
rect 146 38462 152 39238
rect 106 38450 152 38462
rect -96 38403 96 38409
rect -96 38369 -84 38403
rect 84 38369 96 38403
rect -96 38363 96 38369
rect -96 38295 96 38301
rect -96 38261 -84 38295
rect 84 38261 96 38295
rect -96 38255 96 38261
rect -152 38202 -106 38214
rect -152 37426 -146 38202
rect -112 37426 -106 38202
rect -152 37414 -106 37426
rect 106 38202 152 38214
rect 106 37426 112 38202
rect 146 37426 152 38202
rect 106 37414 152 37426
rect -96 37367 96 37373
rect -96 37333 -84 37367
rect 84 37333 96 37367
rect -96 37327 96 37333
rect -96 37259 96 37265
rect -96 37225 -84 37259
rect 84 37225 96 37259
rect -96 37219 96 37225
rect -152 37166 -106 37178
rect -152 36390 -146 37166
rect -112 36390 -106 37166
rect -152 36378 -106 36390
rect 106 37166 152 37178
rect 106 36390 112 37166
rect 146 36390 152 37166
rect 106 36378 152 36390
rect -96 36331 96 36337
rect -96 36297 -84 36331
rect 84 36297 96 36331
rect -96 36291 96 36297
rect -96 36223 96 36229
rect -96 36189 -84 36223
rect 84 36189 96 36223
rect -96 36183 96 36189
rect -152 36130 -106 36142
rect -152 35354 -146 36130
rect -112 35354 -106 36130
rect -152 35342 -106 35354
rect 106 36130 152 36142
rect 106 35354 112 36130
rect 146 35354 152 36130
rect 106 35342 152 35354
rect -96 35295 96 35301
rect -96 35261 -84 35295
rect 84 35261 96 35295
rect -96 35255 96 35261
rect -96 35187 96 35193
rect -96 35153 -84 35187
rect 84 35153 96 35187
rect -96 35147 96 35153
rect -152 35094 -106 35106
rect -152 34318 -146 35094
rect -112 34318 -106 35094
rect -152 34306 -106 34318
rect 106 35094 152 35106
rect 106 34318 112 35094
rect 146 34318 152 35094
rect 106 34306 152 34318
rect -96 34259 96 34265
rect -96 34225 -84 34259
rect 84 34225 96 34259
rect -96 34219 96 34225
rect -96 34151 96 34157
rect -96 34117 -84 34151
rect 84 34117 96 34151
rect -96 34111 96 34117
rect -152 34058 -106 34070
rect -152 33282 -146 34058
rect -112 33282 -106 34058
rect -152 33270 -106 33282
rect 106 34058 152 34070
rect 106 33282 112 34058
rect 146 33282 152 34058
rect 106 33270 152 33282
rect -96 33223 96 33229
rect -96 33189 -84 33223
rect 84 33189 96 33223
rect -96 33183 96 33189
rect -96 33115 96 33121
rect -96 33081 -84 33115
rect 84 33081 96 33115
rect -96 33075 96 33081
rect -152 33022 -106 33034
rect -152 32246 -146 33022
rect -112 32246 -106 33022
rect -152 32234 -106 32246
rect 106 33022 152 33034
rect 106 32246 112 33022
rect 146 32246 152 33022
rect 106 32234 152 32246
rect -96 32187 96 32193
rect -96 32153 -84 32187
rect 84 32153 96 32187
rect -96 32147 96 32153
rect -96 32079 96 32085
rect -96 32045 -84 32079
rect 84 32045 96 32079
rect -96 32039 96 32045
rect -152 31986 -106 31998
rect -152 31210 -146 31986
rect -112 31210 -106 31986
rect -152 31198 -106 31210
rect 106 31986 152 31998
rect 106 31210 112 31986
rect 146 31210 152 31986
rect 106 31198 152 31210
rect -96 31151 96 31157
rect -96 31117 -84 31151
rect 84 31117 96 31151
rect -96 31111 96 31117
rect -96 31043 96 31049
rect -96 31009 -84 31043
rect 84 31009 96 31043
rect -96 31003 96 31009
rect -152 30950 -106 30962
rect -152 30174 -146 30950
rect -112 30174 -106 30950
rect -152 30162 -106 30174
rect 106 30950 152 30962
rect 106 30174 112 30950
rect 146 30174 152 30950
rect 106 30162 152 30174
rect -96 30115 96 30121
rect -96 30081 -84 30115
rect 84 30081 96 30115
rect -96 30075 96 30081
rect -96 30007 96 30013
rect -96 29973 -84 30007
rect 84 29973 96 30007
rect -96 29967 96 29973
rect -152 29914 -106 29926
rect -152 29138 -146 29914
rect -112 29138 -106 29914
rect -152 29126 -106 29138
rect 106 29914 152 29926
rect 106 29138 112 29914
rect 146 29138 152 29914
rect 106 29126 152 29138
rect -96 29079 96 29085
rect -96 29045 -84 29079
rect 84 29045 96 29079
rect -96 29039 96 29045
rect -96 28971 96 28977
rect -96 28937 -84 28971
rect 84 28937 96 28971
rect -96 28931 96 28937
rect -152 28878 -106 28890
rect -152 28102 -146 28878
rect -112 28102 -106 28878
rect -152 28090 -106 28102
rect 106 28878 152 28890
rect 106 28102 112 28878
rect 146 28102 152 28878
rect 106 28090 152 28102
rect -96 28043 96 28049
rect -96 28009 -84 28043
rect 84 28009 96 28043
rect -96 28003 96 28009
rect -96 27935 96 27941
rect -96 27901 -84 27935
rect 84 27901 96 27935
rect -96 27895 96 27901
rect -152 27842 -106 27854
rect -152 27066 -146 27842
rect -112 27066 -106 27842
rect -152 27054 -106 27066
rect 106 27842 152 27854
rect 106 27066 112 27842
rect 146 27066 152 27842
rect 106 27054 152 27066
rect -96 27007 96 27013
rect -96 26973 -84 27007
rect 84 26973 96 27007
rect -96 26967 96 26973
rect -96 26899 96 26905
rect -96 26865 -84 26899
rect 84 26865 96 26899
rect -96 26859 96 26865
rect -152 26806 -106 26818
rect -152 26030 -146 26806
rect -112 26030 -106 26806
rect -152 26018 -106 26030
rect 106 26806 152 26818
rect 106 26030 112 26806
rect 146 26030 152 26806
rect 106 26018 152 26030
rect -96 25971 96 25977
rect -96 25937 -84 25971
rect 84 25937 96 25971
rect -96 25931 96 25937
rect -96 25863 96 25869
rect -96 25829 -84 25863
rect 84 25829 96 25863
rect -96 25823 96 25829
rect -152 25770 -106 25782
rect -152 24994 -146 25770
rect -112 24994 -106 25770
rect -152 24982 -106 24994
rect 106 25770 152 25782
rect 106 24994 112 25770
rect 146 24994 152 25770
rect 106 24982 152 24994
rect -96 24935 96 24941
rect -96 24901 -84 24935
rect 84 24901 96 24935
rect -96 24895 96 24901
rect -96 24827 96 24833
rect -96 24793 -84 24827
rect 84 24793 96 24827
rect -96 24787 96 24793
rect -152 24734 -106 24746
rect -152 23958 -146 24734
rect -112 23958 -106 24734
rect -152 23946 -106 23958
rect 106 24734 152 24746
rect 106 23958 112 24734
rect 146 23958 152 24734
rect 106 23946 152 23958
rect -96 23899 96 23905
rect -96 23865 -84 23899
rect 84 23865 96 23899
rect -96 23859 96 23865
rect -96 23791 96 23797
rect -96 23757 -84 23791
rect 84 23757 96 23791
rect -96 23751 96 23757
rect -152 23698 -106 23710
rect -152 22922 -146 23698
rect -112 22922 -106 23698
rect -152 22910 -106 22922
rect 106 23698 152 23710
rect 106 22922 112 23698
rect 146 22922 152 23698
rect 106 22910 152 22922
rect -96 22863 96 22869
rect -96 22829 -84 22863
rect 84 22829 96 22863
rect -96 22823 96 22829
rect -96 22755 96 22761
rect -96 22721 -84 22755
rect 84 22721 96 22755
rect -96 22715 96 22721
rect -152 22662 -106 22674
rect -152 21886 -146 22662
rect -112 21886 -106 22662
rect -152 21874 -106 21886
rect 106 22662 152 22674
rect 106 21886 112 22662
rect 146 21886 152 22662
rect 106 21874 152 21886
rect -96 21827 96 21833
rect -96 21793 -84 21827
rect 84 21793 96 21827
rect -96 21787 96 21793
rect -96 21719 96 21725
rect -96 21685 -84 21719
rect 84 21685 96 21719
rect -96 21679 96 21685
rect -152 21626 -106 21638
rect -152 20850 -146 21626
rect -112 20850 -106 21626
rect -152 20838 -106 20850
rect 106 21626 152 21638
rect 106 20850 112 21626
rect 146 20850 152 21626
rect 106 20838 152 20850
rect -96 20791 96 20797
rect -96 20757 -84 20791
rect 84 20757 96 20791
rect -96 20751 96 20757
rect -96 20683 96 20689
rect -96 20649 -84 20683
rect 84 20649 96 20683
rect -96 20643 96 20649
rect -152 20590 -106 20602
rect -152 19814 -146 20590
rect -112 19814 -106 20590
rect -152 19802 -106 19814
rect 106 20590 152 20602
rect 106 19814 112 20590
rect 146 19814 152 20590
rect 106 19802 152 19814
rect -96 19755 96 19761
rect -96 19721 -84 19755
rect 84 19721 96 19755
rect -96 19715 96 19721
rect -96 19647 96 19653
rect -96 19613 -84 19647
rect 84 19613 96 19647
rect -96 19607 96 19613
rect -152 19554 -106 19566
rect -152 18778 -146 19554
rect -112 18778 -106 19554
rect -152 18766 -106 18778
rect 106 19554 152 19566
rect 106 18778 112 19554
rect 146 18778 152 19554
rect 106 18766 152 18778
rect -96 18719 96 18725
rect -96 18685 -84 18719
rect 84 18685 96 18719
rect -96 18679 96 18685
rect -96 18611 96 18617
rect -96 18577 -84 18611
rect 84 18577 96 18611
rect -96 18571 96 18577
rect -152 18518 -106 18530
rect -152 17742 -146 18518
rect -112 17742 -106 18518
rect -152 17730 -106 17742
rect 106 18518 152 18530
rect 106 17742 112 18518
rect 146 17742 152 18518
rect 106 17730 152 17742
rect -96 17683 96 17689
rect -96 17649 -84 17683
rect 84 17649 96 17683
rect -96 17643 96 17649
rect -96 17575 96 17581
rect -96 17541 -84 17575
rect 84 17541 96 17575
rect -96 17535 96 17541
rect -152 17482 -106 17494
rect -152 16706 -146 17482
rect -112 16706 -106 17482
rect -152 16694 -106 16706
rect 106 17482 152 17494
rect 106 16706 112 17482
rect 146 16706 152 17482
rect 106 16694 152 16706
rect -96 16647 96 16653
rect -96 16613 -84 16647
rect 84 16613 96 16647
rect -96 16607 96 16613
rect -96 16539 96 16545
rect -96 16505 -84 16539
rect 84 16505 96 16539
rect -96 16499 96 16505
rect -152 16446 -106 16458
rect -152 15670 -146 16446
rect -112 15670 -106 16446
rect -152 15658 -106 15670
rect 106 16446 152 16458
rect 106 15670 112 16446
rect 146 15670 152 16446
rect 106 15658 152 15670
rect -96 15611 96 15617
rect -96 15577 -84 15611
rect 84 15577 96 15611
rect -96 15571 96 15577
rect -96 15503 96 15509
rect -96 15469 -84 15503
rect 84 15469 96 15503
rect -96 15463 96 15469
rect -152 15410 -106 15422
rect -152 14634 -146 15410
rect -112 14634 -106 15410
rect -152 14622 -106 14634
rect 106 15410 152 15422
rect 106 14634 112 15410
rect 146 14634 152 15410
rect 106 14622 152 14634
rect -96 14575 96 14581
rect -96 14541 -84 14575
rect 84 14541 96 14575
rect -96 14535 96 14541
rect -96 14467 96 14473
rect -96 14433 -84 14467
rect 84 14433 96 14467
rect -96 14427 96 14433
rect -152 14374 -106 14386
rect -152 13598 -146 14374
rect -112 13598 -106 14374
rect -152 13586 -106 13598
rect 106 14374 152 14386
rect 106 13598 112 14374
rect 146 13598 152 14374
rect 106 13586 152 13598
rect -96 13539 96 13545
rect -96 13505 -84 13539
rect 84 13505 96 13539
rect -96 13499 96 13505
rect -96 13431 96 13437
rect -96 13397 -84 13431
rect 84 13397 96 13431
rect -96 13391 96 13397
rect -152 13338 -106 13350
rect -152 12562 -146 13338
rect -112 12562 -106 13338
rect -152 12550 -106 12562
rect 106 13338 152 13350
rect 106 12562 112 13338
rect 146 12562 152 13338
rect 106 12550 152 12562
rect -96 12503 96 12509
rect -96 12469 -84 12503
rect 84 12469 96 12503
rect -96 12463 96 12469
rect -96 12395 96 12401
rect -96 12361 -84 12395
rect 84 12361 96 12395
rect -96 12355 96 12361
rect -152 12302 -106 12314
rect -152 11526 -146 12302
rect -112 11526 -106 12302
rect -152 11514 -106 11526
rect 106 12302 152 12314
rect 106 11526 112 12302
rect 146 11526 152 12302
rect 106 11514 152 11526
rect -96 11467 96 11473
rect -96 11433 -84 11467
rect 84 11433 96 11467
rect -96 11427 96 11433
rect -96 11359 96 11365
rect -96 11325 -84 11359
rect 84 11325 96 11359
rect -96 11319 96 11325
rect -152 11266 -106 11278
rect -152 10490 -146 11266
rect -112 10490 -106 11266
rect -152 10478 -106 10490
rect 106 11266 152 11278
rect 106 10490 112 11266
rect 146 10490 152 11266
rect 106 10478 152 10490
rect -96 10431 96 10437
rect -96 10397 -84 10431
rect 84 10397 96 10431
rect -96 10391 96 10397
rect -96 10323 96 10329
rect -96 10289 -84 10323
rect 84 10289 96 10323
rect -96 10283 96 10289
rect -152 10230 -106 10242
rect -152 9454 -146 10230
rect -112 9454 -106 10230
rect -152 9442 -106 9454
rect 106 10230 152 10242
rect 106 9454 112 10230
rect 146 9454 152 10230
rect 106 9442 152 9454
rect -96 9395 96 9401
rect -96 9361 -84 9395
rect 84 9361 96 9395
rect -96 9355 96 9361
rect -96 9287 96 9293
rect -96 9253 -84 9287
rect 84 9253 96 9287
rect -96 9247 96 9253
rect -152 9194 -106 9206
rect -152 8418 -146 9194
rect -112 8418 -106 9194
rect -152 8406 -106 8418
rect 106 9194 152 9206
rect 106 8418 112 9194
rect 146 8418 152 9194
rect 106 8406 152 8418
rect -96 8359 96 8365
rect -96 8325 -84 8359
rect 84 8325 96 8359
rect -96 8319 96 8325
rect -96 8251 96 8257
rect -96 8217 -84 8251
rect 84 8217 96 8251
rect -96 8211 96 8217
rect -152 8158 -106 8170
rect -152 7382 -146 8158
rect -112 7382 -106 8158
rect -152 7370 -106 7382
rect 106 8158 152 8170
rect 106 7382 112 8158
rect 146 7382 152 8158
rect 106 7370 152 7382
rect -96 7323 96 7329
rect -96 7289 -84 7323
rect 84 7289 96 7323
rect -96 7283 96 7289
rect -96 7215 96 7221
rect -96 7181 -84 7215
rect 84 7181 96 7215
rect -96 7175 96 7181
rect -152 7122 -106 7134
rect -152 6346 -146 7122
rect -112 6346 -106 7122
rect -152 6334 -106 6346
rect 106 7122 152 7134
rect 106 6346 112 7122
rect 146 6346 152 7122
rect 106 6334 152 6346
rect -96 6287 96 6293
rect -96 6253 -84 6287
rect 84 6253 96 6287
rect -96 6247 96 6253
rect -96 6179 96 6185
rect -96 6145 -84 6179
rect 84 6145 96 6179
rect -96 6139 96 6145
rect -152 6086 -106 6098
rect -152 5310 -146 6086
rect -112 5310 -106 6086
rect -152 5298 -106 5310
rect 106 6086 152 6098
rect 106 5310 112 6086
rect 146 5310 152 6086
rect 106 5298 152 5310
rect -96 5251 96 5257
rect -96 5217 -84 5251
rect 84 5217 96 5251
rect -96 5211 96 5217
rect -96 5143 96 5149
rect -96 5109 -84 5143
rect 84 5109 96 5143
rect -96 5103 96 5109
rect -152 5050 -106 5062
rect -152 4274 -146 5050
rect -112 4274 -106 5050
rect -152 4262 -106 4274
rect 106 5050 152 5062
rect 106 4274 112 5050
rect 146 4274 152 5050
rect 106 4262 152 4274
rect -96 4215 96 4221
rect -96 4181 -84 4215
rect 84 4181 96 4215
rect -96 4175 96 4181
rect -96 4107 96 4113
rect -96 4073 -84 4107
rect 84 4073 96 4107
rect -96 4067 96 4073
rect -152 4014 -106 4026
rect -152 3238 -146 4014
rect -112 3238 -106 4014
rect -152 3226 -106 3238
rect 106 4014 152 4026
rect 106 3238 112 4014
rect 146 3238 152 4014
rect 106 3226 152 3238
rect -96 3179 96 3185
rect -96 3145 -84 3179
rect 84 3145 96 3179
rect -96 3139 96 3145
rect -96 3071 96 3077
rect -96 3037 -84 3071
rect 84 3037 96 3071
rect -96 3031 96 3037
rect -152 2978 -106 2990
rect -152 2202 -146 2978
rect -112 2202 -106 2978
rect -152 2190 -106 2202
rect 106 2978 152 2990
rect 106 2202 112 2978
rect 146 2202 152 2978
rect 106 2190 152 2202
rect -96 2143 96 2149
rect -96 2109 -84 2143
rect 84 2109 96 2143
rect -96 2103 96 2109
rect -96 2035 96 2041
rect -96 2001 -84 2035
rect 84 2001 96 2035
rect -96 1995 96 2001
rect -152 1942 -106 1954
rect -152 1166 -146 1942
rect -112 1166 -106 1942
rect -152 1154 -106 1166
rect 106 1942 152 1954
rect 106 1166 112 1942
rect 146 1166 152 1942
rect 106 1154 152 1166
rect -96 1107 96 1113
rect -96 1073 -84 1107
rect 84 1073 96 1107
rect -96 1067 96 1073
rect -96 999 96 1005
rect -96 965 -84 999
rect 84 965 96 999
rect -96 959 96 965
rect -152 906 -106 918
rect -152 130 -146 906
rect -112 130 -106 906
rect -152 118 -106 130
rect 106 906 152 918
rect 106 130 112 906
rect 146 130 152 906
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -906 -146 -130
rect -112 -906 -106 -130
rect -152 -918 -106 -906
rect 106 -130 152 -118
rect 106 -906 112 -130
rect 146 -906 152 -130
rect 106 -918 152 -906
rect -96 -965 96 -959
rect -96 -999 -84 -965
rect 84 -999 96 -965
rect -96 -1005 96 -999
rect -96 -1073 96 -1067
rect -96 -1107 -84 -1073
rect 84 -1107 96 -1073
rect -96 -1113 96 -1107
rect -152 -1166 -106 -1154
rect -152 -1942 -146 -1166
rect -112 -1942 -106 -1166
rect -152 -1954 -106 -1942
rect 106 -1166 152 -1154
rect 106 -1942 112 -1166
rect 146 -1942 152 -1166
rect 106 -1954 152 -1942
rect -96 -2001 96 -1995
rect -96 -2035 -84 -2001
rect 84 -2035 96 -2001
rect -96 -2041 96 -2035
rect -96 -2109 96 -2103
rect -96 -2143 -84 -2109
rect 84 -2143 96 -2109
rect -96 -2149 96 -2143
rect -152 -2202 -106 -2190
rect -152 -2978 -146 -2202
rect -112 -2978 -106 -2202
rect -152 -2990 -106 -2978
rect 106 -2202 152 -2190
rect 106 -2978 112 -2202
rect 146 -2978 152 -2202
rect 106 -2990 152 -2978
rect -96 -3037 96 -3031
rect -96 -3071 -84 -3037
rect 84 -3071 96 -3037
rect -96 -3077 96 -3071
rect -96 -3145 96 -3139
rect -96 -3179 -84 -3145
rect 84 -3179 96 -3145
rect -96 -3185 96 -3179
rect -152 -3238 -106 -3226
rect -152 -4014 -146 -3238
rect -112 -4014 -106 -3238
rect -152 -4026 -106 -4014
rect 106 -3238 152 -3226
rect 106 -4014 112 -3238
rect 146 -4014 152 -3238
rect 106 -4026 152 -4014
rect -96 -4073 96 -4067
rect -96 -4107 -84 -4073
rect 84 -4107 96 -4073
rect -96 -4113 96 -4107
rect -96 -4181 96 -4175
rect -96 -4215 -84 -4181
rect 84 -4215 96 -4181
rect -96 -4221 96 -4215
rect -152 -4274 -106 -4262
rect -152 -5050 -146 -4274
rect -112 -5050 -106 -4274
rect -152 -5062 -106 -5050
rect 106 -4274 152 -4262
rect 106 -5050 112 -4274
rect 146 -5050 152 -4274
rect 106 -5062 152 -5050
rect -96 -5109 96 -5103
rect -96 -5143 -84 -5109
rect 84 -5143 96 -5109
rect -96 -5149 96 -5143
rect -96 -5217 96 -5211
rect -96 -5251 -84 -5217
rect 84 -5251 96 -5217
rect -96 -5257 96 -5251
rect -152 -5310 -106 -5298
rect -152 -6086 -146 -5310
rect -112 -6086 -106 -5310
rect -152 -6098 -106 -6086
rect 106 -5310 152 -5298
rect 106 -6086 112 -5310
rect 146 -6086 152 -5310
rect 106 -6098 152 -6086
rect -96 -6145 96 -6139
rect -96 -6179 -84 -6145
rect 84 -6179 96 -6145
rect -96 -6185 96 -6179
rect -96 -6253 96 -6247
rect -96 -6287 -84 -6253
rect 84 -6287 96 -6253
rect -96 -6293 96 -6287
rect -152 -6346 -106 -6334
rect -152 -7122 -146 -6346
rect -112 -7122 -106 -6346
rect -152 -7134 -106 -7122
rect 106 -6346 152 -6334
rect 106 -7122 112 -6346
rect 146 -7122 152 -6346
rect 106 -7134 152 -7122
rect -96 -7181 96 -7175
rect -96 -7215 -84 -7181
rect 84 -7215 96 -7181
rect -96 -7221 96 -7215
rect -96 -7289 96 -7283
rect -96 -7323 -84 -7289
rect 84 -7323 96 -7289
rect -96 -7329 96 -7323
rect -152 -7382 -106 -7370
rect -152 -8158 -146 -7382
rect -112 -8158 -106 -7382
rect -152 -8170 -106 -8158
rect 106 -7382 152 -7370
rect 106 -8158 112 -7382
rect 146 -8158 152 -7382
rect 106 -8170 152 -8158
rect -96 -8217 96 -8211
rect -96 -8251 -84 -8217
rect 84 -8251 96 -8217
rect -96 -8257 96 -8251
rect -96 -8325 96 -8319
rect -96 -8359 -84 -8325
rect 84 -8359 96 -8325
rect -96 -8365 96 -8359
rect -152 -8418 -106 -8406
rect -152 -9194 -146 -8418
rect -112 -9194 -106 -8418
rect -152 -9206 -106 -9194
rect 106 -8418 152 -8406
rect 106 -9194 112 -8418
rect 146 -9194 152 -8418
rect 106 -9206 152 -9194
rect -96 -9253 96 -9247
rect -96 -9287 -84 -9253
rect 84 -9287 96 -9253
rect -96 -9293 96 -9287
rect -96 -9361 96 -9355
rect -96 -9395 -84 -9361
rect 84 -9395 96 -9361
rect -96 -9401 96 -9395
rect -152 -9454 -106 -9442
rect -152 -10230 -146 -9454
rect -112 -10230 -106 -9454
rect -152 -10242 -106 -10230
rect 106 -9454 152 -9442
rect 106 -10230 112 -9454
rect 146 -10230 152 -9454
rect 106 -10242 152 -10230
rect -96 -10289 96 -10283
rect -96 -10323 -84 -10289
rect 84 -10323 96 -10289
rect -96 -10329 96 -10323
rect -96 -10397 96 -10391
rect -96 -10431 -84 -10397
rect 84 -10431 96 -10397
rect -96 -10437 96 -10431
rect -152 -10490 -106 -10478
rect -152 -11266 -146 -10490
rect -112 -11266 -106 -10490
rect -152 -11278 -106 -11266
rect 106 -10490 152 -10478
rect 106 -11266 112 -10490
rect 146 -11266 152 -10490
rect 106 -11278 152 -11266
rect -96 -11325 96 -11319
rect -96 -11359 -84 -11325
rect 84 -11359 96 -11325
rect -96 -11365 96 -11359
rect -96 -11433 96 -11427
rect -96 -11467 -84 -11433
rect 84 -11467 96 -11433
rect -96 -11473 96 -11467
rect -152 -11526 -106 -11514
rect -152 -12302 -146 -11526
rect -112 -12302 -106 -11526
rect -152 -12314 -106 -12302
rect 106 -11526 152 -11514
rect 106 -12302 112 -11526
rect 146 -12302 152 -11526
rect 106 -12314 152 -12302
rect -96 -12361 96 -12355
rect -96 -12395 -84 -12361
rect 84 -12395 96 -12361
rect -96 -12401 96 -12395
rect -96 -12469 96 -12463
rect -96 -12503 -84 -12469
rect 84 -12503 96 -12469
rect -96 -12509 96 -12503
rect -152 -12562 -106 -12550
rect -152 -13338 -146 -12562
rect -112 -13338 -106 -12562
rect -152 -13350 -106 -13338
rect 106 -12562 152 -12550
rect 106 -13338 112 -12562
rect 146 -13338 152 -12562
rect 106 -13350 152 -13338
rect -96 -13397 96 -13391
rect -96 -13431 -84 -13397
rect 84 -13431 96 -13397
rect -96 -13437 96 -13431
rect -96 -13505 96 -13499
rect -96 -13539 -84 -13505
rect 84 -13539 96 -13505
rect -96 -13545 96 -13539
rect -152 -13598 -106 -13586
rect -152 -14374 -146 -13598
rect -112 -14374 -106 -13598
rect -152 -14386 -106 -14374
rect 106 -13598 152 -13586
rect 106 -14374 112 -13598
rect 146 -14374 152 -13598
rect 106 -14386 152 -14374
rect -96 -14433 96 -14427
rect -96 -14467 -84 -14433
rect 84 -14467 96 -14433
rect -96 -14473 96 -14467
rect -96 -14541 96 -14535
rect -96 -14575 -84 -14541
rect 84 -14575 96 -14541
rect -96 -14581 96 -14575
rect -152 -14634 -106 -14622
rect -152 -15410 -146 -14634
rect -112 -15410 -106 -14634
rect -152 -15422 -106 -15410
rect 106 -14634 152 -14622
rect 106 -15410 112 -14634
rect 146 -15410 152 -14634
rect 106 -15422 152 -15410
rect -96 -15469 96 -15463
rect -96 -15503 -84 -15469
rect 84 -15503 96 -15469
rect -96 -15509 96 -15503
rect -96 -15577 96 -15571
rect -96 -15611 -84 -15577
rect 84 -15611 96 -15577
rect -96 -15617 96 -15611
rect -152 -15670 -106 -15658
rect -152 -16446 -146 -15670
rect -112 -16446 -106 -15670
rect -152 -16458 -106 -16446
rect 106 -15670 152 -15658
rect 106 -16446 112 -15670
rect 146 -16446 152 -15670
rect 106 -16458 152 -16446
rect -96 -16505 96 -16499
rect -96 -16539 -84 -16505
rect 84 -16539 96 -16505
rect -96 -16545 96 -16539
rect -96 -16613 96 -16607
rect -96 -16647 -84 -16613
rect 84 -16647 96 -16613
rect -96 -16653 96 -16647
rect -152 -16706 -106 -16694
rect -152 -17482 -146 -16706
rect -112 -17482 -106 -16706
rect -152 -17494 -106 -17482
rect 106 -16706 152 -16694
rect 106 -17482 112 -16706
rect 146 -17482 152 -16706
rect 106 -17494 152 -17482
rect -96 -17541 96 -17535
rect -96 -17575 -84 -17541
rect 84 -17575 96 -17541
rect -96 -17581 96 -17575
rect -96 -17649 96 -17643
rect -96 -17683 -84 -17649
rect 84 -17683 96 -17649
rect -96 -17689 96 -17683
rect -152 -17742 -106 -17730
rect -152 -18518 -146 -17742
rect -112 -18518 -106 -17742
rect -152 -18530 -106 -18518
rect 106 -17742 152 -17730
rect 106 -18518 112 -17742
rect 146 -18518 152 -17742
rect 106 -18530 152 -18518
rect -96 -18577 96 -18571
rect -96 -18611 -84 -18577
rect 84 -18611 96 -18577
rect -96 -18617 96 -18611
rect -96 -18685 96 -18679
rect -96 -18719 -84 -18685
rect 84 -18719 96 -18685
rect -96 -18725 96 -18719
rect -152 -18778 -106 -18766
rect -152 -19554 -146 -18778
rect -112 -19554 -106 -18778
rect -152 -19566 -106 -19554
rect 106 -18778 152 -18766
rect 106 -19554 112 -18778
rect 146 -19554 152 -18778
rect 106 -19566 152 -19554
rect -96 -19613 96 -19607
rect -96 -19647 -84 -19613
rect 84 -19647 96 -19613
rect -96 -19653 96 -19647
rect -96 -19721 96 -19715
rect -96 -19755 -84 -19721
rect 84 -19755 96 -19721
rect -96 -19761 96 -19755
rect -152 -19814 -106 -19802
rect -152 -20590 -146 -19814
rect -112 -20590 -106 -19814
rect -152 -20602 -106 -20590
rect 106 -19814 152 -19802
rect 106 -20590 112 -19814
rect 146 -20590 152 -19814
rect 106 -20602 152 -20590
rect -96 -20649 96 -20643
rect -96 -20683 -84 -20649
rect 84 -20683 96 -20649
rect -96 -20689 96 -20683
rect -96 -20757 96 -20751
rect -96 -20791 -84 -20757
rect 84 -20791 96 -20757
rect -96 -20797 96 -20791
rect -152 -20850 -106 -20838
rect -152 -21626 -146 -20850
rect -112 -21626 -106 -20850
rect -152 -21638 -106 -21626
rect 106 -20850 152 -20838
rect 106 -21626 112 -20850
rect 146 -21626 152 -20850
rect 106 -21638 152 -21626
rect -96 -21685 96 -21679
rect -96 -21719 -84 -21685
rect 84 -21719 96 -21685
rect -96 -21725 96 -21719
rect -96 -21793 96 -21787
rect -96 -21827 -84 -21793
rect 84 -21827 96 -21793
rect -96 -21833 96 -21827
rect -152 -21886 -106 -21874
rect -152 -22662 -146 -21886
rect -112 -22662 -106 -21886
rect -152 -22674 -106 -22662
rect 106 -21886 152 -21874
rect 106 -22662 112 -21886
rect 146 -22662 152 -21886
rect 106 -22674 152 -22662
rect -96 -22721 96 -22715
rect -96 -22755 -84 -22721
rect 84 -22755 96 -22721
rect -96 -22761 96 -22755
rect -96 -22829 96 -22823
rect -96 -22863 -84 -22829
rect 84 -22863 96 -22829
rect -96 -22869 96 -22863
rect -152 -22922 -106 -22910
rect -152 -23698 -146 -22922
rect -112 -23698 -106 -22922
rect -152 -23710 -106 -23698
rect 106 -22922 152 -22910
rect 106 -23698 112 -22922
rect 146 -23698 152 -22922
rect 106 -23710 152 -23698
rect -96 -23757 96 -23751
rect -96 -23791 -84 -23757
rect 84 -23791 96 -23757
rect -96 -23797 96 -23791
rect -96 -23865 96 -23859
rect -96 -23899 -84 -23865
rect 84 -23899 96 -23865
rect -96 -23905 96 -23899
rect -152 -23958 -106 -23946
rect -152 -24734 -146 -23958
rect -112 -24734 -106 -23958
rect -152 -24746 -106 -24734
rect 106 -23958 152 -23946
rect 106 -24734 112 -23958
rect 146 -24734 152 -23958
rect 106 -24746 152 -24734
rect -96 -24793 96 -24787
rect -96 -24827 -84 -24793
rect 84 -24827 96 -24793
rect -96 -24833 96 -24827
rect -96 -24901 96 -24895
rect -96 -24935 -84 -24901
rect 84 -24935 96 -24901
rect -96 -24941 96 -24935
rect -152 -24994 -106 -24982
rect -152 -25770 -146 -24994
rect -112 -25770 -106 -24994
rect -152 -25782 -106 -25770
rect 106 -24994 152 -24982
rect 106 -25770 112 -24994
rect 146 -25770 152 -24994
rect 106 -25782 152 -25770
rect -96 -25829 96 -25823
rect -96 -25863 -84 -25829
rect 84 -25863 96 -25829
rect -96 -25869 96 -25863
rect -96 -25937 96 -25931
rect -96 -25971 -84 -25937
rect 84 -25971 96 -25937
rect -96 -25977 96 -25971
rect -152 -26030 -106 -26018
rect -152 -26806 -146 -26030
rect -112 -26806 -106 -26030
rect -152 -26818 -106 -26806
rect 106 -26030 152 -26018
rect 106 -26806 112 -26030
rect 146 -26806 152 -26030
rect 106 -26818 152 -26806
rect -96 -26865 96 -26859
rect -96 -26899 -84 -26865
rect 84 -26899 96 -26865
rect -96 -26905 96 -26899
rect -96 -26973 96 -26967
rect -96 -27007 -84 -26973
rect 84 -27007 96 -26973
rect -96 -27013 96 -27007
rect -152 -27066 -106 -27054
rect -152 -27842 -146 -27066
rect -112 -27842 -106 -27066
rect -152 -27854 -106 -27842
rect 106 -27066 152 -27054
rect 106 -27842 112 -27066
rect 146 -27842 152 -27066
rect 106 -27854 152 -27842
rect -96 -27901 96 -27895
rect -96 -27935 -84 -27901
rect 84 -27935 96 -27901
rect -96 -27941 96 -27935
rect -96 -28009 96 -28003
rect -96 -28043 -84 -28009
rect 84 -28043 96 -28009
rect -96 -28049 96 -28043
rect -152 -28102 -106 -28090
rect -152 -28878 -146 -28102
rect -112 -28878 -106 -28102
rect -152 -28890 -106 -28878
rect 106 -28102 152 -28090
rect 106 -28878 112 -28102
rect 146 -28878 152 -28102
rect 106 -28890 152 -28878
rect -96 -28937 96 -28931
rect -96 -28971 -84 -28937
rect 84 -28971 96 -28937
rect -96 -28977 96 -28971
rect -96 -29045 96 -29039
rect -96 -29079 -84 -29045
rect 84 -29079 96 -29045
rect -96 -29085 96 -29079
rect -152 -29138 -106 -29126
rect -152 -29914 -146 -29138
rect -112 -29914 -106 -29138
rect -152 -29926 -106 -29914
rect 106 -29138 152 -29126
rect 106 -29914 112 -29138
rect 146 -29914 152 -29138
rect 106 -29926 152 -29914
rect -96 -29973 96 -29967
rect -96 -30007 -84 -29973
rect 84 -30007 96 -29973
rect -96 -30013 96 -30007
rect -96 -30081 96 -30075
rect -96 -30115 -84 -30081
rect 84 -30115 96 -30081
rect -96 -30121 96 -30115
rect -152 -30174 -106 -30162
rect -152 -30950 -146 -30174
rect -112 -30950 -106 -30174
rect -152 -30962 -106 -30950
rect 106 -30174 152 -30162
rect 106 -30950 112 -30174
rect 146 -30950 152 -30174
rect 106 -30962 152 -30950
rect -96 -31009 96 -31003
rect -96 -31043 -84 -31009
rect 84 -31043 96 -31009
rect -96 -31049 96 -31043
rect -96 -31117 96 -31111
rect -96 -31151 -84 -31117
rect 84 -31151 96 -31117
rect -96 -31157 96 -31151
rect -152 -31210 -106 -31198
rect -152 -31986 -146 -31210
rect -112 -31986 -106 -31210
rect -152 -31998 -106 -31986
rect 106 -31210 152 -31198
rect 106 -31986 112 -31210
rect 146 -31986 152 -31210
rect 106 -31998 152 -31986
rect -96 -32045 96 -32039
rect -96 -32079 -84 -32045
rect 84 -32079 96 -32045
rect -96 -32085 96 -32079
rect -96 -32153 96 -32147
rect -96 -32187 -84 -32153
rect 84 -32187 96 -32153
rect -96 -32193 96 -32187
rect -152 -32246 -106 -32234
rect -152 -33022 -146 -32246
rect -112 -33022 -106 -32246
rect -152 -33034 -106 -33022
rect 106 -32246 152 -32234
rect 106 -33022 112 -32246
rect 146 -33022 152 -32246
rect 106 -33034 152 -33022
rect -96 -33081 96 -33075
rect -96 -33115 -84 -33081
rect 84 -33115 96 -33081
rect -96 -33121 96 -33115
rect -96 -33189 96 -33183
rect -96 -33223 -84 -33189
rect 84 -33223 96 -33189
rect -96 -33229 96 -33223
rect -152 -33282 -106 -33270
rect -152 -34058 -146 -33282
rect -112 -34058 -106 -33282
rect -152 -34070 -106 -34058
rect 106 -33282 152 -33270
rect 106 -34058 112 -33282
rect 146 -34058 152 -33282
rect 106 -34070 152 -34058
rect -96 -34117 96 -34111
rect -96 -34151 -84 -34117
rect 84 -34151 96 -34117
rect -96 -34157 96 -34151
rect -96 -34225 96 -34219
rect -96 -34259 -84 -34225
rect 84 -34259 96 -34225
rect -96 -34265 96 -34259
rect -152 -34318 -106 -34306
rect -152 -35094 -146 -34318
rect -112 -35094 -106 -34318
rect -152 -35106 -106 -35094
rect 106 -34318 152 -34306
rect 106 -35094 112 -34318
rect 146 -35094 152 -34318
rect 106 -35106 152 -35094
rect -96 -35153 96 -35147
rect -96 -35187 -84 -35153
rect 84 -35187 96 -35153
rect -96 -35193 96 -35187
rect -96 -35261 96 -35255
rect -96 -35295 -84 -35261
rect 84 -35295 96 -35261
rect -96 -35301 96 -35295
rect -152 -35354 -106 -35342
rect -152 -36130 -146 -35354
rect -112 -36130 -106 -35354
rect -152 -36142 -106 -36130
rect 106 -35354 152 -35342
rect 106 -36130 112 -35354
rect 146 -36130 152 -35354
rect 106 -36142 152 -36130
rect -96 -36189 96 -36183
rect -96 -36223 -84 -36189
rect 84 -36223 96 -36189
rect -96 -36229 96 -36223
rect -96 -36297 96 -36291
rect -96 -36331 -84 -36297
rect 84 -36331 96 -36297
rect -96 -36337 96 -36331
rect -152 -36390 -106 -36378
rect -152 -37166 -146 -36390
rect -112 -37166 -106 -36390
rect -152 -37178 -106 -37166
rect 106 -36390 152 -36378
rect 106 -37166 112 -36390
rect 146 -37166 152 -36390
rect 106 -37178 152 -37166
rect -96 -37225 96 -37219
rect -96 -37259 -84 -37225
rect 84 -37259 96 -37225
rect -96 -37265 96 -37259
rect -96 -37333 96 -37327
rect -96 -37367 -84 -37333
rect 84 -37367 96 -37333
rect -96 -37373 96 -37367
rect -152 -37426 -106 -37414
rect -152 -38202 -146 -37426
rect -112 -38202 -106 -37426
rect -152 -38214 -106 -38202
rect 106 -37426 152 -37414
rect 106 -38202 112 -37426
rect 146 -38202 152 -37426
rect 106 -38214 152 -38202
rect -96 -38261 96 -38255
rect -96 -38295 -84 -38261
rect 84 -38295 96 -38261
rect -96 -38301 96 -38295
rect -96 -38369 96 -38363
rect -96 -38403 -84 -38369
rect 84 -38403 96 -38369
rect -96 -38409 96 -38403
rect -152 -38462 -106 -38450
rect -152 -39238 -146 -38462
rect -112 -39238 -106 -38462
rect -152 -39250 -106 -39238
rect 106 -38462 152 -38450
rect 106 -39238 112 -38462
rect 146 -39238 152 -38462
rect 106 -39250 152 -39238
rect -96 -39297 96 -39291
rect -96 -39331 -84 -39297
rect 84 -39331 96 -39297
rect -96 -39337 96 -39331
rect -96 -39405 96 -39399
rect -96 -39439 -84 -39405
rect 84 -39439 96 -39405
rect -96 -39445 96 -39439
rect -152 -39498 -106 -39486
rect -152 -40274 -146 -39498
rect -112 -40274 -106 -39498
rect -152 -40286 -106 -40274
rect 106 -39498 152 -39486
rect 106 -40274 112 -39498
rect 146 -40274 152 -39498
rect 106 -40286 152 -40274
rect -96 -40333 96 -40327
rect -96 -40367 -84 -40333
rect 84 -40367 96 -40333
rect -96 -40373 96 -40367
rect -96 -40441 96 -40435
rect -96 -40475 -84 -40441
rect 84 -40475 96 -40441
rect -96 -40481 96 -40475
rect -152 -40534 -106 -40522
rect -152 -41310 -146 -40534
rect -112 -41310 -106 -40534
rect -152 -41322 -106 -41310
rect 106 -40534 152 -40522
rect 106 -41310 112 -40534
rect 146 -41310 152 -40534
rect 106 -41322 152 -41310
rect -96 -41369 96 -41363
rect -96 -41403 -84 -41369
rect 84 -41403 96 -41369
rect -96 -41409 96 -41403
rect -96 -41477 96 -41471
rect -96 -41511 -84 -41477
rect 84 -41511 96 -41477
rect -96 -41517 96 -41511
rect -152 -41570 -106 -41558
rect -152 -42346 -146 -41570
rect -112 -42346 -106 -41570
rect -152 -42358 -106 -42346
rect 106 -41570 152 -41558
rect 106 -42346 112 -41570
rect 146 -42346 152 -41570
rect 106 -42358 152 -42346
rect -96 -42405 96 -42399
rect -96 -42439 -84 -42405
rect 84 -42439 96 -42405
rect -96 -42445 96 -42439
rect -96 -42513 96 -42507
rect -96 -42547 -84 -42513
rect 84 -42547 96 -42513
rect -96 -42553 96 -42547
rect -152 -42606 -106 -42594
rect -152 -43382 -146 -42606
rect -112 -43382 -106 -42606
rect -152 -43394 -106 -43382
rect 106 -42606 152 -42594
rect 106 -43382 112 -42606
rect 146 -43382 152 -42606
rect 106 -43394 152 -43382
rect -96 -43441 96 -43435
rect -96 -43475 -84 -43441
rect 84 -43475 96 -43441
rect -96 -43481 96 -43475
rect -96 -43549 96 -43543
rect -96 -43583 -84 -43549
rect 84 -43583 96 -43549
rect -96 -43589 96 -43583
rect -152 -43642 -106 -43630
rect -152 -44418 -146 -43642
rect -112 -44418 -106 -43642
rect -152 -44430 -106 -44418
rect 106 -43642 152 -43630
rect 106 -44418 112 -43642
rect 146 -44418 152 -43642
rect 106 -44430 152 -44418
rect -96 -44477 96 -44471
rect -96 -44511 -84 -44477
rect 84 -44511 96 -44477
rect -96 -44517 96 -44511
rect -96 -44585 96 -44579
rect -96 -44619 -84 -44585
rect 84 -44619 96 -44585
rect -96 -44625 96 -44619
rect -152 -44678 -106 -44666
rect -152 -45454 -146 -44678
rect -112 -45454 -106 -44678
rect -152 -45466 -106 -45454
rect 106 -44678 152 -44666
rect 106 -45454 112 -44678
rect 146 -45454 152 -44678
rect 106 -45466 152 -45454
rect -96 -45513 96 -45507
rect -96 -45547 -84 -45513
rect 84 -45547 96 -45513
rect -96 -45553 96 -45547
rect -96 -45621 96 -45615
rect -96 -45655 -84 -45621
rect 84 -45655 96 -45621
rect -96 -45661 96 -45655
rect -152 -45714 -106 -45702
rect -152 -46490 -146 -45714
rect -112 -46490 -106 -45714
rect -152 -46502 -106 -46490
rect 106 -45714 152 -45702
rect 106 -46490 112 -45714
rect 146 -46490 152 -45714
rect 106 -46502 152 -46490
rect -96 -46549 96 -46543
rect -96 -46583 -84 -46549
rect 84 -46583 96 -46549
rect -96 -46589 96 -46583
rect -96 -46657 96 -46651
rect -96 -46691 -84 -46657
rect 84 -46691 96 -46657
rect -96 -46697 96 -46691
rect -152 -46750 -106 -46738
rect -152 -47526 -146 -46750
rect -112 -47526 -106 -46750
rect -152 -47538 -106 -47526
rect 106 -46750 152 -46738
rect 106 -47526 112 -46750
rect 146 -47526 152 -46750
rect 106 -47538 152 -47526
rect -96 -47585 96 -47579
rect -96 -47619 -84 -47585
rect 84 -47619 96 -47585
rect -96 -47625 96 -47619
rect -96 -47693 96 -47687
rect -96 -47727 -84 -47693
rect 84 -47727 96 -47693
rect -96 -47733 96 -47727
rect -152 -47786 -106 -47774
rect -152 -48562 -146 -47786
rect -112 -48562 -106 -47786
rect -152 -48574 -106 -48562
rect 106 -47786 152 -47774
rect 106 -48562 112 -47786
rect 146 -48562 152 -47786
rect 106 -48574 152 -48562
rect -96 -48621 96 -48615
rect -96 -48655 -84 -48621
rect 84 -48655 96 -48621
rect -96 -48661 96 -48655
rect -96 -48729 96 -48723
rect -96 -48763 -84 -48729
rect 84 -48763 96 -48729
rect -96 -48769 96 -48763
rect -152 -48822 -106 -48810
rect -152 -49598 -146 -48822
rect -112 -49598 -106 -48822
rect -152 -49610 -106 -49598
rect 106 -48822 152 -48810
rect 106 -49598 112 -48822
rect 146 -49598 152 -48822
rect 106 -49610 152 -49598
rect -96 -49657 96 -49651
rect -96 -49691 -84 -49657
rect 84 -49691 96 -49657
rect -96 -49697 96 -49691
rect -96 -49765 96 -49759
rect -96 -49799 -84 -49765
rect 84 -49799 96 -49765
rect -96 -49805 96 -49799
rect -152 -49858 -106 -49846
rect -152 -50634 -146 -49858
rect -112 -50634 -106 -49858
rect -152 -50646 -106 -50634
rect 106 -49858 152 -49846
rect 106 -50634 112 -49858
rect 146 -50634 152 -49858
rect 106 -50646 152 -50634
rect -96 -50693 96 -50687
rect -96 -50727 -84 -50693
rect 84 -50727 96 -50693
rect -96 -50733 96 -50727
rect -96 -50801 96 -50795
rect -96 -50835 -84 -50801
rect 84 -50835 96 -50801
rect -96 -50841 96 -50835
rect -152 -50894 -106 -50882
rect -152 -51670 -146 -50894
rect -112 -51670 -106 -50894
rect -152 -51682 -106 -51670
rect 106 -50894 152 -50882
rect 106 -51670 112 -50894
rect 146 -51670 152 -50894
rect 106 -51682 152 -51670
rect -96 -51729 96 -51723
rect -96 -51763 -84 -51729
rect 84 -51763 96 -51729
rect -96 -51769 96 -51763
rect -96 -51837 96 -51831
rect -96 -51871 -84 -51837
rect 84 -51871 96 -51837
rect -96 -51877 96 -51871
rect -152 -51930 -106 -51918
rect -152 -52706 -146 -51930
rect -112 -52706 -106 -51930
rect -152 -52718 -106 -52706
rect 106 -51930 152 -51918
rect 106 -52706 112 -51930
rect 146 -52706 152 -51930
rect 106 -52718 152 -52706
rect -96 -52765 96 -52759
rect -96 -52799 -84 -52765
rect 84 -52799 96 -52765
rect -96 -52805 96 -52799
rect -96 -52873 96 -52867
rect -96 -52907 -84 -52873
rect 84 -52907 96 -52873
rect -96 -52913 96 -52907
rect -152 -52966 -106 -52954
rect -152 -53742 -146 -52966
rect -112 -53742 -106 -52966
rect -152 -53754 -106 -53742
rect 106 -52966 152 -52954
rect 106 -53742 112 -52966
rect 146 -53742 152 -52966
rect 106 -53754 152 -53742
rect -96 -53801 96 -53795
rect -96 -53835 -84 -53801
rect 84 -53835 96 -53801
rect -96 -53841 96 -53835
rect -96 -53909 96 -53903
rect -96 -53943 -84 -53909
rect 84 -53943 96 -53909
rect -96 -53949 96 -53943
rect -152 -54002 -106 -53990
rect -152 -54778 -146 -54002
rect -112 -54778 -106 -54002
rect -152 -54790 -106 -54778
rect 106 -54002 152 -53990
rect 106 -54778 112 -54002
rect 146 -54778 152 -54002
rect 106 -54790 152 -54778
rect -96 -54837 96 -54831
rect -96 -54871 -84 -54837
rect 84 -54871 96 -54837
rect -96 -54877 96 -54871
rect -96 -54945 96 -54939
rect -96 -54979 -84 -54945
rect 84 -54979 96 -54945
rect -96 -54985 96 -54979
rect -152 -55038 -106 -55026
rect -152 -55814 -146 -55038
rect -112 -55814 -106 -55038
rect -152 -55826 -106 -55814
rect 106 -55038 152 -55026
rect 106 -55814 112 -55038
rect 146 -55814 152 -55038
rect 106 -55826 152 -55814
rect -96 -55873 96 -55867
rect -96 -55907 -84 -55873
rect 84 -55907 96 -55873
rect -96 -55913 96 -55907
rect -96 -55981 96 -55975
rect -96 -56015 -84 -55981
rect 84 -56015 96 -55981
rect -96 -56021 96 -56015
rect -152 -56074 -106 -56062
rect -152 -56850 -146 -56074
rect -112 -56850 -106 -56074
rect -152 -56862 -106 -56850
rect 106 -56074 152 -56062
rect 106 -56850 112 -56074
rect 146 -56850 152 -56074
rect 106 -56862 152 -56850
rect -96 -56909 96 -56903
rect -96 -56943 -84 -56909
rect 84 -56943 96 -56909
rect -96 -56949 96 -56943
rect -96 -57017 96 -57011
rect -96 -57051 -84 -57017
rect 84 -57051 96 -57017
rect -96 -57057 96 -57051
rect -152 -57110 -106 -57098
rect -152 -57886 -146 -57110
rect -112 -57886 -106 -57110
rect -152 -57898 -106 -57886
rect 106 -57110 152 -57098
rect 106 -57886 112 -57110
rect 146 -57886 152 -57110
rect 106 -57898 152 -57886
rect -96 -57945 96 -57939
rect -96 -57979 -84 -57945
rect 84 -57979 96 -57945
rect -96 -57985 96 -57979
rect -96 -58053 96 -58047
rect -96 -58087 -84 -58053
rect 84 -58087 96 -58053
rect -96 -58093 96 -58087
rect -152 -58146 -106 -58134
rect -152 -58922 -146 -58146
rect -112 -58922 -106 -58146
rect -152 -58934 -106 -58922
rect 106 -58146 152 -58134
rect 106 -58922 112 -58146
rect 146 -58922 152 -58146
rect 106 -58934 152 -58922
rect -96 -58981 96 -58975
rect -96 -59015 -84 -58981
rect 84 -59015 96 -58981
rect -96 -59021 96 -59015
rect -96 -59089 96 -59083
rect -96 -59123 -84 -59089
rect 84 -59123 96 -59089
rect -96 -59129 96 -59123
rect -152 -59182 -106 -59170
rect -152 -59958 -146 -59182
rect -112 -59958 -106 -59182
rect -152 -59970 -106 -59958
rect 106 -59182 152 -59170
rect 106 -59958 112 -59182
rect 146 -59958 152 -59182
rect 106 -59970 152 -59958
rect -96 -60017 96 -60011
rect -96 -60051 -84 -60017
rect 84 -60051 96 -60017
rect -96 -60057 96 -60051
rect -96 -60125 96 -60119
rect -96 -60159 -84 -60125
rect 84 -60159 96 -60125
rect -96 -60165 96 -60159
rect -152 -60218 -106 -60206
rect -152 -60994 -146 -60218
rect -112 -60994 -106 -60218
rect -152 -61006 -106 -60994
rect 106 -60218 152 -60206
rect 106 -60994 112 -60218
rect 146 -60994 152 -60218
rect 106 -61006 152 -60994
rect -96 -61053 96 -61047
rect -96 -61087 -84 -61053
rect 84 -61087 96 -61053
rect -96 -61093 96 -61087
rect -96 -61161 96 -61155
rect -96 -61195 -84 -61161
rect 84 -61195 96 -61161
rect -96 -61201 96 -61195
rect -152 -61254 -106 -61242
rect -152 -62030 -146 -61254
rect -112 -62030 -106 -61254
rect -152 -62042 -106 -62030
rect 106 -61254 152 -61242
rect 106 -62030 112 -61254
rect 146 -62030 152 -61254
rect 106 -62042 152 -62030
rect -96 -62089 96 -62083
rect -96 -62123 -84 -62089
rect 84 -62123 96 -62089
rect -96 -62129 96 -62123
rect -96 -62197 96 -62191
rect -96 -62231 -84 -62197
rect 84 -62231 96 -62197
rect -96 -62237 96 -62231
rect -152 -62290 -106 -62278
rect -152 -63066 -146 -62290
rect -112 -63066 -106 -62290
rect -152 -63078 -106 -63066
rect 106 -62290 152 -62278
rect 106 -63066 112 -62290
rect 146 -63066 152 -62290
rect 106 -63078 152 -63066
rect -96 -63125 96 -63119
rect -96 -63159 -84 -63125
rect 84 -63159 96 -63125
rect -96 -63165 96 -63159
rect -96 -63233 96 -63227
rect -96 -63267 -84 -63233
rect 84 -63267 96 -63233
rect -96 -63273 96 -63267
rect -152 -63326 -106 -63314
rect -152 -64102 -146 -63326
rect -112 -64102 -106 -63326
rect -152 -64114 -106 -64102
rect 106 -63326 152 -63314
rect 106 -64102 112 -63326
rect 146 -64102 152 -63326
rect 106 -64114 152 -64102
rect -96 -64161 96 -64155
rect -96 -64195 -84 -64161
rect 84 -64195 96 -64161
rect -96 -64201 96 -64195
rect -96 -64269 96 -64263
rect -96 -64303 -84 -64269
rect 84 -64303 96 -64269
rect -96 -64309 96 -64303
rect -152 -64362 -106 -64350
rect -152 -65138 -146 -64362
rect -112 -65138 -106 -64362
rect -152 -65150 -106 -65138
rect 106 -64362 152 -64350
rect 106 -65138 112 -64362
rect 146 -65138 152 -64362
rect 106 -65150 152 -65138
rect -96 -65197 96 -65191
rect -96 -65231 -84 -65197
rect 84 -65231 96 -65197
rect -96 -65237 96 -65231
rect -96 -65305 96 -65299
rect -96 -65339 -84 -65305
rect 84 -65339 96 -65305
rect -96 -65345 96 -65339
rect -152 -65398 -106 -65386
rect -152 -66174 -146 -65398
rect -112 -66174 -106 -65398
rect -152 -66186 -106 -66174
rect 106 -65398 152 -65386
rect 106 -66174 112 -65398
rect 146 -66174 152 -65398
rect 106 -66186 152 -66174
rect -96 -66233 96 -66227
rect -96 -66267 -84 -66233
rect 84 -66267 96 -66233
rect -96 -66273 96 -66267
rect -96 -66341 96 -66335
rect -96 -66375 -84 -66341
rect 84 -66375 96 -66341
rect -96 -66381 96 -66375
rect -152 -66434 -106 -66422
rect -152 -67210 -146 -66434
rect -112 -67210 -106 -66434
rect -152 -67222 -106 -67210
rect 106 -66434 152 -66422
rect 106 -67210 112 -66434
rect 146 -67210 152 -66434
rect 106 -67222 152 -67210
rect -96 -67269 96 -67263
rect -96 -67303 -84 -67269
rect 84 -67303 96 -67269
rect -96 -67309 96 -67303
rect -96 -67377 96 -67371
rect -96 -67411 -84 -67377
rect 84 -67411 96 -67377
rect -96 -67417 96 -67411
rect -152 -67470 -106 -67458
rect -152 -68246 -146 -67470
rect -112 -68246 -106 -67470
rect -152 -68258 -106 -68246
rect 106 -67470 152 -67458
rect 106 -68246 112 -67470
rect 146 -68246 152 -67470
rect 106 -68258 152 -68246
rect -96 -68305 96 -68299
rect -96 -68339 -84 -68305
rect 84 -68339 96 -68305
rect -96 -68345 96 -68339
rect -96 -68413 96 -68407
rect -96 -68447 -84 -68413
rect 84 -68447 96 -68413
rect -96 -68453 96 -68447
rect -152 -68506 -106 -68494
rect -152 -69282 -146 -68506
rect -112 -69282 -106 -68506
rect -152 -69294 -106 -69282
rect 106 -68506 152 -68494
rect 106 -69282 112 -68506
rect 146 -69282 152 -68506
rect 106 -69294 152 -69282
rect -96 -69341 96 -69335
rect -96 -69375 -84 -69341
rect 84 -69375 96 -69341
rect -96 -69381 96 -69375
rect -96 -69449 96 -69443
rect -96 -69483 -84 -69449
rect 84 -69483 96 -69449
rect -96 -69489 96 -69483
rect -152 -69542 -106 -69530
rect -152 -70318 -146 -69542
rect -112 -70318 -106 -69542
rect -152 -70330 -106 -70318
rect 106 -69542 152 -69530
rect 106 -70318 112 -69542
rect 146 -70318 152 -69542
rect 106 -70330 152 -70318
rect -96 -70377 96 -70371
rect -96 -70411 -84 -70377
rect 84 -70411 96 -70377
rect -96 -70417 96 -70411
rect -96 -70485 96 -70479
rect -96 -70519 -84 -70485
rect 84 -70519 96 -70485
rect -96 -70525 96 -70519
rect -152 -70578 -106 -70566
rect -152 -71354 -146 -70578
rect -112 -71354 -106 -70578
rect -152 -71366 -106 -71354
rect 106 -70578 152 -70566
rect 106 -71354 112 -70578
rect 146 -71354 152 -70578
rect 106 -71366 152 -71354
rect -96 -71413 96 -71407
rect -96 -71447 -84 -71413
rect 84 -71447 96 -71413
rect -96 -71453 96 -71447
rect -96 -71521 96 -71515
rect -96 -71555 -84 -71521
rect 84 -71555 96 -71521
rect -96 -71561 96 -71555
rect -152 -71614 -106 -71602
rect -152 -72390 -146 -71614
rect -112 -72390 -106 -71614
rect -152 -72402 -106 -72390
rect 106 -71614 152 -71602
rect 106 -72390 112 -71614
rect 146 -72390 152 -71614
rect 106 -72402 152 -72390
rect -96 -72449 96 -72443
rect -96 -72483 -84 -72449
rect 84 -72483 96 -72449
rect -96 -72489 96 -72483
rect -96 -72557 96 -72551
rect -96 -72591 -84 -72557
rect 84 -72591 96 -72557
rect -96 -72597 96 -72591
rect -152 -72650 -106 -72638
rect -152 -73426 -146 -72650
rect -112 -73426 -106 -72650
rect -152 -73438 -106 -73426
rect 106 -72650 152 -72638
rect 106 -73426 112 -72650
rect 146 -73426 152 -72650
rect 106 -73438 152 -73426
rect -96 -73485 96 -73479
rect -96 -73519 -84 -73485
rect 84 -73519 96 -73485
rect -96 -73525 96 -73519
rect -96 -73593 96 -73587
rect -96 -73627 -84 -73593
rect 84 -73627 96 -73593
rect -96 -73633 96 -73627
rect -152 -73686 -106 -73674
rect -152 -74462 -146 -73686
rect -112 -74462 -106 -73686
rect -152 -74474 -106 -74462
rect 106 -73686 152 -73674
rect 106 -74462 112 -73686
rect 146 -74462 152 -73686
rect 106 -74474 152 -74462
rect -96 -74521 96 -74515
rect -96 -74555 -84 -74521
rect 84 -74555 96 -74521
rect -96 -74561 96 -74555
rect -96 -74629 96 -74623
rect -96 -74663 -84 -74629
rect 84 -74663 96 -74629
rect -96 -74669 96 -74663
rect -152 -74722 -106 -74710
rect -152 -75498 -146 -74722
rect -112 -75498 -106 -74722
rect -152 -75510 -106 -75498
rect 106 -74722 152 -74710
rect 106 -75498 112 -74722
rect 146 -75498 152 -74722
rect 106 -75510 152 -75498
rect -96 -75557 96 -75551
rect -96 -75591 -84 -75557
rect 84 -75591 96 -75557
rect -96 -75597 96 -75591
rect -96 -75665 96 -75659
rect -96 -75699 -84 -75665
rect 84 -75699 96 -75665
rect -96 -75705 96 -75699
rect -152 -75758 -106 -75746
rect -152 -76534 -146 -75758
rect -112 -76534 -106 -75758
rect -152 -76546 -106 -76534
rect 106 -75758 152 -75746
rect 106 -76534 112 -75758
rect 146 -76534 152 -75758
rect 106 -76546 152 -76534
rect -96 -76593 96 -76587
rect -96 -76627 -84 -76593
rect 84 -76627 96 -76593
rect -96 -76633 96 -76627
rect -96 -76701 96 -76695
rect -96 -76735 -84 -76701
rect 84 -76735 96 -76701
rect -96 -76741 96 -76735
rect -152 -76794 -106 -76782
rect -152 -77570 -146 -76794
rect -112 -77570 -106 -76794
rect -152 -77582 -106 -77570
rect 106 -76794 152 -76782
rect 106 -77570 112 -76794
rect 146 -77570 152 -76794
rect 106 -77582 152 -77570
rect -96 -77629 96 -77623
rect -96 -77663 -84 -77629
rect 84 -77663 96 -77629
rect -96 -77669 96 -77663
rect -96 -77737 96 -77731
rect -96 -77771 -84 -77737
rect 84 -77771 96 -77737
rect -96 -77777 96 -77771
rect -152 -77830 -106 -77818
rect -152 -78606 -146 -77830
rect -112 -78606 -106 -77830
rect -152 -78618 -106 -78606
rect 106 -77830 152 -77818
rect 106 -78606 112 -77830
rect 146 -78606 152 -77830
rect 106 -78618 152 -78606
rect -96 -78665 96 -78659
rect -96 -78699 -84 -78665
rect 84 -78699 96 -78665
rect -96 -78705 96 -78699
rect -96 -78773 96 -78767
rect -96 -78807 -84 -78773
rect 84 -78807 96 -78773
rect -96 -78813 96 -78807
rect -152 -78866 -106 -78854
rect -152 -79642 -146 -78866
rect -112 -79642 -106 -78866
rect -152 -79654 -106 -79642
rect 106 -78866 152 -78854
rect 106 -79642 112 -78866
rect 146 -79642 152 -78866
rect 106 -79654 152 -79642
rect -96 -79701 96 -79695
rect -96 -79735 -84 -79701
rect 84 -79735 96 -79701
rect -96 -79741 96 -79735
rect -96 -79809 96 -79803
rect -96 -79843 -84 -79809
rect 84 -79843 96 -79809
rect -96 -79849 96 -79843
rect -152 -79902 -106 -79890
rect -152 -80678 -146 -79902
rect -112 -80678 -106 -79902
rect -152 -80690 -106 -80678
rect 106 -79902 152 -79890
rect 106 -80678 112 -79902
rect 146 -80678 152 -79902
rect 106 -80690 152 -80678
rect -96 -80737 96 -80731
rect -96 -80771 -84 -80737
rect 84 -80771 96 -80737
rect -96 -80777 96 -80771
rect -96 -80845 96 -80839
rect -96 -80879 -84 -80845
rect 84 -80879 96 -80845
rect -96 -80885 96 -80879
rect -152 -80938 -106 -80926
rect -152 -81714 -146 -80938
rect -112 -81714 -106 -80938
rect -152 -81726 -106 -81714
rect 106 -80938 152 -80926
rect 106 -81714 112 -80938
rect 146 -81714 152 -80938
rect 106 -81726 152 -81714
rect -96 -81773 96 -81767
rect -96 -81807 -84 -81773
rect 84 -81807 96 -81773
rect -96 -81813 96 -81807
rect -96 -81881 96 -81875
rect -96 -81915 -84 -81881
rect 84 -81915 96 -81881
rect -96 -81921 96 -81915
rect -152 -81974 -106 -81962
rect -152 -82750 -146 -81974
rect -112 -82750 -106 -81974
rect -152 -82762 -106 -82750
rect 106 -81974 152 -81962
rect 106 -82750 112 -81974
rect 146 -82750 152 -81974
rect 106 -82762 152 -82750
rect -96 -82809 96 -82803
rect -96 -82843 -84 -82809
rect 84 -82843 96 -82809
rect -96 -82849 96 -82843
rect -96 -82917 96 -82911
rect -96 -82951 -84 -82917
rect 84 -82951 96 -82917
rect -96 -82957 96 -82951
rect -152 -83010 -106 -82998
rect -152 -83786 -146 -83010
rect -112 -83786 -106 -83010
rect -152 -83798 -106 -83786
rect 106 -83010 152 -82998
rect 106 -83786 112 -83010
rect 146 -83786 152 -83010
rect 106 -83798 152 -83786
rect -96 -83845 96 -83839
rect -96 -83879 -84 -83845
rect 84 -83879 96 -83845
rect -96 -83885 96 -83879
rect -96 -83953 96 -83947
rect -96 -83987 -84 -83953
rect 84 -83987 96 -83953
rect -96 -83993 96 -83987
rect -152 -84046 -106 -84034
rect -152 -84822 -146 -84046
rect -112 -84822 -106 -84046
rect -152 -84834 -106 -84822
rect 106 -84046 152 -84034
rect 106 -84822 112 -84046
rect 146 -84822 152 -84046
rect 106 -84834 152 -84822
rect -96 -84881 96 -84875
rect -96 -84915 -84 -84881
rect 84 -84915 96 -84881
rect -96 -84921 96 -84915
rect -96 -84989 96 -84983
rect -96 -85023 -84 -84989
rect 84 -85023 96 -84989
rect -96 -85029 96 -85023
rect -152 -85082 -106 -85070
rect -152 -85858 -146 -85082
rect -112 -85858 -106 -85082
rect -152 -85870 -106 -85858
rect 106 -85082 152 -85070
rect 106 -85858 112 -85082
rect 146 -85858 152 -85082
rect 106 -85870 152 -85858
rect -96 -85917 96 -85911
rect -96 -85951 -84 -85917
rect 84 -85951 96 -85917
rect -96 -85957 96 -85951
rect -96 -86025 96 -86019
rect -96 -86059 -84 -86025
rect 84 -86059 96 -86025
rect -96 -86065 96 -86059
rect -152 -86118 -106 -86106
rect -152 -86894 -146 -86118
rect -112 -86894 -106 -86118
rect -152 -86906 -106 -86894
rect 106 -86118 152 -86106
rect 106 -86894 112 -86118
rect 146 -86894 152 -86118
rect 106 -86906 152 -86894
rect -96 -86953 96 -86947
rect -96 -86987 -84 -86953
rect 84 -86987 96 -86953
rect -96 -86993 96 -86987
rect -96 -87061 96 -87055
rect -96 -87095 -84 -87061
rect 84 -87095 96 -87061
rect -96 -87101 96 -87095
rect -152 -87154 -106 -87142
rect -152 -87930 -146 -87154
rect -112 -87930 -106 -87154
rect -152 -87942 -106 -87930
rect 106 -87154 152 -87142
rect 106 -87930 112 -87154
rect 146 -87930 152 -87154
rect 106 -87942 152 -87930
rect -96 -87989 96 -87983
rect -96 -88023 -84 -87989
rect 84 -88023 96 -87989
rect -96 -88029 96 -88023
rect -96 -88097 96 -88091
rect -96 -88131 -84 -88097
rect 84 -88131 96 -88097
rect -96 -88137 96 -88131
rect -152 -88190 -106 -88178
rect -152 -88966 -146 -88190
rect -112 -88966 -106 -88190
rect -152 -88978 -106 -88966
rect 106 -88190 152 -88178
rect 106 -88966 112 -88190
rect 146 -88966 152 -88190
rect 106 -88978 152 -88966
rect -96 -89025 96 -89019
rect -96 -89059 -84 -89025
rect 84 -89059 96 -89025
rect -96 -89065 96 -89059
rect -96 -89133 96 -89127
rect -96 -89167 -84 -89133
rect 84 -89167 96 -89133
rect -96 -89173 96 -89167
rect -152 -89226 -106 -89214
rect -152 -90002 -146 -89226
rect -112 -90002 -106 -89226
rect -152 -90014 -106 -90002
rect 106 -89226 152 -89214
rect 106 -90002 112 -89226
rect 146 -90002 152 -89226
rect 106 -90014 152 -90002
rect -96 -90061 96 -90055
rect -96 -90095 -84 -90061
rect 84 -90095 96 -90061
rect -96 -90101 96 -90095
rect -96 -90169 96 -90163
rect -96 -90203 -84 -90169
rect 84 -90203 96 -90169
rect -96 -90209 96 -90203
rect -152 -90262 -106 -90250
rect -152 -91038 -146 -90262
rect -112 -91038 -106 -90262
rect -152 -91050 -106 -91038
rect 106 -90262 152 -90250
rect 106 -91038 112 -90262
rect 146 -91038 152 -90262
rect 106 -91050 152 -91038
rect -96 -91097 96 -91091
rect -96 -91131 -84 -91097
rect 84 -91131 96 -91097
rect -96 -91137 96 -91131
rect -96 -91205 96 -91199
rect -96 -91239 -84 -91205
rect 84 -91239 96 -91205
rect -96 -91245 96 -91239
rect -152 -91298 -106 -91286
rect -152 -92074 -146 -91298
rect -112 -92074 -106 -91298
rect -152 -92086 -106 -92074
rect 106 -91298 152 -91286
rect 106 -92074 112 -91298
rect 146 -92074 152 -91298
rect 106 -92086 152 -92074
rect -96 -92133 96 -92127
rect -96 -92167 -84 -92133
rect 84 -92167 96 -92133
rect -96 -92173 96 -92167
rect -96 -92241 96 -92235
rect -96 -92275 -84 -92241
rect 84 -92275 96 -92241
rect -96 -92281 96 -92275
rect -152 -92334 -106 -92322
rect -152 -93110 -146 -92334
rect -112 -93110 -106 -92334
rect -152 -93122 -106 -93110
rect 106 -92334 152 -92322
rect 106 -93110 112 -92334
rect 146 -93110 152 -92334
rect 106 -93122 152 -93110
rect -96 -93169 96 -93163
rect -96 -93203 -84 -93169
rect 84 -93203 96 -93169
rect -96 -93209 96 -93203
rect -96 -93277 96 -93271
rect -96 -93311 -84 -93277
rect 84 -93311 96 -93277
rect -96 -93317 96 -93311
rect -152 -93370 -106 -93358
rect -152 -94146 -146 -93370
rect -112 -94146 -106 -93370
rect -152 -94158 -106 -94146
rect 106 -93370 152 -93358
rect 106 -94146 112 -93370
rect 146 -94146 152 -93370
rect 106 -94158 152 -94146
rect -96 -94205 96 -94199
rect -96 -94239 -84 -94205
rect 84 -94239 96 -94205
rect -96 -94245 96 -94239
rect -96 -94313 96 -94307
rect -96 -94347 -84 -94313
rect 84 -94347 96 -94313
rect -96 -94353 96 -94347
rect -152 -94406 -106 -94394
rect -152 -95182 -146 -94406
rect -112 -95182 -106 -94406
rect -152 -95194 -106 -95182
rect 106 -94406 152 -94394
rect 106 -95182 112 -94406
rect 146 -95182 152 -94406
rect 106 -95194 152 -95182
rect -96 -95241 96 -95235
rect -96 -95275 -84 -95241
rect 84 -95275 96 -95241
rect -96 -95281 96 -95275
rect -96 -95349 96 -95343
rect -96 -95383 -84 -95349
rect 84 -95383 96 -95349
rect -96 -95389 96 -95383
rect -152 -95442 -106 -95430
rect -152 -96218 -146 -95442
rect -112 -96218 -106 -95442
rect -152 -96230 -106 -96218
rect 106 -95442 152 -95430
rect 106 -96218 112 -95442
rect 146 -96218 152 -95442
rect 106 -96230 152 -96218
rect -96 -96277 96 -96271
rect -96 -96311 -84 -96277
rect 84 -96311 96 -96277
rect -96 -96317 96 -96311
rect -96 -96385 96 -96379
rect -96 -96419 -84 -96385
rect 84 -96419 96 -96385
rect -96 -96425 96 -96419
rect -152 -96478 -106 -96466
rect -152 -97254 -146 -96478
rect -112 -97254 -106 -96478
rect -152 -97266 -106 -97254
rect 106 -96478 152 -96466
rect 106 -97254 112 -96478
rect 146 -97254 152 -96478
rect 106 -97266 152 -97254
rect -96 -97313 96 -97307
rect -96 -97347 -84 -97313
rect 84 -97347 96 -97313
rect -96 -97353 96 -97347
rect -96 -97421 96 -97415
rect -96 -97455 -84 -97421
rect 84 -97455 96 -97421
rect -96 -97461 96 -97455
rect -152 -97514 -106 -97502
rect -152 -98290 -146 -97514
rect -112 -98290 -106 -97514
rect -152 -98302 -106 -98290
rect 106 -97514 152 -97502
rect 106 -98290 112 -97514
rect 146 -98290 152 -97514
rect 106 -98302 152 -98290
rect -96 -98349 96 -98343
rect -96 -98383 -84 -98349
rect 84 -98383 96 -98349
rect -96 -98389 96 -98383
rect -96 -98457 96 -98451
rect -96 -98491 -84 -98457
rect 84 -98491 96 -98457
rect -96 -98497 96 -98491
rect -152 -98550 -106 -98538
rect -152 -99326 -146 -98550
rect -112 -99326 -106 -98550
rect -152 -99338 -106 -99326
rect 106 -98550 152 -98538
rect 106 -99326 112 -98550
rect 146 -99326 152 -98550
rect 106 -99338 152 -99326
rect -96 -99385 96 -99379
rect -96 -99419 -84 -99385
rect 84 -99419 96 -99385
rect -96 -99425 96 -99419
rect -96 -99493 96 -99487
rect -96 -99527 -84 -99493
rect 84 -99527 96 -99493
rect -96 -99533 96 -99527
rect -152 -99586 -106 -99574
rect -152 -100362 -146 -99586
rect -112 -100362 -106 -99586
rect -152 -100374 -106 -100362
rect 106 -99586 152 -99574
rect 106 -100362 112 -99586
rect 146 -100362 152 -99586
rect 106 -100374 152 -100362
rect -96 -100421 96 -100415
rect -96 -100455 -84 -100421
rect 84 -100455 96 -100421
rect -96 -100461 96 -100455
rect -96 -100529 96 -100523
rect -96 -100563 -84 -100529
rect 84 -100563 96 -100529
rect -96 -100569 96 -100563
rect -152 -100622 -106 -100610
rect -152 -101398 -146 -100622
rect -112 -101398 -106 -100622
rect -152 -101410 -106 -101398
rect 106 -100622 152 -100610
rect 106 -101398 112 -100622
rect 146 -101398 152 -100622
rect 106 -101410 152 -101398
rect -96 -101457 96 -101451
rect -96 -101491 -84 -101457
rect 84 -101491 96 -101457
rect -96 -101497 96 -101491
rect -96 -101565 96 -101559
rect -96 -101599 -84 -101565
rect 84 -101599 96 -101565
rect -96 -101605 96 -101599
rect -152 -101658 -106 -101646
rect -152 -102434 -146 -101658
rect -112 -102434 -106 -101658
rect -152 -102446 -106 -102434
rect 106 -101658 152 -101646
rect 106 -102434 112 -101658
rect 146 -102434 152 -101658
rect 106 -102446 152 -102434
rect -96 -102493 96 -102487
rect -96 -102527 -84 -102493
rect 84 -102527 96 -102493
rect -96 -102533 96 -102527
rect -96 -102601 96 -102595
rect -96 -102635 -84 -102601
rect 84 -102635 96 -102601
rect -96 -102641 96 -102635
rect -152 -102694 -106 -102682
rect -152 -103470 -146 -102694
rect -112 -103470 -106 -102694
rect -152 -103482 -106 -103470
rect 106 -102694 152 -102682
rect 106 -103470 112 -102694
rect 146 -103470 152 -102694
rect 106 -103482 152 -103470
rect -96 -103529 96 -103523
rect -96 -103563 -84 -103529
rect 84 -103563 96 -103529
rect -96 -103569 96 -103563
rect -96 -103637 96 -103631
rect -96 -103671 -84 -103637
rect 84 -103671 96 -103637
rect -96 -103677 96 -103671
rect -152 -103730 -106 -103718
rect -152 -104506 -146 -103730
rect -112 -104506 -106 -103730
rect -152 -104518 -106 -104506
rect 106 -103730 152 -103718
rect 106 -104506 112 -103730
rect 146 -104506 152 -103730
rect 106 -104518 152 -104506
rect -96 -104565 96 -104559
rect -96 -104599 -84 -104565
rect 84 -104599 96 -104565
rect -96 -104605 96 -104599
rect -96 -104673 96 -104667
rect -96 -104707 -84 -104673
rect 84 -104707 96 -104673
rect -96 -104713 96 -104707
rect -152 -104766 -106 -104754
rect -152 -105542 -146 -104766
rect -112 -105542 -106 -104766
rect -152 -105554 -106 -105542
rect 106 -104766 152 -104754
rect 106 -105542 112 -104766
rect 146 -105542 152 -104766
rect 106 -105554 152 -105542
rect -96 -105601 96 -105595
rect -96 -105635 -84 -105601
rect 84 -105635 96 -105601
rect -96 -105641 96 -105635
rect -96 -105709 96 -105703
rect -96 -105743 -84 -105709
rect 84 -105743 96 -105709
rect -96 -105749 96 -105743
rect -152 -105802 -106 -105790
rect -152 -106578 -146 -105802
rect -112 -106578 -106 -105802
rect -152 -106590 -106 -106578
rect 106 -105802 152 -105790
rect 106 -106578 112 -105802
rect 146 -106578 152 -105802
rect 106 -106590 152 -106578
rect -96 -106637 96 -106631
rect -96 -106671 -84 -106637
rect 84 -106671 96 -106637
rect -96 -106677 96 -106671
rect -96 -106745 96 -106739
rect -96 -106779 -84 -106745
rect 84 -106779 96 -106745
rect -96 -106785 96 -106779
rect -152 -106838 -106 -106826
rect -152 -107614 -146 -106838
rect -112 -107614 -106 -106838
rect -152 -107626 -106 -107614
rect 106 -106838 152 -106826
rect 106 -107614 112 -106838
rect 146 -107614 152 -106838
rect 106 -107626 152 -107614
rect -96 -107673 96 -107667
rect -96 -107707 -84 -107673
rect 84 -107707 96 -107673
rect -96 -107713 96 -107707
rect -96 -107781 96 -107775
rect -96 -107815 -84 -107781
rect 84 -107815 96 -107781
rect -96 -107821 96 -107815
rect -152 -107874 -106 -107862
rect -152 -108650 -146 -107874
rect -112 -108650 -106 -107874
rect -152 -108662 -106 -108650
rect 106 -107874 152 -107862
rect 106 -108650 112 -107874
rect 146 -108650 152 -107874
rect 106 -108662 152 -108650
rect -96 -108709 96 -108703
rect -96 -108743 -84 -108709
rect 84 -108743 96 -108709
rect -96 -108749 96 -108743
rect -96 -108817 96 -108811
rect -96 -108851 -84 -108817
rect 84 -108851 96 -108817
rect -96 -108857 96 -108851
rect -152 -108910 -106 -108898
rect -152 -109686 -146 -108910
rect -112 -109686 -106 -108910
rect -152 -109698 -106 -109686
rect 106 -108910 152 -108898
rect 106 -109686 112 -108910
rect 146 -109686 152 -108910
rect 106 -109698 152 -109686
rect -96 -109745 96 -109739
rect -96 -109779 -84 -109745
rect 84 -109779 96 -109745
rect -96 -109785 96 -109779
rect -96 -109853 96 -109847
rect -96 -109887 -84 -109853
rect 84 -109887 96 -109853
rect -96 -109893 96 -109887
rect -152 -109946 -106 -109934
rect -152 -110722 -146 -109946
rect -112 -110722 -106 -109946
rect -152 -110734 -106 -110722
rect 106 -109946 152 -109934
rect 106 -110722 112 -109946
rect 146 -110722 152 -109946
rect 106 -110734 152 -110722
rect -96 -110781 96 -110775
rect -96 -110815 -84 -110781
rect 84 -110815 96 -110781
rect -96 -110821 96 -110815
rect -96 -110889 96 -110883
rect -96 -110923 -84 -110889
rect 84 -110923 96 -110889
rect -96 -110929 96 -110923
rect -152 -110982 -106 -110970
rect -152 -111758 -146 -110982
rect -112 -111758 -106 -110982
rect -152 -111770 -106 -111758
rect 106 -110982 152 -110970
rect 106 -111758 112 -110982
rect 146 -111758 152 -110982
rect 106 -111770 152 -111758
rect -96 -111817 96 -111811
rect -96 -111851 -84 -111817
rect 84 -111851 96 -111817
rect -96 -111857 96 -111851
rect -96 -111925 96 -111919
rect -96 -111959 -84 -111925
rect 84 -111959 96 -111925
rect -96 -111965 96 -111959
rect -152 -112018 -106 -112006
rect -152 -112794 -146 -112018
rect -112 -112794 -106 -112018
rect -152 -112806 -106 -112794
rect 106 -112018 152 -112006
rect 106 -112794 112 -112018
rect 146 -112794 152 -112018
rect 106 -112806 152 -112794
rect -96 -112853 96 -112847
rect -96 -112887 -84 -112853
rect 84 -112887 96 -112853
rect -96 -112893 96 -112887
rect -96 -112961 96 -112955
rect -96 -112995 -84 -112961
rect 84 -112995 96 -112961
rect -96 -113001 96 -112995
rect -152 -113054 -106 -113042
rect -152 -113830 -146 -113054
rect -112 -113830 -106 -113054
rect -152 -113842 -106 -113830
rect 106 -113054 152 -113042
rect 106 -113830 112 -113054
rect 146 -113830 152 -113054
rect 106 -113842 152 -113830
rect -96 -113889 96 -113883
rect -96 -113923 -84 -113889
rect 84 -113923 96 -113889
rect -96 -113929 96 -113923
rect -96 -113997 96 -113991
rect -96 -114031 -84 -113997
rect 84 -114031 96 -113997
rect -96 -114037 96 -114031
rect -152 -114090 -106 -114078
rect -152 -114866 -146 -114090
rect -112 -114866 -106 -114090
rect -152 -114878 -106 -114866
rect 106 -114090 152 -114078
rect 106 -114866 112 -114090
rect 146 -114866 152 -114090
rect 106 -114878 152 -114866
rect -96 -114925 96 -114919
rect -96 -114959 -84 -114925
rect 84 -114959 96 -114925
rect -96 -114965 96 -114959
rect -96 -115033 96 -115027
rect -96 -115067 -84 -115033
rect 84 -115067 96 -115033
rect -96 -115073 96 -115067
rect -152 -115126 -106 -115114
rect -152 -115902 -146 -115126
rect -112 -115902 -106 -115126
rect -152 -115914 -106 -115902
rect 106 -115126 152 -115114
rect 106 -115902 112 -115126
rect 146 -115902 152 -115126
rect 106 -115914 152 -115902
rect -96 -115961 96 -115955
rect -96 -115995 -84 -115961
rect 84 -115995 96 -115961
rect -96 -116001 96 -115995
rect -96 -116069 96 -116063
rect -96 -116103 -84 -116069
rect 84 -116103 96 -116069
rect -96 -116109 96 -116103
rect -152 -116162 -106 -116150
rect -152 -116938 -146 -116162
rect -112 -116938 -106 -116162
rect -152 -116950 -106 -116938
rect 106 -116162 152 -116150
rect 106 -116938 112 -116162
rect 146 -116938 152 -116162
rect 106 -116950 152 -116938
rect -96 -116997 96 -116991
rect -96 -117031 -84 -116997
rect 84 -117031 96 -116997
rect -96 -117037 96 -117031
rect -96 -117105 96 -117099
rect -96 -117139 -84 -117105
rect 84 -117139 96 -117105
rect -96 -117145 96 -117139
rect -152 -117198 -106 -117186
rect -152 -117974 -146 -117198
rect -112 -117974 -106 -117198
rect -152 -117986 -106 -117974
rect 106 -117198 152 -117186
rect 106 -117974 112 -117198
rect 146 -117974 152 -117198
rect 106 -117986 152 -117974
rect -96 -118033 96 -118027
rect -96 -118067 -84 -118033
rect 84 -118067 96 -118033
rect -96 -118073 96 -118067
rect -96 -118141 96 -118135
rect -96 -118175 -84 -118141
rect 84 -118175 96 -118141
rect -96 -118181 96 -118175
rect -152 -118234 -106 -118222
rect -152 -119010 -146 -118234
rect -112 -119010 -106 -118234
rect -152 -119022 -106 -119010
rect 106 -118234 152 -118222
rect 106 -119010 112 -118234
rect 146 -119010 152 -118234
rect 106 -119022 152 -119010
rect -96 -119069 96 -119063
rect -96 -119103 -84 -119069
rect 84 -119103 96 -119069
rect -96 -119109 96 -119103
rect -96 -119177 96 -119171
rect -96 -119211 -84 -119177
rect 84 -119211 96 -119177
rect -96 -119217 96 -119211
rect -152 -119270 -106 -119258
rect -152 -120046 -146 -119270
rect -112 -120046 -106 -119270
rect -152 -120058 -106 -120046
rect 106 -119270 152 -119258
rect 106 -120046 112 -119270
rect 146 -120046 152 -119270
rect 106 -120058 152 -120046
rect -96 -120105 96 -120099
rect -96 -120139 -84 -120105
rect 84 -120139 96 -120105
rect -96 -120145 96 -120139
rect -96 -120213 96 -120207
rect -96 -120247 -84 -120213
rect 84 -120247 96 -120213
rect -96 -120253 96 -120247
rect -152 -120306 -106 -120294
rect -152 -121082 -146 -120306
rect -112 -121082 -106 -120306
rect -152 -121094 -106 -121082
rect 106 -120306 152 -120294
rect 106 -121082 112 -120306
rect 146 -121082 152 -120306
rect 106 -121094 152 -121082
rect -96 -121141 96 -121135
rect -96 -121175 -84 -121141
rect 84 -121175 96 -121141
rect -96 -121181 96 -121175
rect -96 -121249 96 -121243
rect -96 -121283 -84 -121249
rect 84 -121283 96 -121249
rect -96 -121289 96 -121283
rect -152 -121342 -106 -121330
rect -152 -122118 -146 -121342
rect -112 -122118 -106 -121342
rect -152 -122130 -106 -122118
rect 106 -121342 152 -121330
rect 106 -122118 112 -121342
rect 146 -122118 152 -121342
rect 106 -122130 152 -122118
rect -96 -122177 96 -122171
rect -96 -122211 -84 -122177
rect 84 -122211 96 -122177
rect -96 -122217 96 -122211
rect -96 -122285 96 -122279
rect -96 -122319 -84 -122285
rect 84 -122319 96 -122285
rect -96 -122325 96 -122319
rect -152 -122378 -106 -122366
rect -152 -123154 -146 -122378
rect -112 -123154 -106 -122378
rect -152 -123166 -106 -123154
rect 106 -122378 152 -122366
rect 106 -123154 112 -122378
rect 146 -123154 152 -122378
rect 106 -123166 152 -123154
rect -96 -123213 96 -123207
rect -96 -123247 -84 -123213
rect 84 -123247 96 -123213
rect -96 -123253 96 -123247
rect -96 -123321 96 -123315
rect -96 -123355 -84 -123321
rect 84 -123355 96 -123321
rect -96 -123361 96 -123355
rect -152 -123414 -106 -123402
rect -152 -124190 -146 -123414
rect -112 -124190 -106 -123414
rect -152 -124202 -106 -124190
rect 106 -123414 152 -123402
rect 106 -124190 112 -123414
rect 146 -124190 152 -123414
rect 106 -124202 152 -124190
rect -96 -124249 96 -124243
rect -96 -124283 -84 -124249
rect 84 -124283 96 -124249
rect -96 -124289 96 -124283
rect -96 -124357 96 -124351
rect -96 -124391 -84 -124357
rect 84 -124391 96 -124357
rect -96 -124397 96 -124391
rect -152 -124450 -106 -124438
rect -152 -125226 -146 -124450
rect -112 -125226 -106 -124450
rect -152 -125238 -106 -125226
rect 106 -124450 152 -124438
rect 106 -125226 112 -124450
rect 146 -125226 152 -124450
rect 106 -125238 152 -125226
rect -96 -125285 96 -125279
rect -96 -125319 -84 -125285
rect 84 -125319 96 -125285
rect -96 -125325 96 -125319
rect -96 -125393 96 -125387
rect -96 -125427 -84 -125393
rect 84 -125427 96 -125393
rect -96 -125433 96 -125427
rect -152 -125486 -106 -125474
rect -152 -126262 -146 -125486
rect -112 -126262 -106 -125486
rect -152 -126274 -106 -126262
rect 106 -125486 152 -125474
rect 106 -126262 112 -125486
rect 146 -126262 152 -125486
rect 106 -126274 152 -126262
rect -96 -126321 96 -126315
rect -96 -126355 -84 -126321
rect 84 -126355 96 -126321
rect -96 -126361 96 -126355
rect -96 -126429 96 -126423
rect -96 -126463 -84 -126429
rect 84 -126463 96 -126429
rect -96 -126469 96 -126463
rect -152 -126522 -106 -126510
rect -152 -127298 -146 -126522
rect -112 -127298 -106 -126522
rect -152 -127310 -106 -127298
rect 106 -126522 152 -126510
rect 106 -127298 112 -126522
rect 146 -127298 152 -126522
rect 106 -127310 152 -127298
rect -96 -127357 96 -127351
rect -96 -127391 -84 -127357
rect 84 -127391 96 -127357
rect -96 -127397 96 -127391
rect -96 -127465 96 -127459
rect -96 -127499 -84 -127465
rect 84 -127499 96 -127465
rect -96 -127505 96 -127499
rect -152 -127558 -106 -127546
rect -152 -128334 -146 -127558
rect -112 -128334 -106 -127558
rect -152 -128346 -106 -128334
rect 106 -127558 152 -127546
rect 106 -128334 112 -127558
rect 146 -128334 152 -127558
rect 106 -128346 152 -128334
rect -96 -128393 96 -128387
rect -96 -128427 -84 -128393
rect 84 -128427 96 -128393
rect -96 -128433 96 -128427
rect -96 -128501 96 -128495
rect -96 -128535 -84 -128501
rect 84 -128535 96 -128501
rect -96 -128541 96 -128535
rect -152 -128594 -106 -128582
rect -152 -129370 -146 -128594
rect -112 -129370 -106 -128594
rect -152 -129382 -106 -129370
rect 106 -128594 152 -128582
rect 106 -129370 112 -128594
rect 146 -129370 152 -128594
rect 106 -129382 152 -129370
rect -96 -129429 96 -129423
rect -96 -129463 -84 -129429
rect 84 -129463 96 -129429
rect -96 -129469 96 -129463
rect -96 -129537 96 -129531
rect -96 -129571 -84 -129537
rect 84 -129571 96 -129537
rect -96 -129577 96 -129571
rect -152 -129630 -106 -129618
rect -152 -130406 -146 -129630
rect -112 -130406 -106 -129630
rect -152 -130418 -106 -130406
rect 106 -129630 152 -129618
rect 106 -130406 112 -129630
rect 146 -130406 152 -129630
rect 106 -130418 152 -130406
rect -96 -130465 96 -130459
rect -96 -130499 -84 -130465
rect 84 -130499 96 -130465
rect -96 -130505 96 -130499
rect -96 -130573 96 -130567
rect -96 -130607 -84 -130573
rect 84 -130607 96 -130573
rect -96 -130613 96 -130607
rect -152 -130666 -106 -130654
rect -152 -131442 -146 -130666
rect -112 -131442 -106 -130666
rect -152 -131454 -106 -131442
rect 106 -130666 152 -130654
rect 106 -131442 112 -130666
rect 146 -131442 152 -130666
rect 106 -131454 152 -131442
rect -96 -131501 96 -131495
rect -96 -131535 -84 -131501
rect 84 -131535 96 -131501
rect -96 -131541 96 -131535
rect -96 -131609 96 -131603
rect -96 -131643 -84 -131609
rect 84 -131643 96 -131609
rect -96 -131649 96 -131643
rect -152 -131702 -106 -131690
rect -152 -132478 -146 -131702
rect -112 -132478 -106 -131702
rect -152 -132490 -106 -132478
rect 106 -131702 152 -131690
rect 106 -132478 112 -131702
rect 146 -132478 152 -131702
rect 106 -132490 152 -132478
rect -96 -132537 96 -132531
rect -96 -132571 -84 -132537
rect 84 -132571 96 -132537
rect -96 -132577 96 -132571
<< properties >>
string FIXED_BBOX -263 -132692 263 132692
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 1.0 m 256 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
