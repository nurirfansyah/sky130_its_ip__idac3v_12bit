magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 3344 -2965 3460 -2899
rect 6688 -2965 6804 -2899
rect 10032 -2965 10148 -2899
rect 13376 -2965 13492 -2899
rect 16720 -2965 16836 -2899
rect 20064 -2965 20180 -2899
rect 23408 -2965 23524 -2899
rect 26752 -2965 26868 -2899
rect 30096 -2965 30212 -2899
rect 33440 -2965 33556 -2899
rect 36784 -2965 36900 -2899
rect 40128 -2965 40244 -2899
rect 43472 -2965 43588 -2899
rect 46816 -2965 46932 -2899
rect 50160 -2965 50276 -2899
rect 56848 -2965 56964 -2899
rect 60192 -2965 60308 -2899
rect 63536 -2965 63652 -2899
rect 66880 -2965 66996 -2899
rect 70224 -2965 70340 -2899
rect 73568 -2965 73684 -2899
rect 76912 -2965 77028 -2899
rect 80256 -2965 80372 -2899
rect 83600 -2965 83716 -2899
rect 86944 -2965 87060 -2899
rect 90288 -2965 90404 -2899
rect 93632 -2965 93748 -2899
rect 96976 -2965 97092 -2899
rect 100320 -2965 100436 -2899
rect 103664 -2965 103780 -2899
rect 3460 -3219 3846 -3153
rect 6804 -3219 7190 -3153
rect 10148 -3219 10534 -3153
rect 13492 -3219 13878 -3153
rect 16836 -3219 17222 -3153
rect 20180 -3219 20566 -3153
rect 23524 -3219 23910 -3153
rect 26868 -3219 27254 -3153
rect 30212 -3219 30598 -3153
rect 33556 -3219 33942 -3153
rect 36900 -3219 37286 -3153
rect 40244 -3219 40630 -3153
rect 43588 -3219 43974 -3153
rect 46932 -3219 47318 -3153
rect 50276 -3219 50662 -3153
rect 3196 -3232 3206 -3219
rect 3130 -3274 3206 -3232
rect 3258 -3274 3846 -3219
rect 6540 -3232 6550 -3219
rect 3130 -3277 3846 -3274
rect 3130 -3514 3274 -3277
rect 3460 -3299 3846 -3277
rect 3384 -3385 3846 -3299
rect 6474 -3274 6550 -3232
rect 6602 -3274 7190 -3219
rect 9884 -3232 9894 -3219
rect 6474 -3277 7190 -3274
rect 3388 -3393 3588 -3385
rect 3404 -3397 3572 -3393
rect 3130 -3600 3304 -3514
rect 3330 -3574 3430 -3450
rect 6474 -3514 6618 -3277
rect 6804 -3299 7190 -3277
rect 6728 -3385 7190 -3299
rect 9818 -3274 9894 -3232
rect 9946 -3274 10534 -3219
rect 13228 -3232 13238 -3219
rect 9818 -3277 10534 -3274
rect 6732 -3393 6932 -3385
rect 6748 -3397 6916 -3393
rect 3330 -3628 3332 -3574
rect 6474 -3600 6648 -3514
rect 6674 -3574 6774 -3450
rect 9818 -3514 9962 -3277
rect 10148 -3299 10534 -3277
rect 10072 -3385 10534 -3299
rect 13162 -3274 13238 -3232
rect 13290 -3274 13878 -3219
rect 16572 -3232 16582 -3219
rect 13162 -3277 13878 -3274
rect 10076 -3393 10276 -3385
rect 10092 -3397 10260 -3393
rect 6674 -3628 6676 -3574
rect 9818 -3600 9992 -3514
rect 10018 -3574 10118 -3450
rect 13162 -3514 13306 -3277
rect 13492 -3299 13878 -3277
rect 13416 -3385 13878 -3299
rect 16506 -3274 16582 -3232
rect 16634 -3274 17222 -3219
rect 19916 -3232 19926 -3219
rect 16506 -3277 17222 -3274
rect 13420 -3393 13620 -3385
rect 13436 -3397 13604 -3393
rect 10018 -3628 10020 -3574
rect 13162 -3600 13336 -3514
rect 13362 -3574 13462 -3450
rect 16506 -3514 16650 -3277
rect 16836 -3299 17222 -3277
rect 16760 -3385 17222 -3299
rect 19850 -3274 19926 -3232
rect 19978 -3274 20566 -3219
rect 23260 -3232 23270 -3219
rect 19850 -3277 20566 -3274
rect 16764 -3393 16964 -3385
rect 16780 -3397 16948 -3393
rect 13362 -3628 13364 -3574
rect 16506 -3600 16680 -3514
rect 16706 -3574 16806 -3450
rect 19850 -3514 19994 -3277
rect 20180 -3299 20566 -3277
rect 20104 -3385 20566 -3299
rect 23194 -3274 23270 -3232
rect 23322 -3274 23910 -3219
rect 26604 -3232 26614 -3219
rect 23194 -3277 23910 -3274
rect 20108 -3393 20308 -3385
rect 20124 -3397 20292 -3393
rect 16706 -3628 16708 -3574
rect 19850 -3600 20024 -3514
rect 20050 -3574 20150 -3450
rect 23194 -3514 23338 -3277
rect 23524 -3299 23910 -3277
rect 23448 -3385 23910 -3299
rect 26538 -3274 26614 -3232
rect 26666 -3274 27254 -3219
rect 29948 -3232 29958 -3219
rect 26538 -3277 27254 -3274
rect 23452 -3393 23652 -3385
rect 23468 -3397 23636 -3393
rect 20050 -3628 20052 -3574
rect 23194 -3600 23368 -3514
rect 23394 -3574 23494 -3450
rect 26538 -3514 26682 -3277
rect 26868 -3299 27254 -3277
rect 26792 -3385 27254 -3299
rect 29882 -3274 29958 -3232
rect 30010 -3274 30598 -3219
rect 33292 -3232 33302 -3219
rect 29882 -3277 30598 -3274
rect 26796 -3393 26996 -3385
rect 26812 -3397 26980 -3393
rect 23394 -3628 23396 -3574
rect 26538 -3600 26712 -3514
rect 26738 -3574 26838 -3450
rect 29882 -3514 30026 -3277
rect 30212 -3299 30598 -3277
rect 30136 -3385 30598 -3299
rect 33226 -3274 33302 -3232
rect 33354 -3274 33942 -3219
rect 36636 -3232 36646 -3219
rect 33226 -3277 33942 -3274
rect 30140 -3393 30340 -3385
rect 30156 -3397 30324 -3393
rect 26738 -3628 26740 -3574
rect 29882 -3600 30056 -3514
rect 30082 -3574 30182 -3450
rect 33226 -3514 33370 -3277
rect 33556 -3299 33942 -3277
rect 33480 -3385 33942 -3299
rect 36570 -3274 36646 -3232
rect 36698 -3274 37286 -3219
rect 39980 -3232 39990 -3219
rect 36570 -3277 37286 -3274
rect 33484 -3393 33684 -3385
rect 33500 -3397 33668 -3393
rect 30082 -3628 30084 -3574
rect 33226 -3600 33400 -3514
rect 33426 -3574 33526 -3450
rect 36570 -3514 36714 -3277
rect 36900 -3299 37286 -3277
rect 36824 -3385 37286 -3299
rect 39914 -3274 39990 -3232
rect 40042 -3274 40630 -3219
rect 43324 -3232 43334 -3219
rect 39914 -3277 40630 -3274
rect 36828 -3393 37028 -3385
rect 36844 -3397 37012 -3393
rect 33426 -3628 33428 -3574
rect 36570 -3600 36744 -3514
rect 36770 -3574 36870 -3450
rect 39914 -3514 40058 -3277
rect 40244 -3299 40630 -3277
rect 40168 -3385 40630 -3299
rect 43258 -3274 43334 -3232
rect 43386 -3274 43974 -3219
rect 46668 -3232 46678 -3219
rect 43258 -3277 43974 -3274
rect 40172 -3393 40372 -3385
rect 40188 -3397 40356 -3393
rect 36770 -3628 36772 -3574
rect 39914 -3600 40088 -3514
rect 40114 -3574 40214 -3450
rect 43258 -3514 43402 -3277
rect 43588 -3299 43974 -3277
rect 43512 -3385 43974 -3299
rect 46602 -3274 46678 -3232
rect 46730 -3274 47318 -3219
rect 50012 -3232 50022 -3219
rect 46602 -3277 47318 -3274
rect 43516 -3393 43716 -3385
rect 43532 -3397 43700 -3393
rect 40114 -3628 40116 -3574
rect 43258 -3600 43432 -3514
rect 43458 -3574 43558 -3450
rect 46602 -3514 46746 -3277
rect 46932 -3299 47318 -3277
rect 46856 -3385 47318 -3299
rect 49946 -3274 50022 -3232
rect 50074 -3274 50662 -3219
rect 49946 -3277 50662 -3274
rect 46860 -3393 47060 -3385
rect 46876 -3397 47044 -3393
rect 43458 -3628 43460 -3574
rect 46602 -3600 46776 -3514
rect 46802 -3574 46902 -3450
rect 49946 -3514 50090 -3277
rect 50276 -3299 50662 -3277
rect 50200 -3385 50662 -3299
rect 56700 -3232 56710 -3219
rect 50204 -3393 50404 -3385
rect 50220 -3397 50388 -3393
rect 46802 -3628 46804 -3574
rect 49946 -3600 50120 -3514
rect 50146 -3574 50246 -3450
rect 56634 -3274 56710 -3232
rect 56762 -3274 56964 -3219
rect 50146 -3628 50148 -3574
rect 56778 -3277 56964 -3274
rect 60308 -3219 60694 -3153
rect 63652 -3219 64038 -3153
rect 66996 -3219 67382 -3153
rect 70340 -3219 70726 -3153
rect 73684 -3219 74070 -3153
rect 77028 -3219 77414 -3153
rect 80372 -3219 80758 -3153
rect 83716 -3219 84102 -3153
rect 87060 -3219 87446 -3153
rect 90404 -3219 90790 -3153
rect 93748 -3219 94134 -3153
rect 97092 -3219 97478 -3153
rect 100436 -3219 100822 -3153
rect 103780 -3219 104166 -3153
rect 60044 -3232 60054 -3219
rect 59978 -3274 60054 -3232
rect 60106 -3274 60694 -3219
rect 63388 -3232 63398 -3219
rect 59978 -3277 60694 -3274
rect 56892 -3393 57092 -3385
rect 56908 -3397 57076 -3393
rect 56834 -3574 56934 -3450
rect 59978 -3514 60122 -3277
rect 60308 -3299 60694 -3277
rect 60232 -3385 60694 -3299
rect 63322 -3274 63398 -3232
rect 63450 -3274 64038 -3219
rect 66732 -3232 66742 -3219
rect 63322 -3277 64038 -3274
rect 60236 -3393 60436 -3385
rect 60252 -3397 60420 -3393
rect 56834 -3628 56836 -3574
rect 59978 -3600 60152 -3514
rect 60178 -3574 60278 -3450
rect 63322 -3514 63466 -3277
rect 63652 -3299 64038 -3277
rect 63576 -3385 64038 -3299
rect 66666 -3274 66742 -3232
rect 66794 -3274 67382 -3219
rect 70076 -3232 70086 -3219
rect 66666 -3277 67382 -3274
rect 63580 -3393 63780 -3385
rect 63596 -3397 63764 -3393
rect 60178 -3628 60180 -3574
rect 63322 -3600 63496 -3514
rect 63522 -3574 63622 -3450
rect 66666 -3514 66810 -3277
rect 66996 -3299 67382 -3277
rect 66920 -3385 67382 -3299
rect 70010 -3274 70086 -3232
rect 70138 -3274 70726 -3219
rect 73420 -3232 73430 -3219
rect 70010 -3277 70726 -3274
rect 66924 -3393 67124 -3385
rect 66940 -3397 67108 -3393
rect 63522 -3628 63524 -3574
rect 66666 -3600 66840 -3514
rect 66866 -3574 66966 -3450
rect 70010 -3514 70154 -3277
rect 70340 -3299 70726 -3277
rect 70264 -3385 70726 -3299
rect 73354 -3274 73430 -3232
rect 73482 -3274 74070 -3219
rect 76764 -3232 76774 -3219
rect 73354 -3277 74070 -3274
rect 70268 -3393 70468 -3385
rect 70284 -3397 70452 -3393
rect 66866 -3628 66868 -3574
rect 70010 -3600 70184 -3514
rect 70210 -3574 70310 -3450
rect 73354 -3514 73498 -3277
rect 73684 -3299 74070 -3277
rect 73608 -3385 74070 -3299
rect 76698 -3274 76774 -3232
rect 76826 -3274 77414 -3219
rect 80108 -3232 80118 -3219
rect 76698 -3277 77414 -3274
rect 73612 -3393 73812 -3385
rect 73628 -3397 73796 -3393
rect 70210 -3628 70212 -3574
rect 73354 -3600 73528 -3514
rect 73554 -3574 73654 -3450
rect 76698 -3514 76842 -3277
rect 77028 -3299 77414 -3277
rect 76952 -3385 77414 -3299
rect 80042 -3274 80118 -3232
rect 80170 -3274 80758 -3219
rect 83452 -3232 83462 -3219
rect 80042 -3277 80758 -3274
rect 76956 -3393 77156 -3385
rect 76972 -3397 77140 -3393
rect 73554 -3628 73556 -3574
rect 76698 -3600 76872 -3514
rect 76898 -3574 76998 -3450
rect 80042 -3514 80186 -3277
rect 80372 -3299 80758 -3277
rect 80296 -3385 80758 -3299
rect 83386 -3274 83462 -3232
rect 83514 -3274 84102 -3219
rect 86796 -3232 86806 -3219
rect 83386 -3277 84102 -3274
rect 80300 -3393 80500 -3385
rect 80316 -3397 80484 -3393
rect 76898 -3628 76900 -3574
rect 80042 -3600 80216 -3514
rect 80242 -3574 80342 -3450
rect 83386 -3514 83530 -3277
rect 83716 -3299 84102 -3277
rect 83640 -3385 84102 -3299
rect 86730 -3274 86806 -3232
rect 86858 -3274 87446 -3219
rect 90140 -3232 90150 -3219
rect 86730 -3277 87446 -3274
rect 83644 -3393 83844 -3385
rect 83660 -3397 83828 -3393
rect 80242 -3628 80244 -3574
rect 83386 -3600 83560 -3514
rect 83586 -3574 83686 -3450
rect 86730 -3514 86874 -3277
rect 87060 -3299 87446 -3277
rect 86984 -3385 87446 -3299
rect 90074 -3274 90150 -3232
rect 90202 -3274 90790 -3219
rect 93484 -3232 93494 -3219
rect 90074 -3277 90790 -3274
rect 86988 -3393 87188 -3385
rect 87004 -3397 87172 -3393
rect 83586 -3628 83588 -3574
rect 86730 -3600 86904 -3514
rect 86930 -3574 87030 -3450
rect 90074 -3514 90218 -3277
rect 90404 -3299 90790 -3277
rect 90328 -3385 90790 -3299
rect 93418 -3274 93494 -3232
rect 93546 -3274 94134 -3219
rect 96828 -3232 96838 -3219
rect 93418 -3277 94134 -3274
rect 90332 -3393 90532 -3385
rect 90348 -3397 90516 -3393
rect 86930 -3628 86932 -3574
rect 90074 -3600 90248 -3514
rect 90274 -3574 90374 -3450
rect 93418 -3514 93562 -3277
rect 93748 -3299 94134 -3277
rect 93672 -3385 94134 -3299
rect 96762 -3274 96838 -3232
rect 96890 -3274 97478 -3219
rect 100172 -3232 100182 -3219
rect 96762 -3277 97478 -3274
rect 93676 -3393 93876 -3385
rect 93692 -3397 93860 -3393
rect 90274 -3628 90276 -3574
rect 93418 -3600 93592 -3514
rect 93618 -3574 93718 -3450
rect 96762 -3514 96906 -3277
rect 97092 -3299 97478 -3277
rect 97016 -3385 97478 -3299
rect 100106 -3274 100182 -3232
rect 100234 -3274 100822 -3219
rect 103516 -3232 103526 -3219
rect 100106 -3277 100822 -3274
rect 97020 -3393 97220 -3385
rect 97036 -3397 97204 -3393
rect 93618 -3628 93620 -3574
rect 96762 -3600 96936 -3514
rect 96962 -3574 97062 -3450
rect 100106 -3514 100250 -3277
rect 100436 -3299 100822 -3277
rect 100360 -3385 100822 -3299
rect 103450 -3274 103526 -3232
rect 103578 -3274 104166 -3219
rect 106860 -3232 106870 -3219
rect 103450 -3277 104166 -3274
rect 100364 -3393 100564 -3385
rect 100380 -3397 100548 -3393
rect 96962 -3628 96964 -3574
rect 100106 -3600 100280 -3514
rect 100306 -3574 100406 -3450
rect 103450 -3514 103594 -3277
rect 103780 -3299 104166 -3277
rect 103704 -3385 104166 -3299
rect 106794 -3274 106870 -3232
rect 103708 -3393 103908 -3385
rect 103724 -3397 103892 -3393
rect 100306 -3628 100308 -3574
rect 103450 -3600 103624 -3514
rect 103650 -3574 103750 -3450
rect 106794 -3514 106938 -3274
rect 103650 -3628 103652 -3574
rect 106794 -3600 106968 -3514
rect 106994 -3574 107094 -3450
rect 106994 -3628 106996 -3574
rect 3015 -4371 3159 -4324
rect 3196 -4371 3213 -4270
rect 6359 -4371 6503 -4324
rect 6540 -4371 6557 -4270
rect 9703 -4371 9847 -4324
rect 9884 -4371 9901 -4270
rect 13047 -4371 13191 -4324
rect 13228 -4371 13245 -4270
rect 16391 -4371 16535 -4324
rect 16572 -4371 16589 -4270
rect 19735 -4371 19879 -4324
rect 19916 -4371 19933 -4270
rect 23079 -4371 23223 -4324
rect 23260 -4371 23277 -4270
rect 26423 -4371 26567 -4324
rect 26604 -4371 26621 -4270
rect 29767 -4371 29911 -4324
rect 29948 -4371 29965 -4270
rect 33111 -4371 33255 -4324
rect 33292 -4371 33309 -4270
rect 36455 -4371 36599 -4324
rect 36636 -4371 36653 -4270
rect 39799 -4371 39943 -4324
rect 39980 -4371 39997 -4270
rect 43143 -4371 43287 -4324
rect 43324 -4371 43341 -4270
rect 46487 -4371 46631 -4324
rect 46668 -4371 46685 -4270
rect 49831 -4371 49975 -4324
rect 50012 -4371 50029 -4270
rect 56519 -4371 56663 -4324
rect 56700 -4371 56717 -4270
rect 59863 -4371 60007 -4324
rect 60044 -4371 60061 -4270
rect 63207 -4371 63351 -4324
rect 63388 -4371 63405 -4270
rect 66551 -4371 66695 -4324
rect 66732 -4371 66749 -4270
rect 69895 -4371 70039 -4324
rect 70076 -4371 70093 -4270
rect 73239 -4371 73383 -4324
rect 73420 -4371 73437 -4270
rect 76583 -4371 76727 -4324
rect 76764 -4371 76781 -4270
rect 79927 -4371 80071 -4324
rect 80108 -4371 80125 -4270
rect 83271 -4371 83415 -4324
rect 83452 -4371 83469 -4270
rect 86615 -4371 86759 -4324
rect 86796 -4371 86813 -4270
rect 89959 -4371 90103 -4324
rect 90140 -4371 90157 -4270
rect 93303 -4371 93447 -4324
rect 93484 -4371 93501 -4270
rect 96647 -4371 96791 -4324
rect 96828 -4371 96845 -4270
rect 99991 -4371 100135 -4324
rect 100172 -4371 100189 -4270
rect 103335 -4371 103479 -4324
rect 103516 -4371 103533 -4270
rect 106679 -4371 106823 -4324
rect 106860 -4371 106877 -4270
rect 3015 -4382 3787 -4371
rect 6359 -4382 7131 -4371
rect 9703 -4382 10475 -4371
rect 13047 -4382 13819 -4371
rect 16391 -4382 17163 -4371
rect 19735 -4382 20507 -4371
rect 23079 -4382 23851 -4371
rect 26423 -4382 27195 -4371
rect 29767 -4382 30539 -4371
rect 33111 -4382 33883 -4371
rect 36455 -4382 37227 -4371
rect 39799 -4382 40571 -4371
rect 43143 -4382 43915 -4371
rect 46487 -4382 47259 -4371
rect 49831 -4382 50603 -4371
rect 56519 -4382 56635 -4371
rect 3101 -4407 3787 -4382
rect 6445 -4407 7131 -4382
rect 9789 -4407 10475 -4382
rect 13133 -4407 13819 -4382
rect 16477 -4407 17163 -4382
rect 19821 -4407 20507 -4382
rect 23165 -4407 23851 -4382
rect 26509 -4407 27195 -4382
rect 29853 -4407 30539 -4382
rect 33197 -4407 33883 -4382
rect 36541 -4407 37227 -4382
rect 39885 -4407 40571 -4382
rect 43229 -4407 43915 -4382
rect 46573 -4407 47259 -4382
rect 49917 -4407 50603 -4382
rect 56605 -4407 56635 -4382
rect 3113 -4436 3787 -4407
rect 6457 -4436 7131 -4407
rect 9801 -4436 10475 -4407
rect 13145 -4436 13819 -4407
rect 16489 -4436 17163 -4407
rect 19833 -4436 20507 -4407
rect 23177 -4436 23851 -4407
rect 26521 -4436 27195 -4407
rect 29865 -4436 30539 -4407
rect 33209 -4436 33883 -4407
rect 36553 -4436 37227 -4407
rect 39897 -4436 40571 -4407
rect 43241 -4436 43915 -4407
rect 46585 -4436 47259 -4407
rect 49929 -4436 50603 -4407
rect 3113 -4848 3846 -4436
rect 4295 -4848 4342 -4483
rect 4349 -4848 4396 -4537
rect 6457 -4848 7190 -4436
rect 7639 -4848 7686 -4483
rect 7693 -4848 7740 -4537
rect 9801 -4848 10534 -4436
rect 10983 -4848 11030 -4483
rect 11037 -4848 11084 -4537
rect 13145 -4848 13878 -4436
rect 14327 -4848 14374 -4483
rect 14381 -4848 14428 -4537
rect 16489 -4848 17222 -4436
rect 17671 -4848 17718 -4483
rect 17725 -4848 17772 -4537
rect 19833 -4848 20566 -4436
rect 21015 -4848 21062 -4483
rect 21069 -4848 21116 -4537
rect 23177 -4848 23910 -4436
rect 24359 -4848 24406 -4483
rect 24413 -4848 24460 -4537
rect 26521 -4848 27254 -4436
rect 27703 -4848 27750 -4483
rect 27757 -4848 27804 -4537
rect 29865 -4848 30598 -4436
rect 31047 -4848 31094 -4483
rect 31101 -4848 31148 -4537
rect 33209 -4848 33942 -4436
rect 34391 -4848 34438 -4483
rect 34445 -4848 34492 -4537
rect 36553 -4848 37286 -4436
rect 37735 -4848 37782 -4483
rect 37789 -4848 37836 -4537
rect 39897 -4848 40630 -4436
rect 41079 -4848 41126 -4483
rect 41133 -4848 41180 -4537
rect 43241 -4848 43974 -4436
rect 44423 -4848 44470 -4483
rect 44477 -4848 44524 -4537
rect 46585 -4848 47318 -4436
rect 47767 -4848 47814 -4483
rect 47821 -4848 47868 -4537
rect 49929 -4848 50662 -4436
rect 51111 -4848 51158 -4483
rect 51165 -4848 51212 -4537
rect 3113 -4906 4467 -4848
rect 6457 -4906 7811 -4848
rect 9801 -4906 11155 -4848
rect 13145 -4906 14499 -4848
rect 16489 -4906 17843 -4848
rect 19833 -4906 21187 -4848
rect 23177 -4906 24531 -4848
rect 26521 -4906 27875 -4848
rect 29865 -4906 31219 -4848
rect 33209 -4906 34563 -4848
rect 36553 -4906 37907 -4848
rect 39897 -4906 41251 -4848
rect 43241 -4906 44595 -4848
rect 46585 -4906 47939 -4848
rect 49929 -4906 50984 -4848
rect 2720 -4943 4467 -4906
rect 5884 -4943 7811 -4906
rect 9228 -4943 11155 -4906
rect 12572 -4943 14499 -4906
rect 15916 -4943 17843 -4906
rect 19260 -4943 21187 -4906
rect 22604 -4943 24531 -4906
rect 25948 -4943 27875 -4906
rect 29292 -4943 31219 -4906
rect 32636 -4943 34563 -4906
rect 35980 -4943 37907 -4906
rect 39324 -4943 41251 -4906
rect 42668 -4943 44595 -4906
rect 46012 -4943 47939 -4906
rect 2720 -5067 4969 -4943
rect 5884 -5067 8313 -4943
rect 9228 -5067 11657 -4943
rect 12572 -5067 15001 -4943
rect 15916 -5067 18345 -4943
rect 19260 -5067 21689 -4943
rect 22604 -5067 25033 -4943
rect 25948 -5067 28377 -4943
rect 29292 -5067 31721 -4943
rect 32636 -5067 35065 -4943
rect 35980 -5067 38409 -4943
rect 39324 -5067 41753 -4943
rect 42668 -5067 45097 -4943
rect 46012 -5067 48441 -4943
rect 2720 -6022 5022 -5067
rect 5884 -6022 8366 -5067
rect 9228 -6022 11710 -5067
rect 12572 -6022 15054 -5067
rect 15916 -6022 18398 -5067
rect 19260 -6022 21742 -5067
rect 22604 -6022 25086 -5067
rect 25948 -6022 28430 -5067
rect 29292 -6022 31774 -5067
rect 32636 -6022 35118 -5067
rect 35980 -6022 38462 -5067
rect 39324 -6022 41806 -5067
rect 42668 -6022 45150 -5067
rect 46012 -6022 48494 -5067
rect 49356 -6022 50984 -4906
rect 56617 -4906 56635 -4407
rect 59863 -4382 60635 -4371
rect 63207 -4382 63979 -4371
rect 66551 -4382 67323 -4371
rect 69895 -4382 70667 -4371
rect 73239 -4382 74011 -4371
rect 76583 -4382 77355 -4371
rect 79927 -4382 80699 -4371
rect 83271 -4382 84043 -4371
rect 86615 -4382 87387 -4371
rect 89959 -4382 90731 -4371
rect 93303 -4382 94075 -4371
rect 96647 -4382 97419 -4371
rect 99991 -4382 100763 -4371
rect 103335 -4382 104107 -4371
rect 106679 -4382 107451 -4371
rect 59949 -4407 60635 -4382
rect 63293 -4407 63979 -4382
rect 66637 -4407 67323 -4382
rect 69981 -4407 70667 -4382
rect 73325 -4407 74011 -4382
rect 76669 -4407 77355 -4382
rect 80013 -4407 80699 -4382
rect 83357 -4407 84043 -4382
rect 86701 -4407 87387 -4382
rect 90045 -4407 90731 -4382
rect 93389 -4407 94075 -4382
rect 96733 -4407 97419 -4382
rect 100077 -4407 100763 -4382
rect 103421 -4407 104107 -4382
rect 106765 -4407 107451 -4382
rect 59961 -4436 60635 -4407
rect 63305 -4436 63979 -4407
rect 66649 -4436 67323 -4407
rect 69993 -4436 70667 -4407
rect 73337 -4436 74011 -4407
rect 76681 -4436 77355 -4407
rect 80025 -4436 80699 -4407
rect 83369 -4436 84043 -4407
rect 86713 -4436 87387 -4407
rect 90057 -4436 90731 -4407
rect 93401 -4436 94075 -4407
rect 96745 -4436 97419 -4407
rect 100089 -4436 100763 -4407
rect 103433 -4436 104107 -4407
rect 106777 -4436 107451 -4407
rect 57799 -4848 57846 -4483
rect 57853 -4848 57900 -4537
rect 59961 -4848 60694 -4436
rect 61143 -4848 61190 -4483
rect 61197 -4848 61244 -4537
rect 63305 -4848 64038 -4436
rect 64487 -4848 64534 -4483
rect 64541 -4848 64588 -4537
rect 66649 -4848 67382 -4436
rect 67831 -4848 67878 -4483
rect 67885 -4848 67932 -4537
rect 69993 -4848 70726 -4436
rect 71175 -4848 71222 -4483
rect 71229 -4848 71276 -4537
rect 73337 -4848 74070 -4436
rect 74519 -4848 74566 -4483
rect 74573 -4848 74620 -4537
rect 76681 -4848 77414 -4436
rect 77863 -4848 77910 -4483
rect 77917 -4848 77964 -4537
rect 80025 -4848 80758 -4436
rect 81207 -4848 81254 -4483
rect 81261 -4848 81308 -4537
rect 83369 -4848 84102 -4436
rect 84551 -4848 84598 -4483
rect 84605 -4848 84652 -4537
rect 86713 -4848 87446 -4436
rect 87895 -4848 87942 -4483
rect 87949 -4848 87996 -4537
rect 90057 -4848 90790 -4436
rect 91239 -4848 91286 -4483
rect 91293 -4848 91340 -4537
rect 93401 -4848 94134 -4436
rect 94583 -4848 94630 -4483
rect 94637 -4848 94684 -4537
rect 96745 -4848 97478 -4436
rect 97927 -4848 97974 -4483
rect 97981 -4848 98028 -4537
rect 100089 -4848 100822 -4436
rect 101271 -4848 101318 -4483
rect 101325 -4848 101372 -4537
rect 103433 -4848 104166 -4436
rect 104615 -4848 104662 -4483
rect 104669 -4848 104716 -4537
rect 106777 -4848 107510 -4436
rect 107959 -4848 108006 -4483
rect 108013 -4848 108060 -4537
rect 3131 -6087 5022 -6022
rect 6475 -6087 8366 -6022
rect 9819 -6087 11710 -6022
rect 13163 -6087 15054 -6022
rect 16507 -6087 18398 -6022
rect 19851 -6087 21742 -6022
rect 23195 -6087 25086 -6022
rect 26539 -6087 28430 -6022
rect 29883 -6087 31774 -6022
rect 33227 -6087 35118 -6022
rect 36571 -6087 38462 -6022
rect 39915 -6087 41806 -6022
rect 43259 -6087 45150 -6022
rect 46603 -6087 48494 -6022
rect 49947 -6087 50984 -6022
rect 3722 -6147 5022 -6087
rect 7066 -6147 8366 -6087
rect 10410 -6147 11710 -6087
rect 13754 -6147 15054 -6087
rect 17098 -6147 18398 -6087
rect 20442 -6147 21742 -6087
rect 23786 -6147 25086 -6087
rect 27130 -6147 28430 -6087
rect 30474 -6147 31774 -6087
rect 33818 -6147 35118 -6087
rect 37162 -6147 38462 -6087
rect 40506 -6147 41806 -6087
rect 43850 -6147 45150 -6087
rect 47194 -6147 48494 -6087
rect 50538 -6147 50984 -6087
rect 3751 -6152 5022 -6147
rect 7095 -6152 8366 -6147
rect 10439 -6152 11710 -6147
rect 13783 -6152 15054 -6147
rect 17127 -6152 18398 -6147
rect 20471 -6152 21742 -6147
rect 23815 -6152 25086 -6147
rect 27159 -6152 28430 -6147
rect 30503 -6152 31774 -6147
rect 33847 -6152 35118 -6147
rect 37191 -6152 38462 -6147
rect 40535 -6152 41806 -6147
rect 43879 -6152 45150 -6147
rect 47223 -6152 48494 -6147
rect 50567 -6152 50984 -6147
rect 3875 -6170 5022 -6152
rect 7219 -6170 8366 -6152
rect 10563 -6170 11710 -6152
rect 13907 -6170 15054 -6152
rect 17251 -6170 18398 -6152
rect 20595 -6170 21742 -6152
rect 23939 -6170 25086 -6152
rect 27283 -6170 28430 -6152
rect 30627 -6170 31774 -6152
rect 33971 -6170 35118 -6152
rect 37315 -6170 38462 -6152
rect 40659 -6170 41806 -6152
rect 44003 -6170 45150 -6152
rect 47347 -6170 48494 -6152
rect 50691 -6170 51129 -6152
rect 4313 -6181 5022 -6170
rect 7657 -6181 8366 -6170
rect 11001 -6181 11710 -6170
rect 14345 -6181 15054 -6170
rect 17689 -6181 18398 -6170
rect 21033 -6181 21742 -6170
rect 24377 -6181 25086 -6170
rect 27721 -6181 28430 -6170
rect 31065 -6181 31774 -6170
rect 34409 -6181 35118 -6170
rect 37753 -6181 38462 -6170
rect 41097 -6181 41806 -6170
rect 44441 -6181 45150 -6170
rect 47785 -6181 48494 -6170
rect 4313 -6217 4987 -6181
rect 7657 -6217 8331 -6181
rect 11001 -6217 11675 -6181
rect 14345 -6217 15019 -6181
rect 17689 -6217 18363 -6181
rect 21033 -6217 21707 -6181
rect 24377 -6217 25051 -6181
rect 27721 -6217 28395 -6181
rect 31065 -6217 31739 -6181
rect 34409 -6217 35083 -6181
rect 37753 -6217 38427 -6181
rect 41097 -6217 41771 -6181
rect 44441 -6217 45115 -6181
rect 47785 -6217 48459 -6181
rect 51785 -6181 51838 -5067
rect 57768 -4943 57971 -4848
rect 59961 -4906 61315 -4848
rect 63305 -4906 64659 -4848
rect 66649 -4906 68003 -4848
rect 69993 -4906 71347 -4848
rect 73337 -4906 74691 -4848
rect 76681 -4906 78035 -4848
rect 80025 -4906 81379 -4848
rect 83369 -4906 84723 -4848
rect 86713 -4906 88067 -4848
rect 90057 -4906 91411 -4848
rect 93401 -4906 94755 -4848
rect 96745 -4906 98099 -4848
rect 100089 -4906 101443 -4848
rect 103433 -4906 104787 -4848
rect 106777 -4906 108131 -4848
rect 59388 -4943 61315 -4906
rect 62732 -4943 64659 -4906
rect 66076 -4943 68003 -4906
rect 69420 -4943 71347 -4906
rect 72764 -4943 74691 -4906
rect 76108 -4943 78035 -4906
rect 79452 -4943 81379 -4906
rect 82796 -4943 84723 -4906
rect 86140 -4943 88067 -4906
rect 89484 -4943 91411 -4906
rect 92828 -4943 94755 -4906
rect 96172 -4943 98099 -4906
rect 99516 -4943 101443 -4906
rect 102860 -4943 104787 -4906
rect 106204 -4943 108131 -4906
rect 57768 -5067 58473 -4943
rect 59388 -5067 61817 -4943
rect 62732 -5067 65161 -4943
rect 66076 -5067 68505 -4943
rect 69420 -5067 71849 -4943
rect 72764 -5067 75193 -4943
rect 76108 -5067 78537 -4943
rect 79452 -5067 81881 -4943
rect 82796 -5067 85225 -4943
rect 86140 -5067 88569 -4943
rect 89484 -5067 91913 -4943
rect 92828 -5067 95257 -4943
rect 96172 -5067 98601 -4943
rect 99516 -5067 101945 -4943
rect 102860 -5067 105289 -4943
rect 106204 -5067 108633 -4943
rect 57768 -6152 58526 -5067
rect 59388 -6022 61870 -5067
rect 62732 -6022 65214 -5067
rect 66076 -6022 68558 -5067
rect 69420 -6022 71902 -5067
rect 72764 -6022 75246 -5067
rect 76108 -6022 78590 -5067
rect 79452 -6022 81934 -5067
rect 82796 -6022 85278 -5067
rect 86140 -6022 88622 -5067
rect 89484 -6022 91966 -5067
rect 92828 -6022 95310 -5067
rect 96172 -6022 98654 -5067
rect 99516 -6022 101998 -5067
rect 102860 -6022 105342 -5067
rect 106204 -6022 108686 -5067
rect 59979 -6087 61870 -6022
rect 63323 -6087 65214 -6022
rect 66667 -6087 68558 -6022
rect 70011 -6087 71902 -6022
rect 73355 -6087 75246 -6022
rect 76699 -6087 78590 -6022
rect 80043 -6087 81934 -6022
rect 83387 -6087 85278 -6022
rect 86731 -6087 88622 -6022
rect 90075 -6087 91966 -6022
rect 93419 -6087 95310 -6022
rect 96763 -6087 98654 -6022
rect 100107 -6087 101998 -6022
rect 103451 -6087 105342 -6022
rect 106795 -6087 108686 -6022
rect 60570 -6147 61870 -6087
rect 63914 -6147 65214 -6087
rect 67258 -6147 68558 -6087
rect 70602 -6147 71902 -6087
rect 73946 -6147 75246 -6087
rect 77290 -6147 78590 -6087
rect 80634 -6147 81934 -6087
rect 83978 -6147 85278 -6087
rect 87322 -6147 88622 -6087
rect 90666 -6147 91966 -6087
rect 94010 -6147 95310 -6087
rect 97354 -6147 98654 -6087
rect 100698 -6147 101998 -6087
rect 104042 -6147 105342 -6087
rect 107386 -6147 108686 -6087
rect 60599 -6152 61870 -6147
rect 63943 -6152 65214 -6147
rect 67287 -6152 68558 -6147
rect 70631 -6152 71902 -6147
rect 73975 -6152 75246 -6147
rect 77319 -6152 78590 -6147
rect 80663 -6152 81934 -6147
rect 84007 -6152 85278 -6147
rect 87351 -6152 88622 -6147
rect 90695 -6152 91966 -6147
rect 94039 -6152 95310 -6147
rect 97383 -6152 98654 -6147
rect 100727 -6152 101998 -6147
rect 104071 -6152 105342 -6147
rect 107415 -6152 108686 -6147
rect 57379 -6170 58526 -6152
rect 60723 -6170 61870 -6152
rect 64067 -6170 65214 -6152
rect 67411 -6170 68558 -6152
rect 70755 -6170 71902 -6152
rect 74099 -6170 75246 -6152
rect 77443 -6170 78590 -6152
rect 80787 -6170 81934 -6152
rect 84131 -6170 85278 -6152
rect 87475 -6170 88622 -6152
rect 90819 -6170 91966 -6152
rect 94163 -6170 95310 -6152
rect 97507 -6170 98654 -6152
rect 100851 -6170 101998 -6152
rect 104195 -6170 105342 -6152
rect 107539 -6170 108686 -6152
rect 57817 -6181 58526 -6170
rect 61161 -6181 61870 -6170
rect 64505 -6181 65214 -6170
rect 67849 -6181 68558 -6170
rect 71193 -6181 71902 -6170
rect 74537 -6181 75246 -6170
rect 77881 -6181 78590 -6170
rect 81225 -6181 81934 -6170
rect 84569 -6181 85278 -6170
rect 87913 -6181 88622 -6170
rect 91257 -6181 91966 -6170
rect 94601 -6181 95310 -6170
rect 97945 -6181 98654 -6170
rect 101289 -6181 101998 -6170
rect 104633 -6181 105342 -6170
rect 107977 -6181 108686 -6170
rect 51785 -6217 51803 -6181
rect 57817 -6217 58491 -6181
rect 61161 -6217 61835 -6181
rect 64505 -6217 65179 -6181
rect 67849 -6217 68523 -6181
rect 71193 -6217 71867 -6181
rect 74537 -6217 75211 -6181
rect 77881 -6217 78555 -6181
rect 81225 -6217 81899 -6181
rect 84569 -6217 85243 -6181
rect 87913 -6217 88587 -6181
rect 91257 -6217 91931 -6181
rect 94601 -6217 95275 -6181
rect 97945 -6217 98619 -6181
rect 101289 -6217 101963 -6181
rect 104633 -6217 105307 -6181
rect 107977 -6217 108651 -6181
rect 4496 -6235 4987 -6217
rect 7840 -6235 8331 -6217
rect 11184 -6235 11675 -6217
rect 14528 -6235 15019 -6217
rect 17872 -6235 18363 -6217
rect 21216 -6235 21707 -6217
rect 24560 -6235 25051 -6217
rect 27904 -6235 28395 -6217
rect 31248 -6235 31739 -6217
rect 34592 -6235 35083 -6217
rect 37936 -6235 38427 -6217
rect 41280 -6235 41771 -6217
rect 44624 -6235 45115 -6217
rect 47968 -6235 48459 -6217
rect 51312 -6235 51803 -6217
rect 58000 -6235 58491 -6217
rect 61344 -6235 61835 -6217
rect 64688 -6235 65179 -6217
rect 68032 -6235 68523 -6217
rect 71376 -6235 71867 -6217
rect 74720 -6235 75211 -6217
rect 78064 -6235 78555 -6217
rect 81408 -6235 81899 -6217
rect 84752 -6235 85243 -6217
rect 88096 -6235 88587 -6217
rect 91440 -6235 91931 -6217
rect 94784 -6235 95275 -6217
rect 98128 -6235 98619 -6217
rect 101472 -6235 101963 -6217
rect 104816 -6235 105307 -6217
rect 108160 -6235 108651 -6217
<< error_s >>
rect 53504 -2965 53620 -2899
rect 53620 -3219 54006 -3153
rect 53356 -3232 53366 -3219
rect 53290 -3274 53366 -3232
rect 53418 -3274 54006 -3219
rect 53290 -3277 54006 -3274
rect 53290 -3514 53434 -3277
rect 53620 -3299 54006 -3277
rect 53544 -3385 54006 -3299
rect 53548 -3393 53748 -3385
rect 53564 -3397 53732 -3393
rect 53290 -3600 53464 -3514
rect 53490 -3574 53590 -3450
rect 53490 -3628 53492 -3574
rect 53175 -4371 53319 -4324
rect 53356 -4371 53373 -4270
rect 53175 -4382 53947 -4371
rect 53261 -4407 53947 -4382
rect 53273 -4436 53947 -4407
rect 53273 -4848 54006 -4436
rect 54455 -4848 54502 -4483
rect 54509 -4848 54556 -4537
rect 53273 -4906 54627 -4848
rect 52700 -4943 54627 -4906
rect 52700 -5067 55129 -4943
rect 52700 -6022 55182 -5067
rect 56044 -6022 56508 -4906
rect 53291 -6087 55182 -6022
rect 53882 -6147 55182 -6087
rect 53911 -6152 55182 -6147
rect 54035 -6170 55182 -6152
rect 54473 -6181 55182 -6170
rect 54473 -6217 55147 -6181
rect 54656 -6235 55147 -6217
<< error_ps >>
rect 56634 -3514 56778 -3274
rect 56964 -3299 57350 -3153
rect 56888 -3385 57350 -3299
rect 56634 -3600 56808 -3514
rect 2540 -6022 2720 -4906
rect 50984 -4943 51283 -4848
rect 56635 -4436 57291 -4371
rect 56635 -4848 57350 -4436
rect 56635 -4906 57768 -4848
rect 50984 -6152 51785 -4943
rect 51129 -6217 51785 -6152
rect 56508 -6022 57768 -4906
rect 56635 -6087 57768 -6022
rect 57226 -6147 57768 -6087
rect 57255 -6152 57768 -6147
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
use icell16scs  x1
timestamp 1717439242
transform 1 0 0 0 1 0
box 0 -6337 55248 458
use icell16scs  x2
timestamp 1717439242
transform 1 0 53504 0 1 0
box 0 -6337 55248 458
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
