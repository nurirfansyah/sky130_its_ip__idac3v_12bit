magic
tech sky130A
magscale 1 2
timestamp 1717425130
<< viali >>
rect 2762 961 2796 995
rect 3051 856 3085 890
rect 2907 821 2941 855
rect 1237 -100 1271 2
rect 2912 -93 2946 -59
rect 4041 -192 4075 -158
<< metal1 >>
rect 722 1152 3602 1229
rect 722 1084 1153 1152
rect 1231 1084 3602 1152
rect 722 1081 3602 1084
rect 2749 995 3097 1007
rect 2749 961 2762 995
rect 2796 961 3097 995
rect 2749 949 3097 961
rect 3039 890 3097 949
rect 2891 865 2957 872
rect 2891 812 2897 865
rect 2951 812 2957 865
rect 3039 856 3051 890
rect 3085 856 3097 890
rect 3039 844 3097 856
rect 2891 806 2957 812
rect 3936 535 4136 676
rect 722 415 3602 517
rect 3936 483 4032 535
rect 4084 483 4136 535
rect 3936 476 4136 483
rect 722 403 4274 415
rect 722 334 1377 403
rect 1455 334 4274 403
rect 722 267 4274 334
rect 1667 231 1759 239
rect 1667 163 1675 231
rect 1753 163 1759 231
rect 1667 156 1759 163
rect 823 18 1023 84
rect 823 2 1283 18
rect 823 -100 1237 2
rect 1271 -100 1283 2
rect 823 -116 1283 -100
rect 2896 -49 2962 -43
rect 2896 -102 2902 -49
rect 2956 -102 2962 -49
rect 2896 -108 2962 -102
rect 4026 -149 4090 -143
rect 4026 -201 4032 -149
rect 4084 -201 4090 -149
rect 4026 -207 4090 -201
rect 722 -300 4274 -297
rect 722 -368 1153 -300
rect 1231 -368 4274 -300
rect 722 -445 4274 -368
rect 722 -514 4274 -473
rect 722 -672 1376 -514
rect 1456 -672 4274 -514
rect 722 -673 4274 -672
rect 722 -743 4274 -701
rect 722 -901 1673 -743
rect 1753 -901 4274 -743
rect 722 -1087 1152 -929
rect 1232 -1087 4274 -929
rect 722 -1129 4274 -1087
<< via1 >>
rect 1153 1084 1231 1152
rect 2897 855 2951 865
rect 2897 821 2907 855
rect 2907 821 2941 855
rect 2941 821 2951 855
rect 2897 812 2951 821
rect 4032 483 4084 535
rect 1377 334 1455 403
rect 1675 163 1753 231
rect 2902 -59 2956 -49
rect 2902 -93 2912 -59
rect 2912 -93 2946 -59
rect 2946 -93 2956 -59
rect 2902 -102 2956 -93
rect 4032 -158 4084 -149
rect 4032 -192 4041 -158
rect 4041 -192 4075 -158
rect 4075 -192 4084 -158
rect 4032 -201 4084 -192
rect 1153 -368 1231 -300
rect 1376 -672 1456 -514
rect 1673 -901 1753 -743
rect 1152 -1087 1232 -929
<< metal2 >>
rect 1146 1152 1238 1155
rect 1146 1084 1153 1152
rect 1231 1084 1238 1152
rect 1146 -300 1238 1084
rect 2889 865 2962 873
rect 2889 812 2897 865
rect 2951 812 2962 865
rect 1146 -368 1153 -300
rect 1231 -368 1238 -300
rect 1146 -929 1238 -368
rect 1370 403 1462 415
rect 1370 334 1377 403
rect 1455 334 1462 403
rect 1370 -514 1462 334
rect 1370 -672 1376 -514
rect 1456 -672 1462 -514
rect 1370 -676 1462 -672
rect 1667 231 1759 239
rect 1667 163 1675 231
rect 1753 163 1759 231
rect 1667 -743 1759 163
rect 2889 -49 2962 812
rect 2889 -102 2902 -49
rect 2956 -102 2962 -49
rect 2889 -108 2962 -102
rect 4026 535 4090 542
rect 4026 483 4032 535
rect 4084 483 4090 535
rect 4026 -149 4090 483
rect 4026 -201 4032 -149
rect 4084 -201 4090 -149
rect 4026 -207 4090 -201
rect 1667 -901 1673 -743
rect 1753 -901 1759 -743
rect 1667 -906 1759 -901
rect 1146 -1087 1152 -929
rect 1232 -1087 1238 -929
rect 1146 -1129 1238 -1087
use sky130_fd_sc_hvl__lsbuflv2hv_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1709947739
transform 1 0 722 0 1 -422
box -66 -43 2178 1671
use sky130_fd_sc_hvl__inv_4  x2 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1709947739
transform -1 0 3602 0 -1 1206
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_8  x3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1709947739
transform 1 0 2834 0 1 -422
box -66 -43 1506 897
<< labels >>
flabel metal1 s 722 -809 722 -809 3 FreeSans 800 0 0 0 dvdd
port 0 e
flabel metal1 s 722 -583 722 -583 3 FreeSans 800 0 0 0 avdd
port 1 e
flabel metal1 s 823 -7 823 -7 3 FreeSans 800 0 0 0 blv_in
port 2 e
flabel metal1 s 3935 573 3936 573 3 FreeSans 800 0 0 0 bhv_out
port 3 e
flabel metal1 s 722 -1028 722 -1028 3 FreeSans 800 0 0 0 dvss
port 4 e
<< end >>
