magic
tech sky130A
timestamp 1717438951
<< metal1 >>
rect 5878 -657 6339 -557
use icell2scs  x1
timestamp 1717438951
transform 1 0 0 0 1 0
box 2431 -2580 6083 1395
use icell2scs  x2
timestamp 1717438951
transform 1 0 3630 0 1 0
box 2431 -2580 6083 1395
<< end >>
