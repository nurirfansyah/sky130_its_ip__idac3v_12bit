magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< pwell >>
rect -328 -181653 328 181653
<< mvnmos >>
rect -100 180195 100 181395
rect -100 178777 100 179977
rect -100 177359 100 178559
rect -100 175941 100 177141
rect -100 174523 100 175723
rect -100 173105 100 174305
rect -100 171687 100 172887
rect -100 170269 100 171469
rect -100 168851 100 170051
rect -100 167433 100 168633
rect -100 166015 100 167215
rect -100 164597 100 165797
rect -100 163179 100 164379
rect -100 161761 100 162961
rect -100 160343 100 161543
rect -100 158925 100 160125
rect -100 157507 100 158707
rect -100 156089 100 157289
rect -100 154671 100 155871
rect -100 153253 100 154453
rect -100 151835 100 153035
rect -100 150417 100 151617
rect -100 148999 100 150199
rect -100 147581 100 148781
rect -100 146163 100 147363
rect -100 144745 100 145945
rect -100 143327 100 144527
rect -100 141909 100 143109
rect -100 140491 100 141691
rect -100 139073 100 140273
rect -100 137655 100 138855
rect -100 136237 100 137437
rect -100 134819 100 136019
rect -100 133401 100 134601
rect -100 131983 100 133183
rect -100 130565 100 131765
rect -100 129147 100 130347
rect -100 127729 100 128929
rect -100 126311 100 127511
rect -100 124893 100 126093
rect -100 123475 100 124675
rect -100 122057 100 123257
rect -100 120639 100 121839
rect -100 119221 100 120421
rect -100 117803 100 119003
rect -100 116385 100 117585
rect -100 114967 100 116167
rect -100 113549 100 114749
rect -100 112131 100 113331
rect -100 110713 100 111913
rect -100 109295 100 110495
rect -100 107877 100 109077
rect -100 106459 100 107659
rect -100 105041 100 106241
rect -100 103623 100 104823
rect -100 102205 100 103405
rect -100 100787 100 101987
rect -100 99369 100 100569
rect -100 97951 100 99151
rect -100 96533 100 97733
rect -100 95115 100 96315
rect -100 93697 100 94897
rect -100 92279 100 93479
rect -100 90861 100 92061
rect -100 89443 100 90643
rect -100 88025 100 89225
rect -100 86607 100 87807
rect -100 85189 100 86389
rect -100 83771 100 84971
rect -100 82353 100 83553
rect -100 80935 100 82135
rect -100 79517 100 80717
rect -100 78099 100 79299
rect -100 76681 100 77881
rect -100 75263 100 76463
rect -100 73845 100 75045
rect -100 72427 100 73627
rect -100 71009 100 72209
rect -100 69591 100 70791
rect -100 68173 100 69373
rect -100 66755 100 67955
rect -100 65337 100 66537
rect -100 63919 100 65119
rect -100 62501 100 63701
rect -100 61083 100 62283
rect -100 59665 100 60865
rect -100 58247 100 59447
rect -100 56829 100 58029
rect -100 55411 100 56611
rect -100 53993 100 55193
rect -100 52575 100 53775
rect -100 51157 100 52357
rect -100 49739 100 50939
rect -100 48321 100 49521
rect -100 46903 100 48103
rect -100 45485 100 46685
rect -100 44067 100 45267
rect -100 42649 100 43849
rect -100 41231 100 42431
rect -100 39813 100 41013
rect -100 38395 100 39595
rect -100 36977 100 38177
rect -100 35559 100 36759
rect -100 34141 100 35341
rect -100 32723 100 33923
rect -100 31305 100 32505
rect -100 29887 100 31087
rect -100 28469 100 29669
rect -100 27051 100 28251
rect -100 25633 100 26833
rect -100 24215 100 25415
rect -100 22797 100 23997
rect -100 21379 100 22579
rect -100 19961 100 21161
rect -100 18543 100 19743
rect -100 17125 100 18325
rect -100 15707 100 16907
rect -100 14289 100 15489
rect -100 12871 100 14071
rect -100 11453 100 12653
rect -100 10035 100 11235
rect -100 8617 100 9817
rect -100 7199 100 8399
rect -100 5781 100 6981
rect -100 4363 100 5563
rect -100 2945 100 4145
rect -100 1527 100 2727
rect -100 109 100 1309
rect -100 -1309 100 -109
rect -100 -2727 100 -1527
rect -100 -4145 100 -2945
rect -100 -5563 100 -4363
rect -100 -6981 100 -5781
rect -100 -8399 100 -7199
rect -100 -9817 100 -8617
rect -100 -11235 100 -10035
rect -100 -12653 100 -11453
rect -100 -14071 100 -12871
rect -100 -15489 100 -14289
rect -100 -16907 100 -15707
rect -100 -18325 100 -17125
rect -100 -19743 100 -18543
rect -100 -21161 100 -19961
rect -100 -22579 100 -21379
rect -100 -23997 100 -22797
rect -100 -25415 100 -24215
rect -100 -26833 100 -25633
rect -100 -28251 100 -27051
rect -100 -29669 100 -28469
rect -100 -31087 100 -29887
rect -100 -32505 100 -31305
rect -100 -33923 100 -32723
rect -100 -35341 100 -34141
rect -100 -36759 100 -35559
rect -100 -38177 100 -36977
rect -100 -39595 100 -38395
rect -100 -41013 100 -39813
rect -100 -42431 100 -41231
rect -100 -43849 100 -42649
rect -100 -45267 100 -44067
rect -100 -46685 100 -45485
rect -100 -48103 100 -46903
rect -100 -49521 100 -48321
rect -100 -50939 100 -49739
rect -100 -52357 100 -51157
rect -100 -53775 100 -52575
rect -100 -55193 100 -53993
rect -100 -56611 100 -55411
rect -100 -58029 100 -56829
rect -100 -59447 100 -58247
rect -100 -60865 100 -59665
rect -100 -62283 100 -61083
rect -100 -63701 100 -62501
rect -100 -65119 100 -63919
rect -100 -66537 100 -65337
rect -100 -67955 100 -66755
rect -100 -69373 100 -68173
rect -100 -70791 100 -69591
rect -100 -72209 100 -71009
rect -100 -73627 100 -72427
rect -100 -75045 100 -73845
rect -100 -76463 100 -75263
rect -100 -77881 100 -76681
rect -100 -79299 100 -78099
rect -100 -80717 100 -79517
rect -100 -82135 100 -80935
rect -100 -83553 100 -82353
rect -100 -84971 100 -83771
rect -100 -86389 100 -85189
rect -100 -87807 100 -86607
rect -100 -89225 100 -88025
rect -100 -90643 100 -89443
rect -100 -92061 100 -90861
rect -100 -93479 100 -92279
rect -100 -94897 100 -93697
rect -100 -96315 100 -95115
rect -100 -97733 100 -96533
rect -100 -99151 100 -97951
rect -100 -100569 100 -99369
rect -100 -101987 100 -100787
rect -100 -103405 100 -102205
rect -100 -104823 100 -103623
rect -100 -106241 100 -105041
rect -100 -107659 100 -106459
rect -100 -109077 100 -107877
rect -100 -110495 100 -109295
rect -100 -111913 100 -110713
rect -100 -113331 100 -112131
rect -100 -114749 100 -113549
rect -100 -116167 100 -114967
rect -100 -117585 100 -116385
rect -100 -119003 100 -117803
rect -100 -120421 100 -119221
rect -100 -121839 100 -120639
rect -100 -123257 100 -122057
rect -100 -124675 100 -123475
rect -100 -126093 100 -124893
rect -100 -127511 100 -126311
rect -100 -128929 100 -127729
rect -100 -130347 100 -129147
rect -100 -131765 100 -130565
rect -100 -133183 100 -131983
rect -100 -134601 100 -133401
rect -100 -136019 100 -134819
rect -100 -137437 100 -136237
rect -100 -138855 100 -137655
rect -100 -140273 100 -139073
rect -100 -141691 100 -140491
rect -100 -143109 100 -141909
rect -100 -144527 100 -143327
rect -100 -145945 100 -144745
rect -100 -147363 100 -146163
rect -100 -148781 100 -147581
rect -100 -150199 100 -148999
rect -100 -151617 100 -150417
rect -100 -153035 100 -151835
rect -100 -154453 100 -153253
rect -100 -155871 100 -154671
rect -100 -157289 100 -156089
rect -100 -158707 100 -157507
rect -100 -160125 100 -158925
rect -100 -161543 100 -160343
rect -100 -162961 100 -161761
rect -100 -164379 100 -163179
rect -100 -165797 100 -164597
rect -100 -167215 100 -166015
rect -100 -168633 100 -167433
rect -100 -170051 100 -168851
rect -100 -171469 100 -170269
rect -100 -172887 100 -171687
rect -100 -174305 100 -173105
rect -100 -175723 100 -174523
rect -100 -177141 100 -175941
rect -100 -178559 100 -177359
rect -100 -179977 100 -178777
rect -100 -181395 100 -180195
<< mvndiff >>
rect -158 181383 -100 181395
rect -158 180207 -146 181383
rect -112 180207 -100 181383
rect -158 180195 -100 180207
rect 100 181383 158 181395
rect 100 180207 112 181383
rect 146 180207 158 181383
rect 100 180195 158 180207
rect -158 179965 -100 179977
rect -158 178789 -146 179965
rect -112 178789 -100 179965
rect -158 178777 -100 178789
rect 100 179965 158 179977
rect 100 178789 112 179965
rect 146 178789 158 179965
rect 100 178777 158 178789
rect -158 178547 -100 178559
rect -158 177371 -146 178547
rect -112 177371 -100 178547
rect -158 177359 -100 177371
rect 100 178547 158 178559
rect 100 177371 112 178547
rect 146 177371 158 178547
rect 100 177359 158 177371
rect -158 177129 -100 177141
rect -158 175953 -146 177129
rect -112 175953 -100 177129
rect -158 175941 -100 175953
rect 100 177129 158 177141
rect 100 175953 112 177129
rect 146 175953 158 177129
rect 100 175941 158 175953
rect -158 175711 -100 175723
rect -158 174535 -146 175711
rect -112 174535 -100 175711
rect -158 174523 -100 174535
rect 100 175711 158 175723
rect 100 174535 112 175711
rect 146 174535 158 175711
rect 100 174523 158 174535
rect -158 174293 -100 174305
rect -158 173117 -146 174293
rect -112 173117 -100 174293
rect -158 173105 -100 173117
rect 100 174293 158 174305
rect 100 173117 112 174293
rect 146 173117 158 174293
rect 100 173105 158 173117
rect -158 172875 -100 172887
rect -158 171699 -146 172875
rect -112 171699 -100 172875
rect -158 171687 -100 171699
rect 100 172875 158 172887
rect 100 171699 112 172875
rect 146 171699 158 172875
rect 100 171687 158 171699
rect -158 171457 -100 171469
rect -158 170281 -146 171457
rect -112 170281 -100 171457
rect -158 170269 -100 170281
rect 100 171457 158 171469
rect 100 170281 112 171457
rect 146 170281 158 171457
rect 100 170269 158 170281
rect -158 170039 -100 170051
rect -158 168863 -146 170039
rect -112 168863 -100 170039
rect -158 168851 -100 168863
rect 100 170039 158 170051
rect 100 168863 112 170039
rect 146 168863 158 170039
rect 100 168851 158 168863
rect -158 168621 -100 168633
rect -158 167445 -146 168621
rect -112 167445 -100 168621
rect -158 167433 -100 167445
rect 100 168621 158 168633
rect 100 167445 112 168621
rect 146 167445 158 168621
rect 100 167433 158 167445
rect -158 167203 -100 167215
rect -158 166027 -146 167203
rect -112 166027 -100 167203
rect -158 166015 -100 166027
rect 100 167203 158 167215
rect 100 166027 112 167203
rect 146 166027 158 167203
rect 100 166015 158 166027
rect -158 165785 -100 165797
rect -158 164609 -146 165785
rect -112 164609 -100 165785
rect -158 164597 -100 164609
rect 100 165785 158 165797
rect 100 164609 112 165785
rect 146 164609 158 165785
rect 100 164597 158 164609
rect -158 164367 -100 164379
rect -158 163191 -146 164367
rect -112 163191 -100 164367
rect -158 163179 -100 163191
rect 100 164367 158 164379
rect 100 163191 112 164367
rect 146 163191 158 164367
rect 100 163179 158 163191
rect -158 162949 -100 162961
rect -158 161773 -146 162949
rect -112 161773 -100 162949
rect -158 161761 -100 161773
rect 100 162949 158 162961
rect 100 161773 112 162949
rect 146 161773 158 162949
rect 100 161761 158 161773
rect -158 161531 -100 161543
rect -158 160355 -146 161531
rect -112 160355 -100 161531
rect -158 160343 -100 160355
rect 100 161531 158 161543
rect 100 160355 112 161531
rect 146 160355 158 161531
rect 100 160343 158 160355
rect -158 160113 -100 160125
rect -158 158937 -146 160113
rect -112 158937 -100 160113
rect -158 158925 -100 158937
rect 100 160113 158 160125
rect 100 158937 112 160113
rect 146 158937 158 160113
rect 100 158925 158 158937
rect -158 158695 -100 158707
rect -158 157519 -146 158695
rect -112 157519 -100 158695
rect -158 157507 -100 157519
rect 100 158695 158 158707
rect 100 157519 112 158695
rect 146 157519 158 158695
rect 100 157507 158 157519
rect -158 157277 -100 157289
rect -158 156101 -146 157277
rect -112 156101 -100 157277
rect -158 156089 -100 156101
rect 100 157277 158 157289
rect 100 156101 112 157277
rect 146 156101 158 157277
rect 100 156089 158 156101
rect -158 155859 -100 155871
rect -158 154683 -146 155859
rect -112 154683 -100 155859
rect -158 154671 -100 154683
rect 100 155859 158 155871
rect 100 154683 112 155859
rect 146 154683 158 155859
rect 100 154671 158 154683
rect -158 154441 -100 154453
rect -158 153265 -146 154441
rect -112 153265 -100 154441
rect -158 153253 -100 153265
rect 100 154441 158 154453
rect 100 153265 112 154441
rect 146 153265 158 154441
rect 100 153253 158 153265
rect -158 153023 -100 153035
rect -158 151847 -146 153023
rect -112 151847 -100 153023
rect -158 151835 -100 151847
rect 100 153023 158 153035
rect 100 151847 112 153023
rect 146 151847 158 153023
rect 100 151835 158 151847
rect -158 151605 -100 151617
rect -158 150429 -146 151605
rect -112 150429 -100 151605
rect -158 150417 -100 150429
rect 100 151605 158 151617
rect 100 150429 112 151605
rect 146 150429 158 151605
rect 100 150417 158 150429
rect -158 150187 -100 150199
rect -158 149011 -146 150187
rect -112 149011 -100 150187
rect -158 148999 -100 149011
rect 100 150187 158 150199
rect 100 149011 112 150187
rect 146 149011 158 150187
rect 100 148999 158 149011
rect -158 148769 -100 148781
rect -158 147593 -146 148769
rect -112 147593 -100 148769
rect -158 147581 -100 147593
rect 100 148769 158 148781
rect 100 147593 112 148769
rect 146 147593 158 148769
rect 100 147581 158 147593
rect -158 147351 -100 147363
rect -158 146175 -146 147351
rect -112 146175 -100 147351
rect -158 146163 -100 146175
rect 100 147351 158 147363
rect 100 146175 112 147351
rect 146 146175 158 147351
rect 100 146163 158 146175
rect -158 145933 -100 145945
rect -158 144757 -146 145933
rect -112 144757 -100 145933
rect -158 144745 -100 144757
rect 100 145933 158 145945
rect 100 144757 112 145933
rect 146 144757 158 145933
rect 100 144745 158 144757
rect -158 144515 -100 144527
rect -158 143339 -146 144515
rect -112 143339 -100 144515
rect -158 143327 -100 143339
rect 100 144515 158 144527
rect 100 143339 112 144515
rect 146 143339 158 144515
rect 100 143327 158 143339
rect -158 143097 -100 143109
rect -158 141921 -146 143097
rect -112 141921 -100 143097
rect -158 141909 -100 141921
rect 100 143097 158 143109
rect 100 141921 112 143097
rect 146 141921 158 143097
rect 100 141909 158 141921
rect -158 141679 -100 141691
rect -158 140503 -146 141679
rect -112 140503 -100 141679
rect -158 140491 -100 140503
rect 100 141679 158 141691
rect 100 140503 112 141679
rect 146 140503 158 141679
rect 100 140491 158 140503
rect -158 140261 -100 140273
rect -158 139085 -146 140261
rect -112 139085 -100 140261
rect -158 139073 -100 139085
rect 100 140261 158 140273
rect 100 139085 112 140261
rect 146 139085 158 140261
rect 100 139073 158 139085
rect -158 138843 -100 138855
rect -158 137667 -146 138843
rect -112 137667 -100 138843
rect -158 137655 -100 137667
rect 100 138843 158 138855
rect 100 137667 112 138843
rect 146 137667 158 138843
rect 100 137655 158 137667
rect -158 137425 -100 137437
rect -158 136249 -146 137425
rect -112 136249 -100 137425
rect -158 136237 -100 136249
rect 100 137425 158 137437
rect 100 136249 112 137425
rect 146 136249 158 137425
rect 100 136237 158 136249
rect -158 136007 -100 136019
rect -158 134831 -146 136007
rect -112 134831 -100 136007
rect -158 134819 -100 134831
rect 100 136007 158 136019
rect 100 134831 112 136007
rect 146 134831 158 136007
rect 100 134819 158 134831
rect -158 134589 -100 134601
rect -158 133413 -146 134589
rect -112 133413 -100 134589
rect -158 133401 -100 133413
rect 100 134589 158 134601
rect 100 133413 112 134589
rect 146 133413 158 134589
rect 100 133401 158 133413
rect -158 133171 -100 133183
rect -158 131995 -146 133171
rect -112 131995 -100 133171
rect -158 131983 -100 131995
rect 100 133171 158 133183
rect 100 131995 112 133171
rect 146 131995 158 133171
rect 100 131983 158 131995
rect -158 131753 -100 131765
rect -158 130577 -146 131753
rect -112 130577 -100 131753
rect -158 130565 -100 130577
rect 100 131753 158 131765
rect 100 130577 112 131753
rect 146 130577 158 131753
rect 100 130565 158 130577
rect -158 130335 -100 130347
rect -158 129159 -146 130335
rect -112 129159 -100 130335
rect -158 129147 -100 129159
rect 100 130335 158 130347
rect 100 129159 112 130335
rect 146 129159 158 130335
rect 100 129147 158 129159
rect -158 128917 -100 128929
rect -158 127741 -146 128917
rect -112 127741 -100 128917
rect -158 127729 -100 127741
rect 100 128917 158 128929
rect 100 127741 112 128917
rect 146 127741 158 128917
rect 100 127729 158 127741
rect -158 127499 -100 127511
rect -158 126323 -146 127499
rect -112 126323 -100 127499
rect -158 126311 -100 126323
rect 100 127499 158 127511
rect 100 126323 112 127499
rect 146 126323 158 127499
rect 100 126311 158 126323
rect -158 126081 -100 126093
rect -158 124905 -146 126081
rect -112 124905 -100 126081
rect -158 124893 -100 124905
rect 100 126081 158 126093
rect 100 124905 112 126081
rect 146 124905 158 126081
rect 100 124893 158 124905
rect -158 124663 -100 124675
rect -158 123487 -146 124663
rect -112 123487 -100 124663
rect -158 123475 -100 123487
rect 100 124663 158 124675
rect 100 123487 112 124663
rect 146 123487 158 124663
rect 100 123475 158 123487
rect -158 123245 -100 123257
rect -158 122069 -146 123245
rect -112 122069 -100 123245
rect -158 122057 -100 122069
rect 100 123245 158 123257
rect 100 122069 112 123245
rect 146 122069 158 123245
rect 100 122057 158 122069
rect -158 121827 -100 121839
rect -158 120651 -146 121827
rect -112 120651 -100 121827
rect -158 120639 -100 120651
rect 100 121827 158 121839
rect 100 120651 112 121827
rect 146 120651 158 121827
rect 100 120639 158 120651
rect -158 120409 -100 120421
rect -158 119233 -146 120409
rect -112 119233 -100 120409
rect -158 119221 -100 119233
rect 100 120409 158 120421
rect 100 119233 112 120409
rect 146 119233 158 120409
rect 100 119221 158 119233
rect -158 118991 -100 119003
rect -158 117815 -146 118991
rect -112 117815 -100 118991
rect -158 117803 -100 117815
rect 100 118991 158 119003
rect 100 117815 112 118991
rect 146 117815 158 118991
rect 100 117803 158 117815
rect -158 117573 -100 117585
rect -158 116397 -146 117573
rect -112 116397 -100 117573
rect -158 116385 -100 116397
rect 100 117573 158 117585
rect 100 116397 112 117573
rect 146 116397 158 117573
rect 100 116385 158 116397
rect -158 116155 -100 116167
rect -158 114979 -146 116155
rect -112 114979 -100 116155
rect -158 114967 -100 114979
rect 100 116155 158 116167
rect 100 114979 112 116155
rect 146 114979 158 116155
rect 100 114967 158 114979
rect -158 114737 -100 114749
rect -158 113561 -146 114737
rect -112 113561 -100 114737
rect -158 113549 -100 113561
rect 100 114737 158 114749
rect 100 113561 112 114737
rect 146 113561 158 114737
rect 100 113549 158 113561
rect -158 113319 -100 113331
rect -158 112143 -146 113319
rect -112 112143 -100 113319
rect -158 112131 -100 112143
rect 100 113319 158 113331
rect 100 112143 112 113319
rect 146 112143 158 113319
rect 100 112131 158 112143
rect -158 111901 -100 111913
rect -158 110725 -146 111901
rect -112 110725 -100 111901
rect -158 110713 -100 110725
rect 100 111901 158 111913
rect 100 110725 112 111901
rect 146 110725 158 111901
rect 100 110713 158 110725
rect -158 110483 -100 110495
rect -158 109307 -146 110483
rect -112 109307 -100 110483
rect -158 109295 -100 109307
rect 100 110483 158 110495
rect 100 109307 112 110483
rect 146 109307 158 110483
rect 100 109295 158 109307
rect -158 109065 -100 109077
rect -158 107889 -146 109065
rect -112 107889 -100 109065
rect -158 107877 -100 107889
rect 100 109065 158 109077
rect 100 107889 112 109065
rect 146 107889 158 109065
rect 100 107877 158 107889
rect -158 107647 -100 107659
rect -158 106471 -146 107647
rect -112 106471 -100 107647
rect -158 106459 -100 106471
rect 100 107647 158 107659
rect 100 106471 112 107647
rect 146 106471 158 107647
rect 100 106459 158 106471
rect -158 106229 -100 106241
rect -158 105053 -146 106229
rect -112 105053 -100 106229
rect -158 105041 -100 105053
rect 100 106229 158 106241
rect 100 105053 112 106229
rect 146 105053 158 106229
rect 100 105041 158 105053
rect -158 104811 -100 104823
rect -158 103635 -146 104811
rect -112 103635 -100 104811
rect -158 103623 -100 103635
rect 100 104811 158 104823
rect 100 103635 112 104811
rect 146 103635 158 104811
rect 100 103623 158 103635
rect -158 103393 -100 103405
rect -158 102217 -146 103393
rect -112 102217 -100 103393
rect -158 102205 -100 102217
rect 100 103393 158 103405
rect 100 102217 112 103393
rect 146 102217 158 103393
rect 100 102205 158 102217
rect -158 101975 -100 101987
rect -158 100799 -146 101975
rect -112 100799 -100 101975
rect -158 100787 -100 100799
rect 100 101975 158 101987
rect 100 100799 112 101975
rect 146 100799 158 101975
rect 100 100787 158 100799
rect -158 100557 -100 100569
rect -158 99381 -146 100557
rect -112 99381 -100 100557
rect -158 99369 -100 99381
rect 100 100557 158 100569
rect 100 99381 112 100557
rect 146 99381 158 100557
rect 100 99369 158 99381
rect -158 99139 -100 99151
rect -158 97963 -146 99139
rect -112 97963 -100 99139
rect -158 97951 -100 97963
rect 100 99139 158 99151
rect 100 97963 112 99139
rect 146 97963 158 99139
rect 100 97951 158 97963
rect -158 97721 -100 97733
rect -158 96545 -146 97721
rect -112 96545 -100 97721
rect -158 96533 -100 96545
rect 100 97721 158 97733
rect 100 96545 112 97721
rect 146 96545 158 97721
rect 100 96533 158 96545
rect -158 96303 -100 96315
rect -158 95127 -146 96303
rect -112 95127 -100 96303
rect -158 95115 -100 95127
rect 100 96303 158 96315
rect 100 95127 112 96303
rect 146 95127 158 96303
rect 100 95115 158 95127
rect -158 94885 -100 94897
rect -158 93709 -146 94885
rect -112 93709 -100 94885
rect -158 93697 -100 93709
rect 100 94885 158 94897
rect 100 93709 112 94885
rect 146 93709 158 94885
rect 100 93697 158 93709
rect -158 93467 -100 93479
rect -158 92291 -146 93467
rect -112 92291 -100 93467
rect -158 92279 -100 92291
rect 100 93467 158 93479
rect 100 92291 112 93467
rect 146 92291 158 93467
rect 100 92279 158 92291
rect -158 92049 -100 92061
rect -158 90873 -146 92049
rect -112 90873 -100 92049
rect -158 90861 -100 90873
rect 100 92049 158 92061
rect 100 90873 112 92049
rect 146 90873 158 92049
rect 100 90861 158 90873
rect -158 90631 -100 90643
rect -158 89455 -146 90631
rect -112 89455 -100 90631
rect -158 89443 -100 89455
rect 100 90631 158 90643
rect 100 89455 112 90631
rect 146 89455 158 90631
rect 100 89443 158 89455
rect -158 89213 -100 89225
rect -158 88037 -146 89213
rect -112 88037 -100 89213
rect -158 88025 -100 88037
rect 100 89213 158 89225
rect 100 88037 112 89213
rect 146 88037 158 89213
rect 100 88025 158 88037
rect -158 87795 -100 87807
rect -158 86619 -146 87795
rect -112 86619 -100 87795
rect -158 86607 -100 86619
rect 100 87795 158 87807
rect 100 86619 112 87795
rect 146 86619 158 87795
rect 100 86607 158 86619
rect -158 86377 -100 86389
rect -158 85201 -146 86377
rect -112 85201 -100 86377
rect -158 85189 -100 85201
rect 100 86377 158 86389
rect 100 85201 112 86377
rect 146 85201 158 86377
rect 100 85189 158 85201
rect -158 84959 -100 84971
rect -158 83783 -146 84959
rect -112 83783 -100 84959
rect -158 83771 -100 83783
rect 100 84959 158 84971
rect 100 83783 112 84959
rect 146 83783 158 84959
rect 100 83771 158 83783
rect -158 83541 -100 83553
rect -158 82365 -146 83541
rect -112 82365 -100 83541
rect -158 82353 -100 82365
rect 100 83541 158 83553
rect 100 82365 112 83541
rect 146 82365 158 83541
rect 100 82353 158 82365
rect -158 82123 -100 82135
rect -158 80947 -146 82123
rect -112 80947 -100 82123
rect -158 80935 -100 80947
rect 100 82123 158 82135
rect 100 80947 112 82123
rect 146 80947 158 82123
rect 100 80935 158 80947
rect -158 80705 -100 80717
rect -158 79529 -146 80705
rect -112 79529 -100 80705
rect -158 79517 -100 79529
rect 100 80705 158 80717
rect 100 79529 112 80705
rect 146 79529 158 80705
rect 100 79517 158 79529
rect -158 79287 -100 79299
rect -158 78111 -146 79287
rect -112 78111 -100 79287
rect -158 78099 -100 78111
rect 100 79287 158 79299
rect 100 78111 112 79287
rect 146 78111 158 79287
rect 100 78099 158 78111
rect -158 77869 -100 77881
rect -158 76693 -146 77869
rect -112 76693 -100 77869
rect -158 76681 -100 76693
rect 100 77869 158 77881
rect 100 76693 112 77869
rect 146 76693 158 77869
rect 100 76681 158 76693
rect -158 76451 -100 76463
rect -158 75275 -146 76451
rect -112 75275 -100 76451
rect -158 75263 -100 75275
rect 100 76451 158 76463
rect 100 75275 112 76451
rect 146 75275 158 76451
rect 100 75263 158 75275
rect -158 75033 -100 75045
rect -158 73857 -146 75033
rect -112 73857 -100 75033
rect -158 73845 -100 73857
rect 100 75033 158 75045
rect 100 73857 112 75033
rect 146 73857 158 75033
rect 100 73845 158 73857
rect -158 73615 -100 73627
rect -158 72439 -146 73615
rect -112 72439 -100 73615
rect -158 72427 -100 72439
rect 100 73615 158 73627
rect 100 72439 112 73615
rect 146 72439 158 73615
rect 100 72427 158 72439
rect -158 72197 -100 72209
rect -158 71021 -146 72197
rect -112 71021 -100 72197
rect -158 71009 -100 71021
rect 100 72197 158 72209
rect 100 71021 112 72197
rect 146 71021 158 72197
rect 100 71009 158 71021
rect -158 70779 -100 70791
rect -158 69603 -146 70779
rect -112 69603 -100 70779
rect -158 69591 -100 69603
rect 100 70779 158 70791
rect 100 69603 112 70779
rect 146 69603 158 70779
rect 100 69591 158 69603
rect -158 69361 -100 69373
rect -158 68185 -146 69361
rect -112 68185 -100 69361
rect -158 68173 -100 68185
rect 100 69361 158 69373
rect 100 68185 112 69361
rect 146 68185 158 69361
rect 100 68173 158 68185
rect -158 67943 -100 67955
rect -158 66767 -146 67943
rect -112 66767 -100 67943
rect -158 66755 -100 66767
rect 100 67943 158 67955
rect 100 66767 112 67943
rect 146 66767 158 67943
rect 100 66755 158 66767
rect -158 66525 -100 66537
rect -158 65349 -146 66525
rect -112 65349 -100 66525
rect -158 65337 -100 65349
rect 100 66525 158 66537
rect 100 65349 112 66525
rect 146 65349 158 66525
rect 100 65337 158 65349
rect -158 65107 -100 65119
rect -158 63931 -146 65107
rect -112 63931 -100 65107
rect -158 63919 -100 63931
rect 100 65107 158 65119
rect 100 63931 112 65107
rect 146 63931 158 65107
rect 100 63919 158 63931
rect -158 63689 -100 63701
rect -158 62513 -146 63689
rect -112 62513 -100 63689
rect -158 62501 -100 62513
rect 100 63689 158 63701
rect 100 62513 112 63689
rect 146 62513 158 63689
rect 100 62501 158 62513
rect -158 62271 -100 62283
rect -158 61095 -146 62271
rect -112 61095 -100 62271
rect -158 61083 -100 61095
rect 100 62271 158 62283
rect 100 61095 112 62271
rect 146 61095 158 62271
rect 100 61083 158 61095
rect -158 60853 -100 60865
rect -158 59677 -146 60853
rect -112 59677 -100 60853
rect -158 59665 -100 59677
rect 100 60853 158 60865
rect 100 59677 112 60853
rect 146 59677 158 60853
rect 100 59665 158 59677
rect -158 59435 -100 59447
rect -158 58259 -146 59435
rect -112 58259 -100 59435
rect -158 58247 -100 58259
rect 100 59435 158 59447
rect 100 58259 112 59435
rect 146 58259 158 59435
rect 100 58247 158 58259
rect -158 58017 -100 58029
rect -158 56841 -146 58017
rect -112 56841 -100 58017
rect -158 56829 -100 56841
rect 100 58017 158 58029
rect 100 56841 112 58017
rect 146 56841 158 58017
rect 100 56829 158 56841
rect -158 56599 -100 56611
rect -158 55423 -146 56599
rect -112 55423 -100 56599
rect -158 55411 -100 55423
rect 100 56599 158 56611
rect 100 55423 112 56599
rect 146 55423 158 56599
rect 100 55411 158 55423
rect -158 55181 -100 55193
rect -158 54005 -146 55181
rect -112 54005 -100 55181
rect -158 53993 -100 54005
rect 100 55181 158 55193
rect 100 54005 112 55181
rect 146 54005 158 55181
rect 100 53993 158 54005
rect -158 53763 -100 53775
rect -158 52587 -146 53763
rect -112 52587 -100 53763
rect -158 52575 -100 52587
rect 100 53763 158 53775
rect 100 52587 112 53763
rect 146 52587 158 53763
rect 100 52575 158 52587
rect -158 52345 -100 52357
rect -158 51169 -146 52345
rect -112 51169 -100 52345
rect -158 51157 -100 51169
rect 100 52345 158 52357
rect 100 51169 112 52345
rect 146 51169 158 52345
rect 100 51157 158 51169
rect -158 50927 -100 50939
rect -158 49751 -146 50927
rect -112 49751 -100 50927
rect -158 49739 -100 49751
rect 100 50927 158 50939
rect 100 49751 112 50927
rect 146 49751 158 50927
rect 100 49739 158 49751
rect -158 49509 -100 49521
rect -158 48333 -146 49509
rect -112 48333 -100 49509
rect -158 48321 -100 48333
rect 100 49509 158 49521
rect 100 48333 112 49509
rect 146 48333 158 49509
rect 100 48321 158 48333
rect -158 48091 -100 48103
rect -158 46915 -146 48091
rect -112 46915 -100 48091
rect -158 46903 -100 46915
rect 100 48091 158 48103
rect 100 46915 112 48091
rect 146 46915 158 48091
rect 100 46903 158 46915
rect -158 46673 -100 46685
rect -158 45497 -146 46673
rect -112 45497 -100 46673
rect -158 45485 -100 45497
rect 100 46673 158 46685
rect 100 45497 112 46673
rect 146 45497 158 46673
rect 100 45485 158 45497
rect -158 45255 -100 45267
rect -158 44079 -146 45255
rect -112 44079 -100 45255
rect -158 44067 -100 44079
rect 100 45255 158 45267
rect 100 44079 112 45255
rect 146 44079 158 45255
rect 100 44067 158 44079
rect -158 43837 -100 43849
rect -158 42661 -146 43837
rect -112 42661 -100 43837
rect -158 42649 -100 42661
rect 100 43837 158 43849
rect 100 42661 112 43837
rect 146 42661 158 43837
rect 100 42649 158 42661
rect -158 42419 -100 42431
rect -158 41243 -146 42419
rect -112 41243 -100 42419
rect -158 41231 -100 41243
rect 100 42419 158 42431
rect 100 41243 112 42419
rect 146 41243 158 42419
rect 100 41231 158 41243
rect -158 41001 -100 41013
rect -158 39825 -146 41001
rect -112 39825 -100 41001
rect -158 39813 -100 39825
rect 100 41001 158 41013
rect 100 39825 112 41001
rect 146 39825 158 41001
rect 100 39813 158 39825
rect -158 39583 -100 39595
rect -158 38407 -146 39583
rect -112 38407 -100 39583
rect -158 38395 -100 38407
rect 100 39583 158 39595
rect 100 38407 112 39583
rect 146 38407 158 39583
rect 100 38395 158 38407
rect -158 38165 -100 38177
rect -158 36989 -146 38165
rect -112 36989 -100 38165
rect -158 36977 -100 36989
rect 100 38165 158 38177
rect 100 36989 112 38165
rect 146 36989 158 38165
rect 100 36977 158 36989
rect -158 36747 -100 36759
rect -158 35571 -146 36747
rect -112 35571 -100 36747
rect -158 35559 -100 35571
rect 100 36747 158 36759
rect 100 35571 112 36747
rect 146 35571 158 36747
rect 100 35559 158 35571
rect -158 35329 -100 35341
rect -158 34153 -146 35329
rect -112 34153 -100 35329
rect -158 34141 -100 34153
rect 100 35329 158 35341
rect 100 34153 112 35329
rect 146 34153 158 35329
rect 100 34141 158 34153
rect -158 33911 -100 33923
rect -158 32735 -146 33911
rect -112 32735 -100 33911
rect -158 32723 -100 32735
rect 100 33911 158 33923
rect 100 32735 112 33911
rect 146 32735 158 33911
rect 100 32723 158 32735
rect -158 32493 -100 32505
rect -158 31317 -146 32493
rect -112 31317 -100 32493
rect -158 31305 -100 31317
rect 100 32493 158 32505
rect 100 31317 112 32493
rect 146 31317 158 32493
rect 100 31305 158 31317
rect -158 31075 -100 31087
rect -158 29899 -146 31075
rect -112 29899 -100 31075
rect -158 29887 -100 29899
rect 100 31075 158 31087
rect 100 29899 112 31075
rect 146 29899 158 31075
rect 100 29887 158 29899
rect -158 29657 -100 29669
rect -158 28481 -146 29657
rect -112 28481 -100 29657
rect -158 28469 -100 28481
rect 100 29657 158 29669
rect 100 28481 112 29657
rect 146 28481 158 29657
rect 100 28469 158 28481
rect -158 28239 -100 28251
rect -158 27063 -146 28239
rect -112 27063 -100 28239
rect -158 27051 -100 27063
rect 100 28239 158 28251
rect 100 27063 112 28239
rect 146 27063 158 28239
rect 100 27051 158 27063
rect -158 26821 -100 26833
rect -158 25645 -146 26821
rect -112 25645 -100 26821
rect -158 25633 -100 25645
rect 100 26821 158 26833
rect 100 25645 112 26821
rect 146 25645 158 26821
rect 100 25633 158 25645
rect -158 25403 -100 25415
rect -158 24227 -146 25403
rect -112 24227 -100 25403
rect -158 24215 -100 24227
rect 100 25403 158 25415
rect 100 24227 112 25403
rect 146 24227 158 25403
rect 100 24215 158 24227
rect -158 23985 -100 23997
rect -158 22809 -146 23985
rect -112 22809 -100 23985
rect -158 22797 -100 22809
rect 100 23985 158 23997
rect 100 22809 112 23985
rect 146 22809 158 23985
rect 100 22797 158 22809
rect -158 22567 -100 22579
rect -158 21391 -146 22567
rect -112 21391 -100 22567
rect -158 21379 -100 21391
rect 100 22567 158 22579
rect 100 21391 112 22567
rect 146 21391 158 22567
rect 100 21379 158 21391
rect -158 21149 -100 21161
rect -158 19973 -146 21149
rect -112 19973 -100 21149
rect -158 19961 -100 19973
rect 100 21149 158 21161
rect 100 19973 112 21149
rect 146 19973 158 21149
rect 100 19961 158 19973
rect -158 19731 -100 19743
rect -158 18555 -146 19731
rect -112 18555 -100 19731
rect -158 18543 -100 18555
rect 100 19731 158 19743
rect 100 18555 112 19731
rect 146 18555 158 19731
rect 100 18543 158 18555
rect -158 18313 -100 18325
rect -158 17137 -146 18313
rect -112 17137 -100 18313
rect -158 17125 -100 17137
rect 100 18313 158 18325
rect 100 17137 112 18313
rect 146 17137 158 18313
rect 100 17125 158 17137
rect -158 16895 -100 16907
rect -158 15719 -146 16895
rect -112 15719 -100 16895
rect -158 15707 -100 15719
rect 100 16895 158 16907
rect 100 15719 112 16895
rect 146 15719 158 16895
rect 100 15707 158 15719
rect -158 15477 -100 15489
rect -158 14301 -146 15477
rect -112 14301 -100 15477
rect -158 14289 -100 14301
rect 100 15477 158 15489
rect 100 14301 112 15477
rect 146 14301 158 15477
rect 100 14289 158 14301
rect -158 14059 -100 14071
rect -158 12883 -146 14059
rect -112 12883 -100 14059
rect -158 12871 -100 12883
rect 100 14059 158 14071
rect 100 12883 112 14059
rect 146 12883 158 14059
rect 100 12871 158 12883
rect -158 12641 -100 12653
rect -158 11465 -146 12641
rect -112 11465 -100 12641
rect -158 11453 -100 11465
rect 100 12641 158 12653
rect 100 11465 112 12641
rect 146 11465 158 12641
rect 100 11453 158 11465
rect -158 11223 -100 11235
rect -158 10047 -146 11223
rect -112 10047 -100 11223
rect -158 10035 -100 10047
rect 100 11223 158 11235
rect 100 10047 112 11223
rect 146 10047 158 11223
rect 100 10035 158 10047
rect -158 9805 -100 9817
rect -158 8629 -146 9805
rect -112 8629 -100 9805
rect -158 8617 -100 8629
rect 100 9805 158 9817
rect 100 8629 112 9805
rect 146 8629 158 9805
rect 100 8617 158 8629
rect -158 8387 -100 8399
rect -158 7211 -146 8387
rect -112 7211 -100 8387
rect -158 7199 -100 7211
rect 100 8387 158 8399
rect 100 7211 112 8387
rect 146 7211 158 8387
rect 100 7199 158 7211
rect -158 6969 -100 6981
rect -158 5793 -146 6969
rect -112 5793 -100 6969
rect -158 5781 -100 5793
rect 100 6969 158 6981
rect 100 5793 112 6969
rect 146 5793 158 6969
rect 100 5781 158 5793
rect -158 5551 -100 5563
rect -158 4375 -146 5551
rect -112 4375 -100 5551
rect -158 4363 -100 4375
rect 100 5551 158 5563
rect 100 4375 112 5551
rect 146 4375 158 5551
rect 100 4363 158 4375
rect -158 4133 -100 4145
rect -158 2957 -146 4133
rect -112 2957 -100 4133
rect -158 2945 -100 2957
rect 100 4133 158 4145
rect 100 2957 112 4133
rect 146 2957 158 4133
rect 100 2945 158 2957
rect -158 2715 -100 2727
rect -158 1539 -146 2715
rect -112 1539 -100 2715
rect -158 1527 -100 1539
rect 100 2715 158 2727
rect 100 1539 112 2715
rect 146 1539 158 2715
rect 100 1527 158 1539
rect -158 1297 -100 1309
rect -158 121 -146 1297
rect -112 121 -100 1297
rect -158 109 -100 121
rect 100 1297 158 1309
rect 100 121 112 1297
rect 146 121 158 1297
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -1297 -146 -121
rect -112 -1297 -100 -121
rect -158 -1309 -100 -1297
rect 100 -121 158 -109
rect 100 -1297 112 -121
rect 146 -1297 158 -121
rect 100 -1309 158 -1297
rect -158 -1539 -100 -1527
rect -158 -2715 -146 -1539
rect -112 -2715 -100 -1539
rect -158 -2727 -100 -2715
rect 100 -1539 158 -1527
rect 100 -2715 112 -1539
rect 146 -2715 158 -1539
rect 100 -2727 158 -2715
rect -158 -2957 -100 -2945
rect -158 -4133 -146 -2957
rect -112 -4133 -100 -2957
rect -158 -4145 -100 -4133
rect 100 -2957 158 -2945
rect 100 -4133 112 -2957
rect 146 -4133 158 -2957
rect 100 -4145 158 -4133
rect -158 -4375 -100 -4363
rect -158 -5551 -146 -4375
rect -112 -5551 -100 -4375
rect -158 -5563 -100 -5551
rect 100 -4375 158 -4363
rect 100 -5551 112 -4375
rect 146 -5551 158 -4375
rect 100 -5563 158 -5551
rect -158 -5793 -100 -5781
rect -158 -6969 -146 -5793
rect -112 -6969 -100 -5793
rect -158 -6981 -100 -6969
rect 100 -5793 158 -5781
rect 100 -6969 112 -5793
rect 146 -6969 158 -5793
rect 100 -6981 158 -6969
rect -158 -7211 -100 -7199
rect -158 -8387 -146 -7211
rect -112 -8387 -100 -7211
rect -158 -8399 -100 -8387
rect 100 -7211 158 -7199
rect 100 -8387 112 -7211
rect 146 -8387 158 -7211
rect 100 -8399 158 -8387
rect -158 -8629 -100 -8617
rect -158 -9805 -146 -8629
rect -112 -9805 -100 -8629
rect -158 -9817 -100 -9805
rect 100 -8629 158 -8617
rect 100 -9805 112 -8629
rect 146 -9805 158 -8629
rect 100 -9817 158 -9805
rect -158 -10047 -100 -10035
rect -158 -11223 -146 -10047
rect -112 -11223 -100 -10047
rect -158 -11235 -100 -11223
rect 100 -10047 158 -10035
rect 100 -11223 112 -10047
rect 146 -11223 158 -10047
rect 100 -11235 158 -11223
rect -158 -11465 -100 -11453
rect -158 -12641 -146 -11465
rect -112 -12641 -100 -11465
rect -158 -12653 -100 -12641
rect 100 -11465 158 -11453
rect 100 -12641 112 -11465
rect 146 -12641 158 -11465
rect 100 -12653 158 -12641
rect -158 -12883 -100 -12871
rect -158 -14059 -146 -12883
rect -112 -14059 -100 -12883
rect -158 -14071 -100 -14059
rect 100 -12883 158 -12871
rect 100 -14059 112 -12883
rect 146 -14059 158 -12883
rect 100 -14071 158 -14059
rect -158 -14301 -100 -14289
rect -158 -15477 -146 -14301
rect -112 -15477 -100 -14301
rect -158 -15489 -100 -15477
rect 100 -14301 158 -14289
rect 100 -15477 112 -14301
rect 146 -15477 158 -14301
rect 100 -15489 158 -15477
rect -158 -15719 -100 -15707
rect -158 -16895 -146 -15719
rect -112 -16895 -100 -15719
rect -158 -16907 -100 -16895
rect 100 -15719 158 -15707
rect 100 -16895 112 -15719
rect 146 -16895 158 -15719
rect 100 -16907 158 -16895
rect -158 -17137 -100 -17125
rect -158 -18313 -146 -17137
rect -112 -18313 -100 -17137
rect -158 -18325 -100 -18313
rect 100 -17137 158 -17125
rect 100 -18313 112 -17137
rect 146 -18313 158 -17137
rect 100 -18325 158 -18313
rect -158 -18555 -100 -18543
rect -158 -19731 -146 -18555
rect -112 -19731 -100 -18555
rect -158 -19743 -100 -19731
rect 100 -18555 158 -18543
rect 100 -19731 112 -18555
rect 146 -19731 158 -18555
rect 100 -19743 158 -19731
rect -158 -19973 -100 -19961
rect -158 -21149 -146 -19973
rect -112 -21149 -100 -19973
rect -158 -21161 -100 -21149
rect 100 -19973 158 -19961
rect 100 -21149 112 -19973
rect 146 -21149 158 -19973
rect 100 -21161 158 -21149
rect -158 -21391 -100 -21379
rect -158 -22567 -146 -21391
rect -112 -22567 -100 -21391
rect -158 -22579 -100 -22567
rect 100 -21391 158 -21379
rect 100 -22567 112 -21391
rect 146 -22567 158 -21391
rect 100 -22579 158 -22567
rect -158 -22809 -100 -22797
rect -158 -23985 -146 -22809
rect -112 -23985 -100 -22809
rect -158 -23997 -100 -23985
rect 100 -22809 158 -22797
rect 100 -23985 112 -22809
rect 146 -23985 158 -22809
rect 100 -23997 158 -23985
rect -158 -24227 -100 -24215
rect -158 -25403 -146 -24227
rect -112 -25403 -100 -24227
rect -158 -25415 -100 -25403
rect 100 -24227 158 -24215
rect 100 -25403 112 -24227
rect 146 -25403 158 -24227
rect 100 -25415 158 -25403
rect -158 -25645 -100 -25633
rect -158 -26821 -146 -25645
rect -112 -26821 -100 -25645
rect -158 -26833 -100 -26821
rect 100 -25645 158 -25633
rect 100 -26821 112 -25645
rect 146 -26821 158 -25645
rect 100 -26833 158 -26821
rect -158 -27063 -100 -27051
rect -158 -28239 -146 -27063
rect -112 -28239 -100 -27063
rect -158 -28251 -100 -28239
rect 100 -27063 158 -27051
rect 100 -28239 112 -27063
rect 146 -28239 158 -27063
rect 100 -28251 158 -28239
rect -158 -28481 -100 -28469
rect -158 -29657 -146 -28481
rect -112 -29657 -100 -28481
rect -158 -29669 -100 -29657
rect 100 -28481 158 -28469
rect 100 -29657 112 -28481
rect 146 -29657 158 -28481
rect 100 -29669 158 -29657
rect -158 -29899 -100 -29887
rect -158 -31075 -146 -29899
rect -112 -31075 -100 -29899
rect -158 -31087 -100 -31075
rect 100 -29899 158 -29887
rect 100 -31075 112 -29899
rect 146 -31075 158 -29899
rect 100 -31087 158 -31075
rect -158 -31317 -100 -31305
rect -158 -32493 -146 -31317
rect -112 -32493 -100 -31317
rect -158 -32505 -100 -32493
rect 100 -31317 158 -31305
rect 100 -32493 112 -31317
rect 146 -32493 158 -31317
rect 100 -32505 158 -32493
rect -158 -32735 -100 -32723
rect -158 -33911 -146 -32735
rect -112 -33911 -100 -32735
rect -158 -33923 -100 -33911
rect 100 -32735 158 -32723
rect 100 -33911 112 -32735
rect 146 -33911 158 -32735
rect 100 -33923 158 -33911
rect -158 -34153 -100 -34141
rect -158 -35329 -146 -34153
rect -112 -35329 -100 -34153
rect -158 -35341 -100 -35329
rect 100 -34153 158 -34141
rect 100 -35329 112 -34153
rect 146 -35329 158 -34153
rect 100 -35341 158 -35329
rect -158 -35571 -100 -35559
rect -158 -36747 -146 -35571
rect -112 -36747 -100 -35571
rect -158 -36759 -100 -36747
rect 100 -35571 158 -35559
rect 100 -36747 112 -35571
rect 146 -36747 158 -35571
rect 100 -36759 158 -36747
rect -158 -36989 -100 -36977
rect -158 -38165 -146 -36989
rect -112 -38165 -100 -36989
rect -158 -38177 -100 -38165
rect 100 -36989 158 -36977
rect 100 -38165 112 -36989
rect 146 -38165 158 -36989
rect 100 -38177 158 -38165
rect -158 -38407 -100 -38395
rect -158 -39583 -146 -38407
rect -112 -39583 -100 -38407
rect -158 -39595 -100 -39583
rect 100 -38407 158 -38395
rect 100 -39583 112 -38407
rect 146 -39583 158 -38407
rect 100 -39595 158 -39583
rect -158 -39825 -100 -39813
rect -158 -41001 -146 -39825
rect -112 -41001 -100 -39825
rect -158 -41013 -100 -41001
rect 100 -39825 158 -39813
rect 100 -41001 112 -39825
rect 146 -41001 158 -39825
rect 100 -41013 158 -41001
rect -158 -41243 -100 -41231
rect -158 -42419 -146 -41243
rect -112 -42419 -100 -41243
rect -158 -42431 -100 -42419
rect 100 -41243 158 -41231
rect 100 -42419 112 -41243
rect 146 -42419 158 -41243
rect 100 -42431 158 -42419
rect -158 -42661 -100 -42649
rect -158 -43837 -146 -42661
rect -112 -43837 -100 -42661
rect -158 -43849 -100 -43837
rect 100 -42661 158 -42649
rect 100 -43837 112 -42661
rect 146 -43837 158 -42661
rect 100 -43849 158 -43837
rect -158 -44079 -100 -44067
rect -158 -45255 -146 -44079
rect -112 -45255 -100 -44079
rect -158 -45267 -100 -45255
rect 100 -44079 158 -44067
rect 100 -45255 112 -44079
rect 146 -45255 158 -44079
rect 100 -45267 158 -45255
rect -158 -45497 -100 -45485
rect -158 -46673 -146 -45497
rect -112 -46673 -100 -45497
rect -158 -46685 -100 -46673
rect 100 -45497 158 -45485
rect 100 -46673 112 -45497
rect 146 -46673 158 -45497
rect 100 -46685 158 -46673
rect -158 -46915 -100 -46903
rect -158 -48091 -146 -46915
rect -112 -48091 -100 -46915
rect -158 -48103 -100 -48091
rect 100 -46915 158 -46903
rect 100 -48091 112 -46915
rect 146 -48091 158 -46915
rect 100 -48103 158 -48091
rect -158 -48333 -100 -48321
rect -158 -49509 -146 -48333
rect -112 -49509 -100 -48333
rect -158 -49521 -100 -49509
rect 100 -48333 158 -48321
rect 100 -49509 112 -48333
rect 146 -49509 158 -48333
rect 100 -49521 158 -49509
rect -158 -49751 -100 -49739
rect -158 -50927 -146 -49751
rect -112 -50927 -100 -49751
rect -158 -50939 -100 -50927
rect 100 -49751 158 -49739
rect 100 -50927 112 -49751
rect 146 -50927 158 -49751
rect 100 -50939 158 -50927
rect -158 -51169 -100 -51157
rect -158 -52345 -146 -51169
rect -112 -52345 -100 -51169
rect -158 -52357 -100 -52345
rect 100 -51169 158 -51157
rect 100 -52345 112 -51169
rect 146 -52345 158 -51169
rect 100 -52357 158 -52345
rect -158 -52587 -100 -52575
rect -158 -53763 -146 -52587
rect -112 -53763 -100 -52587
rect -158 -53775 -100 -53763
rect 100 -52587 158 -52575
rect 100 -53763 112 -52587
rect 146 -53763 158 -52587
rect 100 -53775 158 -53763
rect -158 -54005 -100 -53993
rect -158 -55181 -146 -54005
rect -112 -55181 -100 -54005
rect -158 -55193 -100 -55181
rect 100 -54005 158 -53993
rect 100 -55181 112 -54005
rect 146 -55181 158 -54005
rect 100 -55193 158 -55181
rect -158 -55423 -100 -55411
rect -158 -56599 -146 -55423
rect -112 -56599 -100 -55423
rect -158 -56611 -100 -56599
rect 100 -55423 158 -55411
rect 100 -56599 112 -55423
rect 146 -56599 158 -55423
rect 100 -56611 158 -56599
rect -158 -56841 -100 -56829
rect -158 -58017 -146 -56841
rect -112 -58017 -100 -56841
rect -158 -58029 -100 -58017
rect 100 -56841 158 -56829
rect 100 -58017 112 -56841
rect 146 -58017 158 -56841
rect 100 -58029 158 -58017
rect -158 -58259 -100 -58247
rect -158 -59435 -146 -58259
rect -112 -59435 -100 -58259
rect -158 -59447 -100 -59435
rect 100 -58259 158 -58247
rect 100 -59435 112 -58259
rect 146 -59435 158 -58259
rect 100 -59447 158 -59435
rect -158 -59677 -100 -59665
rect -158 -60853 -146 -59677
rect -112 -60853 -100 -59677
rect -158 -60865 -100 -60853
rect 100 -59677 158 -59665
rect 100 -60853 112 -59677
rect 146 -60853 158 -59677
rect 100 -60865 158 -60853
rect -158 -61095 -100 -61083
rect -158 -62271 -146 -61095
rect -112 -62271 -100 -61095
rect -158 -62283 -100 -62271
rect 100 -61095 158 -61083
rect 100 -62271 112 -61095
rect 146 -62271 158 -61095
rect 100 -62283 158 -62271
rect -158 -62513 -100 -62501
rect -158 -63689 -146 -62513
rect -112 -63689 -100 -62513
rect -158 -63701 -100 -63689
rect 100 -62513 158 -62501
rect 100 -63689 112 -62513
rect 146 -63689 158 -62513
rect 100 -63701 158 -63689
rect -158 -63931 -100 -63919
rect -158 -65107 -146 -63931
rect -112 -65107 -100 -63931
rect -158 -65119 -100 -65107
rect 100 -63931 158 -63919
rect 100 -65107 112 -63931
rect 146 -65107 158 -63931
rect 100 -65119 158 -65107
rect -158 -65349 -100 -65337
rect -158 -66525 -146 -65349
rect -112 -66525 -100 -65349
rect -158 -66537 -100 -66525
rect 100 -65349 158 -65337
rect 100 -66525 112 -65349
rect 146 -66525 158 -65349
rect 100 -66537 158 -66525
rect -158 -66767 -100 -66755
rect -158 -67943 -146 -66767
rect -112 -67943 -100 -66767
rect -158 -67955 -100 -67943
rect 100 -66767 158 -66755
rect 100 -67943 112 -66767
rect 146 -67943 158 -66767
rect 100 -67955 158 -67943
rect -158 -68185 -100 -68173
rect -158 -69361 -146 -68185
rect -112 -69361 -100 -68185
rect -158 -69373 -100 -69361
rect 100 -68185 158 -68173
rect 100 -69361 112 -68185
rect 146 -69361 158 -68185
rect 100 -69373 158 -69361
rect -158 -69603 -100 -69591
rect -158 -70779 -146 -69603
rect -112 -70779 -100 -69603
rect -158 -70791 -100 -70779
rect 100 -69603 158 -69591
rect 100 -70779 112 -69603
rect 146 -70779 158 -69603
rect 100 -70791 158 -70779
rect -158 -71021 -100 -71009
rect -158 -72197 -146 -71021
rect -112 -72197 -100 -71021
rect -158 -72209 -100 -72197
rect 100 -71021 158 -71009
rect 100 -72197 112 -71021
rect 146 -72197 158 -71021
rect 100 -72209 158 -72197
rect -158 -72439 -100 -72427
rect -158 -73615 -146 -72439
rect -112 -73615 -100 -72439
rect -158 -73627 -100 -73615
rect 100 -72439 158 -72427
rect 100 -73615 112 -72439
rect 146 -73615 158 -72439
rect 100 -73627 158 -73615
rect -158 -73857 -100 -73845
rect -158 -75033 -146 -73857
rect -112 -75033 -100 -73857
rect -158 -75045 -100 -75033
rect 100 -73857 158 -73845
rect 100 -75033 112 -73857
rect 146 -75033 158 -73857
rect 100 -75045 158 -75033
rect -158 -75275 -100 -75263
rect -158 -76451 -146 -75275
rect -112 -76451 -100 -75275
rect -158 -76463 -100 -76451
rect 100 -75275 158 -75263
rect 100 -76451 112 -75275
rect 146 -76451 158 -75275
rect 100 -76463 158 -76451
rect -158 -76693 -100 -76681
rect -158 -77869 -146 -76693
rect -112 -77869 -100 -76693
rect -158 -77881 -100 -77869
rect 100 -76693 158 -76681
rect 100 -77869 112 -76693
rect 146 -77869 158 -76693
rect 100 -77881 158 -77869
rect -158 -78111 -100 -78099
rect -158 -79287 -146 -78111
rect -112 -79287 -100 -78111
rect -158 -79299 -100 -79287
rect 100 -78111 158 -78099
rect 100 -79287 112 -78111
rect 146 -79287 158 -78111
rect 100 -79299 158 -79287
rect -158 -79529 -100 -79517
rect -158 -80705 -146 -79529
rect -112 -80705 -100 -79529
rect -158 -80717 -100 -80705
rect 100 -79529 158 -79517
rect 100 -80705 112 -79529
rect 146 -80705 158 -79529
rect 100 -80717 158 -80705
rect -158 -80947 -100 -80935
rect -158 -82123 -146 -80947
rect -112 -82123 -100 -80947
rect -158 -82135 -100 -82123
rect 100 -80947 158 -80935
rect 100 -82123 112 -80947
rect 146 -82123 158 -80947
rect 100 -82135 158 -82123
rect -158 -82365 -100 -82353
rect -158 -83541 -146 -82365
rect -112 -83541 -100 -82365
rect -158 -83553 -100 -83541
rect 100 -82365 158 -82353
rect 100 -83541 112 -82365
rect 146 -83541 158 -82365
rect 100 -83553 158 -83541
rect -158 -83783 -100 -83771
rect -158 -84959 -146 -83783
rect -112 -84959 -100 -83783
rect -158 -84971 -100 -84959
rect 100 -83783 158 -83771
rect 100 -84959 112 -83783
rect 146 -84959 158 -83783
rect 100 -84971 158 -84959
rect -158 -85201 -100 -85189
rect -158 -86377 -146 -85201
rect -112 -86377 -100 -85201
rect -158 -86389 -100 -86377
rect 100 -85201 158 -85189
rect 100 -86377 112 -85201
rect 146 -86377 158 -85201
rect 100 -86389 158 -86377
rect -158 -86619 -100 -86607
rect -158 -87795 -146 -86619
rect -112 -87795 -100 -86619
rect -158 -87807 -100 -87795
rect 100 -86619 158 -86607
rect 100 -87795 112 -86619
rect 146 -87795 158 -86619
rect 100 -87807 158 -87795
rect -158 -88037 -100 -88025
rect -158 -89213 -146 -88037
rect -112 -89213 -100 -88037
rect -158 -89225 -100 -89213
rect 100 -88037 158 -88025
rect 100 -89213 112 -88037
rect 146 -89213 158 -88037
rect 100 -89225 158 -89213
rect -158 -89455 -100 -89443
rect -158 -90631 -146 -89455
rect -112 -90631 -100 -89455
rect -158 -90643 -100 -90631
rect 100 -89455 158 -89443
rect 100 -90631 112 -89455
rect 146 -90631 158 -89455
rect 100 -90643 158 -90631
rect -158 -90873 -100 -90861
rect -158 -92049 -146 -90873
rect -112 -92049 -100 -90873
rect -158 -92061 -100 -92049
rect 100 -90873 158 -90861
rect 100 -92049 112 -90873
rect 146 -92049 158 -90873
rect 100 -92061 158 -92049
rect -158 -92291 -100 -92279
rect -158 -93467 -146 -92291
rect -112 -93467 -100 -92291
rect -158 -93479 -100 -93467
rect 100 -92291 158 -92279
rect 100 -93467 112 -92291
rect 146 -93467 158 -92291
rect 100 -93479 158 -93467
rect -158 -93709 -100 -93697
rect -158 -94885 -146 -93709
rect -112 -94885 -100 -93709
rect -158 -94897 -100 -94885
rect 100 -93709 158 -93697
rect 100 -94885 112 -93709
rect 146 -94885 158 -93709
rect 100 -94897 158 -94885
rect -158 -95127 -100 -95115
rect -158 -96303 -146 -95127
rect -112 -96303 -100 -95127
rect -158 -96315 -100 -96303
rect 100 -95127 158 -95115
rect 100 -96303 112 -95127
rect 146 -96303 158 -95127
rect 100 -96315 158 -96303
rect -158 -96545 -100 -96533
rect -158 -97721 -146 -96545
rect -112 -97721 -100 -96545
rect -158 -97733 -100 -97721
rect 100 -96545 158 -96533
rect 100 -97721 112 -96545
rect 146 -97721 158 -96545
rect 100 -97733 158 -97721
rect -158 -97963 -100 -97951
rect -158 -99139 -146 -97963
rect -112 -99139 -100 -97963
rect -158 -99151 -100 -99139
rect 100 -97963 158 -97951
rect 100 -99139 112 -97963
rect 146 -99139 158 -97963
rect 100 -99151 158 -99139
rect -158 -99381 -100 -99369
rect -158 -100557 -146 -99381
rect -112 -100557 -100 -99381
rect -158 -100569 -100 -100557
rect 100 -99381 158 -99369
rect 100 -100557 112 -99381
rect 146 -100557 158 -99381
rect 100 -100569 158 -100557
rect -158 -100799 -100 -100787
rect -158 -101975 -146 -100799
rect -112 -101975 -100 -100799
rect -158 -101987 -100 -101975
rect 100 -100799 158 -100787
rect 100 -101975 112 -100799
rect 146 -101975 158 -100799
rect 100 -101987 158 -101975
rect -158 -102217 -100 -102205
rect -158 -103393 -146 -102217
rect -112 -103393 -100 -102217
rect -158 -103405 -100 -103393
rect 100 -102217 158 -102205
rect 100 -103393 112 -102217
rect 146 -103393 158 -102217
rect 100 -103405 158 -103393
rect -158 -103635 -100 -103623
rect -158 -104811 -146 -103635
rect -112 -104811 -100 -103635
rect -158 -104823 -100 -104811
rect 100 -103635 158 -103623
rect 100 -104811 112 -103635
rect 146 -104811 158 -103635
rect 100 -104823 158 -104811
rect -158 -105053 -100 -105041
rect -158 -106229 -146 -105053
rect -112 -106229 -100 -105053
rect -158 -106241 -100 -106229
rect 100 -105053 158 -105041
rect 100 -106229 112 -105053
rect 146 -106229 158 -105053
rect 100 -106241 158 -106229
rect -158 -106471 -100 -106459
rect -158 -107647 -146 -106471
rect -112 -107647 -100 -106471
rect -158 -107659 -100 -107647
rect 100 -106471 158 -106459
rect 100 -107647 112 -106471
rect 146 -107647 158 -106471
rect 100 -107659 158 -107647
rect -158 -107889 -100 -107877
rect -158 -109065 -146 -107889
rect -112 -109065 -100 -107889
rect -158 -109077 -100 -109065
rect 100 -107889 158 -107877
rect 100 -109065 112 -107889
rect 146 -109065 158 -107889
rect 100 -109077 158 -109065
rect -158 -109307 -100 -109295
rect -158 -110483 -146 -109307
rect -112 -110483 -100 -109307
rect -158 -110495 -100 -110483
rect 100 -109307 158 -109295
rect 100 -110483 112 -109307
rect 146 -110483 158 -109307
rect 100 -110495 158 -110483
rect -158 -110725 -100 -110713
rect -158 -111901 -146 -110725
rect -112 -111901 -100 -110725
rect -158 -111913 -100 -111901
rect 100 -110725 158 -110713
rect 100 -111901 112 -110725
rect 146 -111901 158 -110725
rect 100 -111913 158 -111901
rect -158 -112143 -100 -112131
rect -158 -113319 -146 -112143
rect -112 -113319 -100 -112143
rect -158 -113331 -100 -113319
rect 100 -112143 158 -112131
rect 100 -113319 112 -112143
rect 146 -113319 158 -112143
rect 100 -113331 158 -113319
rect -158 -113561 -100 -113549
rect -158 -114737 -146 -113561
rect -112 -114737 -100 -113561
rect -158 -114749 -100 -114737
rect 100 -113561 158 -113549
rect 100 -114737 112 -113561
rect 146 -114737 158 -113561
rect 100 -114749 158 -114737
rect -158 -114979 -100 -114967
rect -158 -116155 -146 -114979
rect -112 -116155 -100 -114979
rect -158 -116167 -100 -116155
rect 100 -114979 158 -114967
rect 100 -116155 112 -114979
rect 146 -116155 158 -114979
rect 100 -116167 158 -116155
rect -158 -116397 -100 -116385
rect -158 -117573 -146 -116397
rect -112 -117573 -100 -116397
rect -158 -117585 -100 -117573
rect 100 -116397 158 -116385
rect 100 -117573 112 -116397
rect 146 -117573 158 -116397
rect 100 -117585 158 -117573
rect -158 -117815 -100 -117803
rect -158 -118991 -146 -117815
rect -112 -118991 -100 -117815
rect -158 -119003 -100 -118991
rect 100 -117815 158 -117803
rect 100 -118991 112 -117815
rect 146 -118991 158 -117815
rect 100 -119003 158 -118991
rect -158 -119233 -100 -119221
rect -158 -120409 -146 -119233
rect -112 -120409 -100 -119233
rect -158 -120421 -100 -120409
rect 100 -119233 158 -119221
rect 100 -120409 112 -119233
rect 146 -120409 158 -119233
rect 100 -120421 158 -120409
rect -158 -120651 -100 -120639
rect -158 -121827 -146 -120651
rect -112 -121827 -100 -120651
rect -158 -121839 -100 -121827
rect 100 -120651 158 -120639
rect 100 -121827 112 -120651
rect 146 -121827 158 -120651
rect 100 -121839 158 -121827
rect -158 -122069 -100 -122057
rect -158 -123245 -146 -122069
rect -112 -123245 -100 -122069
rect -158 -123257 -100 -123245
rect 100 -122069 158 -122057
rect 100 -123245 112 -122069
rect 146 -123245 158 -122069
rect 100 -123257 158 -123245
rect -158 -123487 -100 -123475
rect -158 -124663 -146 -123487
rect -112 -124663 -100 -123487
rect -158 -124675 -100 -124663
rect 100 -123487 158 -123475
rect 100 -124663 112 -123487
rect 146 -124663 158 -123487
rect 100 -124675 158 -124663
rect -158 -124905 -100 -124893
rect -158 -126081 -146 -124905
rect -112 -126081 -100 -124905
rect -158 -126093 -100 -126081
rect 100 -124905 158 -124893
rect 100 -126081 112 -124905
rect 146 -126081 158 -124905
rect 100 -126093 158 -126081
rect -158 -126323 -100 -126311
rect -158 -127499 -146 -126323
rect -112 -127499 -100 -126323
rect -158 -127511 -100 -127499
rect 100 -126323 158 -126311
rect 100 -127499 112 -126323
rect 146 -127499 158 -126323
rect 100 -127511 158 -127499
rect -158 -127741 -100 -127729
rect -158 -128917 -146 -127741
rect -112 -128917 -100 -127741
rect -158 -128929 -100 -128917
rect 100 -127741 158 -127729
rect 100 -128917 112 -127741
rect 146 -128917 158 -127741
rect 100 -128929 158 -128917
rect -158 -129159 -100 -129147
rect -158 -130335 -146 -129159
rect -112 -130335 -100 -129159
rect -158 -130347 -100 -130335
rect 100 -129159 158 -129147
rect 100 -130335 112 -129159
rect 146 -130335 158 -129159
rect 100 -130347 158 -130335
rect -158 -130577 -100 -130565
rect -158 -131753 -146 -130577
rect -112 -131753 -100 -130577
rect -158 -131765 -100 -131753
rect 100 -130577 158 -130565
rect 100 -131753 112 -130577
rect 146 -131753 158 -130577
rect 100 -131765 158 -131753
rect -158 -131995 -100 -131983
rect -158 -133171 -146 -131995
rect -112 -133171 -100 -131995
rect -158 -133183 -100 -133171
rect 100 -131995 158 -131983
rect 100 -133171 112 -131995
rect 146 -133171 158 -131995
rect 100 -133183 158 -133171
rect -158 -133413 -100 -133401
rect -158 -134589 -146 -133413
rect -112 -134589 -100 -133413
rect -158 -134601 -100 -134589
rect 100 -133413 158 -133401
rect 100 -134589 112 -133413
rect 146 -134589 158 -133413
rect 100 -134601 158 -134589
rect -158 -134831 -100 -134819
rect -158 -136007 -146 -134831
rect -112 -136007 -100 -134831
rect -158 -136019 -100 -136007
rect 100 -134831 158 -134819
rect 100 -136007 112 -134831
rect 146 -136007 158 -134831
rect 100 -136019 158 -136007
rect -158 -136249 -100 -136237
rect -158 -137425 -146 -136249
rect -112 -137425 -100 -136249
rect -158 -137437 -100 -137425
rect 100 -136249 158 -136237
rect 100 -137425 112 -136249
rect 146 -137425 158 -136249
rect 100 -137437 158 -137425
rect -158 -137667 -100 -137655
rect -158 -138843 -146 -137667
rect -112 -138843 -100 -137667
rect -158 -138855 -100 -138843
rect 100 -137667 158 -137655
rect 100 -138843 112 -137667
rect 146 -138843 158 -137667
rect 100 -138855 158 -138843
rect -158 -139085 -100 -139073
rect -158 -140261 -146 -139085
rect -112 -140261 -100 -139085
rect -158 -140273 -100 -140261
rect 100 -139085 158 -139073
rect 100 -140261 112 -139085
rect 146 -140261 158 -139085
rect 100 -140273 158 -140261
rect -158 -140503 -100 -140491
rect -158 -141679 -146 -140503
rect -112 -141679 -100 -140503
rect -158 -141691 -100 -141679
rect 100 -140503 158 -140491
rect 100 -141679 112 -140503
rect 146 -141679 158 -140503
rect 100 -141691 158 -141679
rect -158 -141921 -100 -141909
rect -158 -143097 -146 -141921
rect -112 -143097 -100 -141921
rect -158 -143109 -100 -143097
rect 100 -141921 158 -141909
rect 100 -143097 112 -141921
rect 146 -143097 158 -141921
rect 100 -143109 158 -143097
rect -158 -143339 -100 -143327
rect -158 -144515 -146 -143339
rect -112 -144515 -100 -143339
rect -158 -144527 -100 -144515
rect 100 -143339 158 -143327
rect 100 -144515 112 -143339
rect 146 -144515 158 -143339
rect 100 -144527 158 -144515
rect -158 -144757 -100 -144745
rect -158 -145933 -146 -144757
rect -112 -145933 -100 -144757
rect -158 -145945 -100 -145933
rect 100 -144757 158 -144745
rect 100 -145933 112 -144757
rect 146 -145933 158 -144757
rect 100 -145945 158 -145933
rect -158 -146175 -100 -146163
rect -158 -147351 -146 -146175
rect -112 -147351 -100 -146175
rect -158 -147363 -100 -147351
rect 100 -146175 158 -146163
rect 100 -147351 112 -146175
rect 146 -147351 158 -146175
rect 100 -147363 158 -147351
rect -158 -147593 -100 -147581
rect -158 -148769 -146 -147593
rect -112 -148769 -100 -147593
rect -158 -148781 -100 -148769
rect 100 -147593 158 -147581
rect 100 -148769 112 -147593
rect 146 -148769 158 -147593
rect 100 -148781 158 -148769
rect -158 -149011 -100 -148999
rect -158 -150187 -146 -149011
rect -112 -150187 -100 -149011
rect -158 -150199 -100 -150187
rect 100 -149011 158 -148999
rect 100 -150187 112 -149011
rect 146 -150187 158 -149011
rect 100 -150199 158 -150187
rect -158 -150429 -100 -150417
rect -158 -151605 -146 -150429
rect -112 -151605 -100 -150429
rect -158 -151617 -100 -151605
rect 100 -150429 158 -150417
rect 100 -151605 112 -150429
rect 146 -151605 158 -150429
rect 100 -151617 158 -151605
rect -158 -151847 -100 -151835
rect -158 -153023 -146 -151847
rect -112 -153023 -100 -151847
rect -158 -153035 -100 -153023
rect 100 -151847 158 -151835
rect 100 -153023 112 -151847
rect 146 -153023 158 -151847
rect 100 -153035 158 -153023
rect -158 -153265 -100 -153253
rect -158 -154441 -146 -153265
rect -112 -154441 -100 -153265
rect -158 -154453 -100 -154441
rect 100 -153265 158 -153253
rect 100 -154441 112 -153265
rect 146 -154441 158 -153265
rect 100 -154453 158 -154441
rect -158 -154683 -100 -154671
rect -158 -155859 -146 -154683
rect -112 -155859 -100 -154683
rect -158 -155871 -100 -155859
rect 100 -154683 158 -154671
rect 100 -155859 112 -154683
rect 146 -155859 158 -154683
rect 100 -155871 158 -155859
rect -158 -156101 -100 -156089
rect -158 -157277 -146 -156101
rect -112 -157277 -100 -156101
rect -158 -157289 -100 -157277
rect 100 -156101 158 -156089
rect 100 -157277 112 -156101
rect 146 -157277 158 -156101
rect 100 -157289 158 -157277
rect -158 -157519 -100 -157507
rect -158 -158695 -146 -157519
rect -112 -158695 -100 -157519
rect -158 -158707 -100 -158695
rect 100 -157519 158 -157507
rect 100 -158695 112 -157519
rect 146 -158695 158 -157519
rect 100 -158707 158 -158695
rect -158 -158937 -100 -158925
rect -158 -160113 -146 -158937
rect -112 -160113 -100 -158937
rect -158 -160125 -100 -160113
rect 100 -158937 158 -158925
rect 100 -160113 112 -158937
rect 146 -160113 158 -158937
rect 100 -160125 158 -160113
rect -158 -160355 -100 -160343
rect -158 -161531 -146 -160355
rect -112 -161531 -100 -160355
rect -158 -161543 -100 -161531
rect 100 -160355 158 -160343
rect 100 -161531 112 -160355
rect 146 -161531 158 -160355
rect 100 -161543 158 -161531
rect -158 -161773 -100 -161761
rect -158 -162949 -146 -161773
rect -112 -162949 -100 -161773
rect -158 -162961 -100 -162949
rect 100 -161773 158 -161761
rect 100 -162949 112 -161773
rect 146 -162949 158 -161773
rect 100 -162961 158 -162949
rect -158 -163191 -100 -163179
rect -158 -164367 -146 -163191
rect -112 -164367 -100 -163191
rect -158 -164379 -100 -164367
rect 100 -163191 158 -163179
rect 100 -164367 112 -163191
rect 146 -164367 158 -163191
rect 100 -164379 158 -164367
rect -158 -164609 -100 -164597
rect -158 -165785 -146 -164609
rect -112 -165785 -100 -164609
rect -158 -165797 -100 -165785
rect 100 -164609 158 -164597
rect 100 -165785 112 -164609
rect 146 -165785 158 -164609
rect 100 -165797 158 -165785
rect -158 -166027 -100 -166015
rect -158 -167203 -146 -166027
rect -112 -167203 -100 -166027
rect -158 -167215 -100 -167203
rect 100 -166027 158 -166015
rect 100 -167203 112 -166027
rect 146 -167203 158 -166027
rect 100 -167215 158 -167203
rect -158 -167445 -100 -167433
rect -158 -168621 -146 -167445
rect -112 -168621 -100 -167445
rect -158 -168633 -100 -168621
rect 100 -167445 158 -167433
rect 100 -168621 112 -167445
rect 146 -168621 158 -167445
rect 100 -168633 158 -168621
rect -158 -168863 -100 -168851
rect -158 -170039 -146 -168863
rect -112 -170039 -100 -168863
rect -158 -170051 -100 -170039
rect 100 -168863 158 -168851
rect 100 -170039 112 -168863
rect 146 -170039 158 -168863
rect 100 -170051 158 -170039
rect -158 -170281 -100 -170269
rect -158 -171457 -146 -170281
rect -112 -171457 -100 -170281
rect -158 -171469 -100 -171457
rect 100 -170281 158 -170269
rect 100 -171457 112 -170281
rect 146 -171457 158 -170281
rect 100 -171469 158 -171457
rect -158 -171699 -100 -171687
rect -158 -172875 -146 -171699
rect -112 -172875 -100 -171699
rect -158 -172887 -100 -172875
rect 100 -171699 158 -171687
rect 100 -172875 112 -171699
rect 146 -172875 158 -171699
rect 100 -172887 158 -172875
rect -158 -173117 -100 -173105
rect -158 -174293 -146 -173117
rect -112 -174293 -100 -173117
rect -158 -174305 -100 -174293
rect 100 -173117 158 -173105
rect 100 -174293 112 -173117
rect 146 -174293 158 -173117
rect 100 -174305 158 -174293
rect -158 -174535 -100 -174523
rect -158 -175711 -146 -174535
rect -112 -175711 -100 -174535
rect -158 -175723 -100 -175711
rect 100 -174535 158 -174523
rect 100 -175711 112 -174535
rect 146 -175711 158 -174535
rect 100 -175723 158 -175711
rect -158 -175953 -100 -175941
rect -158 -177129 -146 -175953
rect -112 -177129 -100 -175953
rect -158 -177141 -100 -177129
rect 100 -175953 158 -175941
rect 100 -177129 112 -175953
rect 146 -177129 158 -175953
rect 100 -177141 158 -177129
rect -158 -177371 -100 -177359
rect -158 -178547 -146 -177371
rect -112 -178547 -100 -177371
rect -158 -178559 -100 -178547
rect 100 -177371 158 -177359
rect 100 -178547 112 -177371
rect 146 -178547 158 -177371
rect 100 -178559 158 -178547
rect -158 -178789 -100 -178777
rect -158 -179965 -146 -178789
rect -112 -179965 -100 -178789
rect -158 -179977 -100 -179965
rect 100 -178789 158 -178777
rect 100 -179965 112 -178789
rect 146 -179965 158 -178789
rect 100 -179977 158 -179965
rect -158 -180207 -100 -180195
rect -158 -181383 -146 -180207
rect -112 -181383 -100 -180207
rect -158 -181395 -100 -181383
rect 100 -180207 158 -180195
rect 100 -181383 112 -180207
rect 146 -181383 158 -180207
rect 100 -181395 158 -181383
<< mvndiffc >>
rect -146 180207 -112 181383
rect 112 180207 146 181383
rect -146 178789 -112 179965
rect 112 178789 146 179965
rect -146 177371 -112 178547
rect 112 177371 146 178547
rect -146 175953 -112 177129
rect 112 175953 146 177129
rect -146 174535 -112 175711
rect 112 174535 146 175711
rect -146 173117 -112 174293
rect 112 173117 146 174293
rect -146 171699 -112 172875
rect 112 171699 146 172875
rect -146 170281 -112 171457
rect 112 170281 146 171457
rect -146 168863 -112 170039
rect 112 168863 146 170039
rect -146 167445 -112 168621
rect 112 167445 146 168621
rect -146 166027 -112 167203
rect 112 166027 146 167203
rect -146 164609 -112 165785
rect 112 164609 146 165785
rect -146 163191 -112 164367
rect 112 163191 146 164367
rect -146 161773 -112 162949
rect 112 161773 146 162949
rect -146 160355 -112 161531
rect 112 160355 146 161531
rect -146 158937 -112 160113
rect 112 158937 146 160113
rect -146 157519 -112 158695
rect 112 157519 146 158695
rect -146 156101 -112 157277
rect 112 156101 146 157277
rect -146 154683 -112 155859
rect 112 154683 146 155859
rect -146 153265 -112 154441
rect 112 153265 146 154441
rect -146 151847 -112 153023
rect 112 151847 146 153023
rect -146 150429 -112 151605
rect 112 150429 146 151605
rect -146 149011 -112 150187
rect 112 149011 146 150187
rect -146 147593 -112 148769
rect 112 147593 146 148769
rect -146 146175 -112 147351
rect 112 146175 146 147351
rect -146 144757 -112 145933
rect 112 144757 146 145933
rect -146 143339 -112 144515
rect 112 143339 146 144515
rect -146 141921 -112 143097
rect 112 141921 146 143097
rect -146 140503 -112 141679
rect 112 140503 146 141679
rect -146 139085 -112 140261
rect 112 139085 146 140261
rect -146 137667 -112 138843
rect 112 137667 146 138843
rect -146 136249 -112 137425
rect 112 136249 146 137425
rect -146 134831 -112 136007
rect 112 134831 146 136007
rect -146 133413 -112 134589
rect 112 133413 146 134589
rect -146 131995 -112 133171
rect 112 131995 146 133171
rect -146 130577 -112 131753
rect 112 130577 146 131753
rect -146 129159 -112 130335
rect 112 129159 146 130335
rect -146 127741 -112 128917
rect 112 127741 146 128917
rect -146 126323 -112 127499
rect 112 126323 146 127499
rect -146 124905 -112 126081
rect 112 124905 146 126081
rect -146 123487 -112 124663
rect 112 123487 146 124663
rect -146 122069 -112 123245
rect 112 122069 146 123245
rect -146 120651 -112 121827
rect 112 120651 146 121827
rect -146 119233 -112 120409
rect 112 119233 146 120409
rect -146 117815 -112 118991
rect 112 117815 146 118991
rect -146 116397 -112 117573
rect 112 116397 146 117573
rect -146 114979 -112 116155
rect 112 114979 146 116155
rect -146 113561 -112 114737
rect 112 113561 146 114737
rect -146 112143 -112 113319
rect 112 112143 146 113319
rect -146 110725 -112 111901
rect 112 110725 146 111901
rect -146 109307 -112 110483
rect 112 109307 146 110483
rect -146 107889 -112 109065
rect 112 107889 146 109065
rect -146 106471 -112 107647
rect 112 106471 146 107647
rect -146 105053 -112 106229
rect 112 105053 146 106229
rect -146 103635 -112 104811
rect 112 103635 146 104811
rect -146 102217 -112 103393
rect 112 102217 146 103393
rect -146 100799 -112 101975
rect 112 100799 146 101975
rect -146 99381 -112 100557
rect 112 99381 146 100557
rect -146 97963 -112 99139
rect 112 97963 146 99139
rect -146 96545 -112 97721
rect 112 96545 146 97721
rect -146 95127 -112 96303
rect 112 95127 146 96303
rect -146 93709 -112 94885
rect 112 93709 146 94885
rect -146 92291 -112 93467
rect 112 92291 146 93467
rect -146 90873 -112 92049
rect 112 90873 146 92049
rect -146 89455 -112 90631
rect 112 89455 146 90631
rect -146 88037 -112 89213
rect 112 88037 146 89213
rect -146 86619 -112 87795
rect 112 86619 146 87795
rect -146 85201 -112 86377
rect 112 85201 146 86377
rect -146 83783 -112 84959
rect 112 83783 146 84959
rect -146 82365 -112 83541
rect 112 82365 146 83541
rect -146 80947 -112 82123
rect 112 80947 146 82123
rect -146 79529 -112 80705
rect 112 79529 146 80705
rect -146 78111 -112 79287
rect 112 78111 146 79287
rect -146 76693 -112 77869
rect 112 76693 146 77869
rect -146 75275 -112 76451
rect 112 75275 146 76451
rect -146 73857 -112 75033
rect 112 73857 146 75033
rect -146 72439 -112 73615
rect 112 72439 146 73615
rect -146 71021 -112 72197
rect 112 71021 146 72197
rect -146 69603 -112 70779
rect 112 69603 146 70779
rect -146 68185 -112 69361
rect 112 68185 146 69361
rect -146 66767 -112 67943
rect 112 66767 146 67943
rect -146 65349 -112 66525
rect 112 65349 146 66525
rect -146 63931 -112 65107
rect 112 63931 146 65107
rect -146 62513 -112 63689
rect 112 62513 146 63689
rect -146 61095 -112 62271
rect 112 61095 146 62271
rect -146 59677 -112 60853
rect 112 59677 146 60853
rect -146 58259 -112 59435
rect 112 58259 146 59435
rect -146 56841 -112 58017
rect 112 56841 146 58017
rect -146 55423 -112 56599
rect 112 55423 146 56599
rect -146 54005 -112 55181
rect 112 54005 146 55181
rect -146 52587 -112 53763
rect 112 52587 146 53763
rect -146 51169 -112 52345
rect 112 51169 146 52345
rect -146 49751 -112 50927
rect 112 49751 146 50927
rect -146 48333 -112 49509
rect 112 48333 146 49509
rect -146 46915 -112 48091
rect 112 46915 146 48091
rect -146 45497 -112 46673
rect 112 45497 146 46673
rect -146 44079 -112 45255
rect 112 44079 146 45255
rect -146 42661 -112 43837
rect 112 42661 146 43837
rect -146 41243 -112 42419
rect 112 41243 146 42419
rect -146 39825 -112 41001
rect 112 39825 146 41001
rect -146 38407 -112 39583
rect 112 38407 146 39583
rect -146 36989 -112 38165
rect 112 36989 146 38165
rect -146 35571 -112 36747
rect 112 35571 146 36747
rect -146 34153 -112 35329
rect 112 34153 146 35329
rect -146 32735 -112 33911
rect 112 32735 146 33911
rect -146 31317 -112 32493
rect 112 31317 146 32493
rect -146 29899 -112 31075
rect 112 29899 146 31075
rect -146 28481 -112 29657
rect 112 28481 146 29657
rect -146 27063 -112 28239
rect 112 27063 146 28239
rect -146 25645 -112 26821
rect 112 25645 146 26821
rect -146 24227 -112 25403
rect 112 24227 146 25403
rect -146 22809 -112 23985
rect 112 22809 146 23985
rect -146 21391 -112 22567
rect 112 21391 146 22567
rect -146 19973 -112 21149
rect 112 19973 146 21149
rect -146 18555 -112 19731
rect 112 18555 146 19731
rect -146 17137 -112 18313
rect 112 17137 146 18313
rect -146 15719 -112 16895
rect 112 15719 146 16895
rect -146 14301 -112 15477
rect 112 14301 146 15477
rect -146 12883 -112 14059
rect 112 12883 146 14059
rect -146 11465 -112 12641
rect 112 11465 146 12641
rect -146 10047 -112 11223
rect 112 10047 146 11223
rect -146 8629 -112 9805
rect 112 8629 146 9805
rect -146 7211 -112 8387
rect 112 7211 146 8387
rect -146 5793 -112 6969
rect 112 5793 146 6969
rect -146 4375 -112 5551
rect 112 4375 146 5551
rect -146 2957 -112 4133
rect 112 2957 146 4133
rect -146 1539 -112 2715
rect 112 1539 146 2715
rect -146 121 -112 1297
rect 112 121 146 1297
rect -146 -1297 -112 -121
rect 112 -1297 146 -121
rect -146 -2715 -112 -1539
rect 112 -2715 146 -1539
rect -146 -4133 -112 -2957
rect 112 -4133 146 -2957
rect -146 -5551 -112 -4375
rect 112 -5551 146 -4375
rect -146 -6969 -112 -5793
rect 112 -6969 146 -5793
rect -146 -8387 -112 -7211
rect 112 -8387 146 -7211
rect -146 -9805 -112 -8629
rect 112 -9805 146 -8629
rect -146 -11223 -112 -10047
rect 112 -11223 146 -10047
rect -146 -12641 -112 -11465
rect 112 -12641 146 -11465
rect -146 -14059 -112 -12883
rect 112 -14059 146 -12883
rect -146 -15477 -112 -14301
rect 112 -15477 146 -14301
rect -146 -16895 -112 -15719
rect 112 -16895 146 -15719
rect -146 -18313 -112 -17137
rect 112 -18313 146 -17137
rect -146 -19731 -112 -18555
rect 112 -19731 146 -18555
rect -146 -21149 -112 -19973
rect 112 -21149 146 -19973
rect -146 -22567 -112 -21391
rect 112 -22567 146 -21391
rect -146 -23985 -112 -22809
rect 112 -23985 146 -22809
rect -146 -25403 -112 -24227
rect 112 -25403 146 -24227
rect -146 -26821 -112 -25645
rect 112 -26821 146 -25645
rect -146 -28239 -112 -27063
rect 112 -28239 146 -27063
rect -146 -29657 -112 -28481
rect 112 -29657 146 -28481
rect -146 -31075 -112 -29899
rect 112 -31075 146 -29899
rect -146 -32493 -112 -31317
rect 112 -32493 146 -31317
rect -146 -33911 -112 -32735
rect 112 -33911 146 -32735
rect -146 -35329 -112 -34153
rect 112 -35329 146 -34153
rect -146 -36747 -112 -35571
rect 112 -36747 146 -35571
rect -146 -38165 -112 -36989
rect 112 -38165 146 -36989
rect -146 -39583 -112 -38407
rect 112 -39583 146 -38407
rect -146 -41001 -112 -39825
rect 112 -41001 146 -39825
rect -146 -42419 -112 -41243
rect 112 -42419 146 -41243
rect -146 -43837 -112 -42661
rect 112 -43837 146 -42661
rect -146 -45255 -112 -44079
rect 112 -45255 146 -44079
rect -146 -46673 -112 -45497
rect 112 -46673 146 -45497
rect -146 -48091 -112 -46915
rect 112 -48091 146 -46915
rect -146 -49509 -112 -48333
rect 112 -49509 146 -48333
rect -146 -50927 -112 -49751
rect 112 -50927 146 -49751
rect -146 -52345 -112 -51169
rect 112 -52345 146 -51169
rect -146 -53763 -112 -52587
rect 112 -53763 146 -52587
rect -146 -55181 -112 -54005
rect 112 -55181 146 -54005
rect -146 -56599 -112 -55423
rect 112 -56599 146 -55423
rect -146 -58017 -112 -56841
rect 112 -58017 146 -56841
rect -146 -59435 -112 -58259
rect 112 -59435 146 -58259
rect -146 -60853 -112 -59677
rect 112 -60853 146 -59677
rect -146 -62271 -112 -61095
rect 112 -62271 146 -61095
rect -146 -63689 -112 -62513
rect 112 -63689 146 -62513
rect -146 -65107 -112 -63931
rect 112 -65107 146 -63931
rect -146 -66525 -112 -65349
rect 112 -66525 146 -65349
rect -146 -67943 -112 -66767
rect 112 -67943 146 -66767
rect -146 -69361 -112 -68185
rect 112 -69361 146 -68185
rect -146 -70779 -112 -69603
rect 112 -70779 146 -69603
rect -146 -72197 -112 -71021
rect 112 -72197 146 -71021
rect -146 -73615 -112 -72439
rect 112 -73615 146 -72439
rect -146 -75033 -112 -73857
rect 112 -75033 146 -73857
rect -146 -76451 -112 -75275
rect 112 -76451 146 -75275
rect -146 -77869 -112 -76693
rect 112 -77869 146 -76693
rect -146 -79287 -112 -78111
rect 112 -79287 146 -78111
rect -146 -80705 -112 -79529
rect 112 -80705 146 -79529
rect -146 -82123 -112 -80947
rect 112 -82123 146 -80947
rect -146 -83541 -112 -82365
rect 112 -83541 146 -82365
rect -146 -84959 -112 -83783
rect 112 -84959 146 -83783
rect -146 -86377 -112 -85201
rect 112 -86377 146 -85201
rect -146 -87795 -112 -86619
rect 112 -87795 146 -86619
rect -146 -89213 -112 -88037
rect 112 -89213 146 -88037
rect -146 -90631 -112 -89455
rect 112 -90631 146 -89455
rect -146 -92049 -112 -90873
rect 112 -92049 146 -90873
rect -146 -93467 -112 -92291
rect 112 -93467 146 -92291
rect -146 -94885 -112 -93709
rect 112 -94885 146 -93709
rect -146 -96303 -112 -95127
rect 112 -96303 146 -95127
rect -146 -97721 -112 -96545
rect 112 -97721 146 -96545
rect -146 -99139 -112 -97963
rect 112 -99139 146 -97963
rect -146 -100557 -112 -99381
rect 112 -100557 146 -99381
rect -146 -101975 -112 -100799
rect 112 -101975 146 -100799
rect -146 -103393 -112 -102217
rect 112 -103393 146 -102217
rect -146 -104811 -112 -103635
rect 112 -104811 146 -103635
rect -146 -106229 -112 -105053
rect 112 -106229 146 -105053
rect -146 -107647 -112 -106471
rect 112 -107647 146 -106471
rect -146 -109065 -112 -107889
rect 112 -109065 146 -107889
rect -146 -110483 -112 -109307
rect 112 -110483 146 -109307
rect -146 -111901 -112 -110725
rect 112 -111901 146 -110725
rect -146 -113319 -112 -112143
rect 112 -113319 146 -112143
rect -146 -114737 -112 -113561
rect 112 -114737 146 -113561
rect -146 -116155 -112 -114979
rect 112 -116155 146 -114979
rect -146 -117573 -112 -116397
rect 112 -117573 146 -116397
rect -146 -118991 -112 -117815
rect 112 -118991 146 -117815
rect -146 -120409 -112 -119233
rect 112 -120409 146 -119233
rect -146 -121827 -112 -120651
rect 112 -121827 146 -120651
rect -146 -123245 -112 -122069
rect 112 -123245 146 -122069
rect -146 -124663 -112 -123487
rect 112 -124663 146 -123487
rect -146 -126081 -112 -124905
rect 112 -126081 146 -124905
rect -146 -127499 -112 -126323
rect 112 -127499 146 -126323
rect -146 -128917 -112 -127741
rect 112 -128917 146 -127741
rect -146 -130335 -112 -129159
rect 112 -130335 146 -129159
rect -146 -131753 -112 -130577
rect 112 -131753 146 -130577
rect -146 -133171 -112 -131995
rect 112 -133171 146 -131995
rect -146 -134589 -112 -133413
rect 112 -134589 146 -133413
rect -146 -136007 -112 -134831
rect 112 -136007 146 -134831
rect -146 -137425 -112 -136249
rect 112 -137425 146 -136249
rect -146 -138843 -112 -137667
rect 112 -138843 146 -137667
rect -146 -140261 -112 -139085
rect 112 -140261 146 -139085
rect -146 -141679 -112 -140503
rect 112 -141679 146 -140503
rect -146 -143097 -112 -141921
rect 112 -143097 146 -141921
rect -146 -144515 -112 -143339
rect 112 -144515 146 -143339
rect -146 -145933 -112 -144757
rect 112 -145933 146 -144757
rect -146 -147351 -112 -146175
rect 112 -147351 146 -146175
rect -146 -148769 -112 -147593
rect 112 -148769 146 -147593
rect -146 -150187 -112 -149011
rect 112 -150187 146 -149011
rect -146 -151605 -112 -150429
rect 112 -151605 146 -150429
rect -146 -153023 -112 -151847
rect 112 -153023 146 -151847
rect -146 -154441 -112 -153265
rect 112 -154441 146 -153265
rect -146 -155859 -112 -154683
rect 112 -155859 146 -154683
rect -146 -157277 -112 -156101
rect 112 -157277 146 -156101
rect -146 -158695 -112 -157519
rect 112 -158695 146 -157519
rect -146 -160113 -112 -158937
rect 112 -160113 146 -158937
rect -146 -161531 -112 -160355
rect 112 -161531 146 -160355
rect -146 -162949 -112 -161773
rect 112 -162949 146 -161773
rect -146 -164367 -112 -163191
rect 112 -164367 146 -163191
rect -146 -165785 -112 -164609
rect 112 -165785 146 -164609
rect -146 -167203 -112 -166027
rect 112 -167203 146 -166027
rect -146 -168621 -112 -167445
rect 112 -168621 146 -167445
rect -146 -170039 -112 -168863
rect 112 -170039 146 -168863
rect -146 -171457 -112 -170281
rect 112 -171457 146 -170281
rect -146 -172875 -112 -171699
rect 112 -172875 146 -171699
rect -146 -174293 -112 -173117
rect 112 -174293 146 -173117
rect -146 -175711 -112 -174535
rect 112 -175711 146 -174535
rect -146 -177129 -112 -175953
rect 112 -177129 146 -175953
rect -146 -178547 -112 -177371
rect 112 -178547 146 -177371
rect -146 -179965 -112 -178789
rect 112 -179965 146 -178789
rect -146 -181383 -112 -180207
rect 112 -181383 146 -180207
<< mvpsubdiff >>
rect -292 181605 292 181617
rect -292 181571 -184 181605
rect 184 181571 292 181605
rect -292 181559 292 181571
rect -292 181509 -234 181559
rect -292 -181509 -280 181509
rect -246 -181509 -234 181509
rect 234 181509 292 181559
rect -292 -181559 -234 -181509
rect 234 -181509 246 181509
rect 280 -181509 292 181509
rect 234 -181559 292 -181509
rect -292 -181571 292 -181559
rect -292 -181605 -184 -181571
rect 184 -181605 292 -181571
rect -292 -181617 292 -181605
<< mvpsubdiffcont >>
rect -184 181571 184 181605
rect -280 -181509 -246 181509
rect 246 -181509 280 181509
rect -184 -181605 184 -181571
<< poly >>
rect -100 181467 100 181483
rect -100 181433 -84 181467
rect 84 181433 100 181467
rect -100 181395 100 181433
rect -100 180157 100 180195
rect -100 180123 -84 180157
rect 84 180123 100 180157
rect -100 180107 100 180123
rect -100 180049 100 180065
rect -100 180015 -84 180049
rect 84 180015 100 180049
rect -100 179977 100 180015
rect -100 178739 100 178777
rect -100 178705 -84 178739
rect 84 178705 100 178739
rect -100 178689 100 178705
rect -100 178631 100 178647
rect -100 178597 -84 178631
rect 84 178597 100 178631
rect -100 178559 100 178597
rect -100 177321 100 177359
rect -100 177287 -84 177321
rect 84 177287 100 177321
rect -100 177271 100 177287
rect -100 177213 100 177229
rect -100 177179 -84 177213
rect 84 177179 100 177213
rect -100 177141 100 177179
rect -100 175903 100 175941
rect -100 175869 -84 175903
rect 84 175869 100 175903
rect -100 175853 100 175869
rect -100 175795 100 175811
rect -100 175761 -84 175795
rect 84 175761 100 175795
rect -100 175723 100 175761
rect -100 174485 100 174523
rect -100 174451 -84 174485
rect 84 174451 100 174485
rect -100 174435 100 174451
rect -100 174377 100 174393
rect -100 174343 -84 174377
rect 84 174343 100 174377
rect -100 174305 100 174343
rect -100 173067 100 173105
rect -100 173033 -84 173067
rect 84 173033 100 173067
rect -100 173017 100 173033
rect -100 172959 100 172975
rect -100 172925 -84 172959
rect 84 172925 100 172959
rect -100 172887 100 172925
rect -100 171649 100 171687
rect -100 171615 -84 171649
rect 84 171615 100 171649
rect -100 171599 100 171615
rect -100 171541 100 171557
rect -100 171507 -84 171541
rect 84 171507 100 171541
rect -100 171469 100 171507
rect -100 170231 100 170269
rect -100 170197 -84 170231
rect 84 170197 100 170231
rect -100 170181 100 170197
rect -100 170123 100 170139
rect -100 170089 -84 170123
rect 84 170089 100 170123
rect -100 170051 100 170089
rect -100 168813 100 168851
rect -100 168779 -84 168813
rect 84 168779 100 168813
rect -100 168763 100 168779
rect -100 168705 100 168721
rect -100 168671 -84 168705
rect 84 168671 100 168705
rect -100 168633 100 168671
rect -100 167395 100 167433
rect -100 167361 -84 167395
rect 84 167361 100 167395
rect -100 167345 100 167361
rect -100 167287 100 167303
rect -100 167253 -84 167287
rect 84 167253 100 167287
rect -100 167215 100 167253
rect -100 165977 100 166015
rect -100 165943 -84 165977
rect 84 165943 100 165977
rect -100 165927 100 165943
rect -100 165869 100 165885
rect -100 165835 -84 165869
rect 84 165835 100 165869
rect -100 165797 100 165835
rect -100 164559 100 164597
rect -100 164525 -84 164559
rect 84 164525 100 164559
rect -100 164509 100 164525
rect -100 164451 100 164467
rect -100 164417 -84 164451
rect 84 164417 100 164451
rect -100 164379 100 164417
rect -100 163141 100 163179
rect -100 163107 -84 163141
rect 84 163107 100 163141
rect -100 163091 100 163107
rect -100 163033 100 163049
rect -100 162999 -84 163033
rect 84 162999 100 163033
rect -100 162961 100 162999
rect -100 161723 100 161761
rect -100 161689 -84 161723
rect 84 161689 100 161723
rect -100 161673 100 161689
rect -100 161615 100 161631
rect -100 161581 -84 161615
rect 84 161581 100 161615
rect -100 161543 100 161581
rect -100 160305 100 160343
rect -100 160271 -84 160305
rect 84 160271 100 160305
rect -100 160255 100 160271
rect -100 160197 100 160213
rect -100 160163 -84 160197
rect 84 160163 100 160197
rect -100 160125 100 160163
rect -100 158887 100 158925
rect -100 158853 -84 158887
rect 84 158853 100 158887
rect -100 158837 100 158853
rect -100 158779 100 158795
rect -100 158745 -84 158779
rect 84 158745 100 158779
rect -100 158707 100 158745
rect -100 157469 100 157507
rect -100 157435 -84 157469
rect 84 157435 100 157469
rect -100 157419 100 157435
rect -100 157361 100 157377
rect -100 157327 -84 157361
rect 84 157327 100 157361
rect -100 157289 100 157327
rect -100 156051 100 156089
rect -100 156017 -84 156051
rect 84 156017 100 156051
rect -100 156001 100 156017
rect -100 155943 100 155959
rect -100 155909 -84 155943
rect 84 155909 100 155943
rect -100 155871 100 155909
rect -100 154633 100 154671
rect -100 154599 -84 154633
rect 84 154599 100 154633
rect -100 154583 100 154599
rect -100 154525 100 154541
rect -100 154491 -84 154525
rect 84 154491 100 154525
rect -100 154453 100 154491
rect -100 153215 100 153253
rect -100 153181 -84 153215
rect 84 153181 100 153215
rect -100 153165 100 153181
rect -100 153107 100 153123
rect -100 153073 -84 153107
rect 84 153073 100 153107
rect -100 153035 100 153073
rect -100 151797 100 151835
rect -100 151763 -84 151797
rect 84 151763 100 151797
rect -100 151747 100 151763
rect -100 151689 100 151705
rect -100 151655 -84 151689
rect 84 151655 100 151689
rect -100 151617 100 151655
rect -100 150379 100 150417
rect -100 150345 -84 150379
rect 84 150345 100 150379
rect -100 150329 100 150345
rect -100 150271 100 150287
rect -100 150237 -84 150271
rect 84 150237 100 150271
rect -100 150199 100 150237
rect -100 148961 100 148999
rect -100 148927 -84 148961
rect 84 148927 100 148961
rect -100 148911 100 148927
rect -100 148853 100 148869
rect -100 148819 -84 148853
rect 84 148819 100 148853
rect -100 148781 100 148819
rect -100 147543 100 147581
rect -100 147509 -84 147543
rect 84 147509 100 147543
rect -100 147493 100 147509
rect -100 147435 100 147451
rect -100 147401 -84 147435
rect 84 147401 100 147435
rect -100 147363 100 147401
rect -100 146125 100 146163
rect -100 146091 -84 146125
rect 84 146091 100 146125
rect -100 146075 100 146091
rect -100 146017 100 146033
rect -100 145983 -84 146017
rect 84 145983 100 146017
rect -100 145945 100 145983
rect -100 144707 100 144745
rect -100 144673 -84 144707
rect 84 144673 100 144707
rect -100 144657 100 144673
rect -100 144599 100 144615
rect -100 144565 -84 144599
rect 84 144565 100 144599
rect -100 144527 100 144565
rect -100 143289 100 143327
rect -100 143255 -84 143289
rect 84 143255 100 143289
rect -100 143239 100 143255
rect -100 143181 100 143197
rect -100 143147 -84 143181
rect 84 143147 100 143181
rect -100 143109 100 143147
rect -100 141871 100 141909
rect -100 141837 -84 141871
rect 84 141837 100 141871
rect -100 141821 100 141837
rect -100 141763 100 141779
rect -100 141729 -84 141763
rect 84 141729 100 141763
rect -100 141691 100 141729
rect -100 140453 100 140491
rect -100 140419 -84 140453
rect 84 140419 100 140453
rect -100 140403 100 140419
rect -100 140345 100 140361
rect -100 140311 -84 140345
rect 84 140311 100 140345
rect -100 140273 100 140311
rect -100 139035 100 139073
rect -100 139001 -84 139035
rect 84 139001 100 139035
rect -100 138985 100 139001
rect -100 138927 100 138943
rect -100 138893 -84 138927
rect 84 138893 100 138927
rect -100 138855 100 138893
rect -100 137617 100 137655
rect -100 137583 -84 137617
rect 84 137583 100 137617
rect -100 137567 100 137583
rect -100 137509 100 137525
rect -100 137475 -84 137509
rect 84 137475 100 137509
rect -100 137437 100 137475
rect -100 136199 100 136237
rect -100 136165 -84 136199
rect 84 136165 100 136199
rect -100 136149 100 136165
rect -100 136091 100 136107
rect -100 136057 -84 136091
rect 84 136057 100 136091
rect -100 136019 100 136057
rect -100 134781 100 134819
rect -100 134747 -84 134781
rect 84 134747 100 134781
rect -100 134731 100 134747
rect -100 134673 100 134689
rect -100 134639 -84 134673
rect 84 134639 100 134673
rect -100 134601 100 134639
rect -100 133363 100 133401
rect -100 133329 -84 133363
rect 84 133329 100 133363
rect -100 133313 100 133329
rect -100 133255 100 133271
rect -100 133221 -84 133255
rect 84 133221 100 133255
rect -100 133183 100 133221
rect -100 131945 100 131983
rect -100 131911 -84 131945
rect 84 131911 100 131945
rect -100 131895 100 131911
rect -100 131837 100 131853
rect -100 131803 -84 131837
rect 84 131803 100 131837
rect -100 131765 100 131803
rect -100 130527 100 130565
rect -100 130493 -84 130527
rect 84 130493 100 130527
rect -100 130477 100 130493
rect -100 130419 100 130435
rect -100 130385 -84 130419
rect 84 130385 100 130419
rect -100 130347 100 130385
rect -100 129109 100 129147
rect -100 129075 -84 129109
rect 84 129075 100 129109
rect -100 129059 100 129075
rect -100 129001 100 129017
rect -100 128967 -84 129001
rect 84 128967 100 129001
rect -100 128929 100 128967
rect -100 127691 100 127729
rect -100 127657 -84 127691
rect 84 127657 100 127691
rect -100 127641 100 127657
rect -100 127583 100 127599
rect -100 127549 -84 127583
rect 84 127549 100 127583
rect -100 127511 100 127549
rect -100 126273 100 126311
rect -100 126239 -84 126273
rect 84 126239 100 126273
rect -100 126223 100 126239
rect -100 126165 100 126181
rect -100 126131 -84 126165
rect 84 126131 100 126165
rect -100 126093 100 126131
rect -100 124855 100 124893
rect -100 124821 -84 124855
rect 84 124821 100 124855
rect -100 124805 100 124821
rect -100 124747 100 124763
rect -100 124713 -84 124747
rect 84 124713 100 124747
rect -100 124675 100 124713
rect -100 123437 100 123475
rect -100 123403 -84 123437
rect 84 123403 100 123437
rect -100 123387 100 123403
rect -100 123329 100 123345
rect -100 123295 -84 123329
rect 84 123295 100 123329
rect -100 123257 100 123295
rect -100 122019 100 122057
rect -100 121985 -84 122019
rect 84 121985 100 122019
rect -100 121969 100 121985
rect -100 121911 100 121927
rect -100 121877 -84 121911
rect 84 121877 100 121911
rect -100 121839 100 121877
rect -100 120601 100 120639
rect -100 120567 -84 120601
rect 84 120567 100 120601
rect -100 120551 100 120567
rect -100 120493 100 120509
rect -100 120459 -84 120493
rect 84 120459 100 120493
rect -100 120421 100 120459
rect -100 119183 100 119221
rect -100 119149 -84 119183
rect 84 119149 100 119183
rect -100 119133 100 119149
rect -100 119075 100 119091
rect -100 119041 -84 119075
rect 84 119041 100 119075
rect -100 119003 100 119041
rect -100 117765 100 117803
rect -100 117731 -84 117765
rect 84 117731 100 117765
rect -100 117715 100 117731
rect -100 117657 100 117673
rect -100 117623 -84 117657
rect 84 117623 100 117657
rect -100 117585 100 117623
rect -100 116347 100 116385
rect -100 116313 -84 116347
rect 84 116313 100 116347
rect -100 116297 100 116313
rect -100 116239 100 116255
rect -100 116205 -84 116239
rect 84 116205 100 116239
rect -100 116167 100 116205
rect -100 114929 100 114967
rect -100 114895 -84 114929
rect 84 114895 100 114929
rect -100 114879 100 114895
rect -100 114821 100 114837
rect -100 114787 -84 114821
rect 84 114787 100 114821
rect -100 114749 100 114787
rect -100 113511 100 113549
rect -100 113477 -84 113511
rect 84 113477 100 113511
rect -100 113461 100 113477
rect -100 113403 100 113419
rect -100 113369 -84 113403
rect 84 113369 100 113403
rect -100 113331 100 113369
rect -100 112093 100 112131
rect -100 112059 -84 112093
rect 84 112059 100 112093
rect -100 112043 100 112059
rect -100 111985 100 112001
rect -100 111951 -84 111985
rect 84 111951 100 111985
rect -100 111913 100 111951
rect -100 110675 100 110713
rect -100 110641 -84 110675
rect 84 110641 100 110675
rect -100 110625 100 110641
rect -100 110567 100 110583
rect -100 110533 -84 110567
rect 84 110533 100 110567
rect -100 110495 100 110533
rect -100 109257 100 109295
rect -100 109223 -84 109257
rect 84 109223 100 109257
rect -100 109207 100 109223
rect -100 109149 100 109165
rect -100 109115 -84 109149
rect 84 109115 100 109149
rect -100 109077 100 109115
rect -100 107839 100 107877
rect -100 107805 -84 107839
rect 84 107805 100 107839
rect -100 107789 100 107805
rect -100 107731 100 107747
rect -100 107697 -84 107731
rect 84 107697 100 107731
rect -100 107659 100 107697
rect -100 106421 100 106459
rect -100 106387 -84 106421
rect 84 106387 100 106421
rect -100 106371 100 106387
rect -100 106313 100 106329
rect -100 106279 -84 106313
rect 84 106279 100 106313
rect -100 106241 100 106279
rect -100 105003 100 105041
rect -100 104969 -84 105003
rect 84 104969 100 105003
rect -100 104953 100 104969
rect -100 104895 100 104911
rect -100 104861 -84 104895
rect 84 104861 100 104895
rect -100 104823 100 104861
rect -100 103585 100 103623
rect -100 103551 -84 103585
rect 84 103551 100 103585
rect -100 103535 100 103551
rect -100 103477 100 103493
rect -100 103443 -84 103477
rect 84 103443 100 103477
rect -100 103405 100 103443
rect -100 102167 100 102205
rect -100 102133 -84 102167
rect 84 102133 100 102167
rect -100 102117 100 102133
rect -100 102059 100 102075
rect -100 102025 -84 102059
rect 84 102025 100 102059
rect -100 101987 100 102025
rect -100 100749 100 100787
rect -100 100715 -84 100749
rect 84 100715 100 100749
rect -100 100699 100 100715
rect -100 100641 100 100657
rect -100 100607 -84 100641
rect 84 100607 100 100641
rect -100 100569 100 100607
rect -100 99331 100 99369
rect -100 99297 -84 99331
rect 84 99297 100 99331
rect -100 99281 100 99297
rect -100 99223 100 99239
rect -100 99189 -84 99223
rect 84 99189 100 99223
rect -100 99151 100 99189
rect -100 97913 100 97951
rect -100 97879 -84 97913
rect 84 97879 100 97913
rect -100 97863 100 97879
rect -100 97805 100 97821
rect -100 97771 -84 97805
rect 84 97771 100 97805
rect -100 97733 100 97771
rect -100 96495 100 96533
rect -100 96461 -84 96495
rect 84 96461 100 96495
rect -100 96445 100 96461
rect -100 96387 100 96403
rect -100 96353 -84 96387
rect 84 96353 100 96387
rect -100 96315 100 96353
rect -100 95077 100 95115
rect -100 95043 -84 95077
rect 84 95043 100 95077
rect -100 95027 100 95043
rect -100 94969 100 94985
rect -100 94935 -84 94969
rect 84 94935 100 94969
rect -100 94897 100 94935
rect -100 93659 100 93697
rect -100 93625 -84 93659
rect 84 93625 100 93659
rect -100 93609 100 93625
rect -100 93551 100 93567
rect -100 93517 -84 93551
rect 84 93517 100 93551
rect -100 93479 100 93517
rect -100 92241 100 92279
rect -100 92207 -84 92241
rect 84 92207 100 92241
rect -100 92191 100 92207
rect -100 92133 100 92149
rect -100 92099 -84 92133
rect 84 92099 100 92133
rect -100 92061 100 92099
rect -100 90823 100 90861
rect -100 90789 -84 90823
rect 84 90789 100 90823
rect -100 90773 100 90789
rect -100 90715 100 90731
rect -100 90681 -84 90715
rect 84 90681 100 90715
rect -100 90643 100 90681
rect -100 89405 100 89443
rect -100 89371 -84 89405
rect 84 89371 100 89405
rect -100 89355 100 89371
rect -100 89297 100 89313
rect -100 89263 -84 89297
rect 84 89263 100 89297
rect -100 89225 100 89263
rect -100 87987 100 88025
rect -100 87953 -84 87987
rect 84 87953 100 87987
rect -100 87937 100 87953
rect -100 87879 100 87895
rect -100 87845 -84 87879
rect 84 87845 100 87879
rect -100 87807 100 87845
rect -100 86569 100 86607
rect -100 86535 -84 86569
rect 84 86535 100 86569
rect -100 86519 100 86535
rect -100 86461 100 86477
rect -100 86427 -84 86461
rect 84 86427 100 86461
rect -100 86389 100 86427
rect -100 85151 100 85189
rect -100 85117 -84 85151
rect 84 85117 100 85151
rect -100 85101 100 85117
rect -100 85043 100 85059
rect -100 85009 -84 85043
rect 84 85009 100 85043
rect -100 84971 100 85009
rect -100 83733 100 83771
rect -100 83699 -84 83733
rect 84 83699 100 83733
rect -100 83683 100 83699
rect -100 83625 100 83641
rect -100 83591 -84 83625
rect 84 83591 100 83625
rect -100 83553 100 83591
rect -100 82315 100 82353
rect -100 82281 -84 82315
rect 84 82281 100 82315
rect -100 82265 100 82281
rect -100 82207 100 82223
rect -100 82173 -84 82207
rect 84 82173 100 82207
rect -100 82135 100 82173
rect -100 80897 100 80935
rect -100 80863 -84 80897
rect 84 80863 100 80897
rect -100 80847 100 80863
rect -100 80789 100 80805
rect -100 80755 -84 80789
rect 84 80755 100 80789
rect -100 80717 100 80755
rect -100 79479 100 79517
rect -100 79445 -84 79479
rect 84 79445 100 79479
rect -100 79429 100 79445
rect -100 79371 100 79387
rect -100 79337 -84 79371
rect 84 79337 100 79371
rect -100 79299 100 79337
rect -100 78061 100 78099
rect -100 78027 -84 78061
rect 84 78027 100 78061
rect -100 78011 100 78027
rect -100 77953 100 77969
rect -100 77919 -84 77953
rect 84 77919 100 77953
rect -100 77881 100 77919
rect -100 76643 100 76681
rect -100 76609 -84 76643
rect 84 76609 100 76643
rect -100 76593 100 76609
rect -100 76535 100 76551
rect -100 76501 -84 76535
rect 84 76501 100 76535
rect -100 76463 100 76501
rect -100 75225 100 75263
rect -100 75191 -84 75225
rect 84 75191 100 75225
rect -100 75175 100 75191
rect -100 75117 100 75133
rect -100 75083 -84 75117
rect 84 75083 100 75117
rect -100 75045 100 75083
rect -100 73807 100 73845
rect -100 73773 -84 73807
rect 84 73773 100 73807
rect -100 73757 100 73773
rect -100 73699 100 73715
rect -100 73665 -84 73699
rect 84 73665 100 73699
rect -100 73627 100 73665
rect -100 72389 100 72427
rect -100 72355 -84 72389
rect 84 72355 100 72389
rect -100 72339 100 72355
rect -100 72281 100 72297
rect -100 72247 -84 72281
rect 84 72247 100 72281
rect -100 72209 100 72247
rect -100 70971 100 71009
rect -100 70937 -84 70971
rect 84 70937 100 70971
rect -100 70921 100 70937
rect -100 70863 100 70879
rect -100 70829 -84 70863
rect 84 70829 100 70863
rect -100 70791 100 70829
rect -100 69553 100 69591
rect -100 69519 -84 69553
rect 84 69519 100 69553
rect -100 69503 100 69519
rect -100 69445 100 69461
rect -100 69411 -84 69445
rect 84 69411 100 69445
rect -100 69373 100 69411
rect -100 68135 100 68173
rect -100 68101 -84 68135
rect 84 68101 100 68135
rect -100 68085 100 68101
rect -100 68027 100 68043
rect -100 67993 -84 68027
rect 84 67993 100 68027
rect -100 67955 100 67993
rect -100 66717 100 66755
rect -100 66683 -84 66717
rect 84 66683 100 66717
rect -100 66667 100 66683
rect -100 66609 100 66625
rect -100 66575 -84 66609
rect 84 66575 100 66609
rect -100 66537 100 66575
rect -100 65299 100 65337
rect -100 65265 -84 65299
rect 84 65265 100 65299
rect -100 65249 100 65265
rect -100 65191 100 65207
rect -100 65157 -84 65191
rect 84 65157 100 65191
rect -100 65119 100 65157
rect -100 63881 100 63919
rect -100 63847 -84 63881
rect 84 63847 100 63881
rect -100 63831 100 63847
rect -100 63773 100 63789
rect -100 63739 -84 63773
rect 84 63739 100 63773
rect -100 63701 100 63739
rect -100 62463 100 62501
rect -100 62429 -84 62463
rect 84 62429 100 62463
rect -100 62413 100 62429
rect -100 62355 100 62371
rect -100 62321 -84 62355
rect 84 62321 100 62355
rect -100 62283 100 62321
rect -100 61045 100 61083
rect -100 61011 -84 61045
rect 84 61011 100 61045
rect -100 60995 100 61011
rect -100 60937 100 60953
rect -100 60903 -84 60937
rect 84 60903 100 60937
rect -100 60865 100 60903
rect -100 59627 100 59665
rect -100 59593 -84 59627
rect 84 59593 100 59627
rect -100 59577 100 59593
rect -100 59519 100 59535
rect -100 59485 -84 59519
rect 84 59485 100 59519
rect -100 59447 100 59485
rect -100 58209 100 58247
rect -100 58175 -84 58209
rect 84 58175 100 58209
rect -100 58159 100 58175
rect -100 58101 100 58117
rect -100 58067 -84 58101
rect 84 58067 100 58101
rect -100 58029 100 58067
rect -100 56791 100 56829
rect -100 56757 -84 56791
rect 84 56757 100 56791
rect -100 56741 100 56757
rect -100 56683 100 56699
rect -100 56649 -84 56683
rect 84 56649 100 56683
rect -100 56611 100 56649
rect -100 55373 100 55411
rect -100 55339 -84 55373
rect 84 55339 100 55373
rect -100 55323 100 55339
rect -100 55265 100 55281
rect -100 55231 -84 55265
rect 84 55231 100 55265
rect -100 55193 100 55231
rect -100 53955 100 53993
rect -100 53921 -84 53955
rect 84 53921 100 53955
rect -100 53905 100 53921
rect -100 53847 100 53863
rect -100 53813 -84 53847
rect 84 53813 100 53847
rect -100 53775 100 53813
rect -100 52537 100 52575
rect -100 52503 -84 52537
rect 84 52503 100 52537
rect -100 52487 100 52503
rect -100 52429 100 52445
rect -100 52395 -84 52429
rect 84 52395 100 52429
rect -100 52357 100 52395
rect -100 51119 100 51157
rect -100 51085 -84 51119
rect 84 51085 100 51119
rect -100 51069 100 51085
rect -100 51011 100 51027
rect -100 50977 -84 51011
rect 84 50977 100 51011
rect -100 50939 100 50977
rect -100 49701 100 49739
rect -100 49667 -84 49701
rect 84 49667 100 49701
rect -100 49651 100 49667
rect -100 49593 100 49609
rect -100 49559 -84 49593
rect 84 49559 100 49593
rect -100 49521 100 49559
rect -100 48283 100 48321
rect -100 48249 -84 48283
rect 84 48249 100 48283
rect -100 48233 100 48249
rect -100 48175 100 48191
rect -100 48141 -84 48175
rect 84 48141 100 48175
rect -100 48103 100 48141
rect -100 46865 100 46903
rect -100 46831 -84 46865
rect 84 46831 100 46865
rect -100 46815 100 46831
rect -100 46757 100 46773
rect -100 46723 -84 46757
rect 84 46723 100 46757
rect -100 46685 100 46723
rect -100 45447 100 45485
rect -100 45413 -84 45447
rect 84 45413 100 45447
rect -100 45397 100 45413
rect -100 45339 100 45355
rect -100 45305 -84 45339
rect 84 45305 100 45339
rect -100 45267 100 45305
rect -100 44029 100 44067
rect -100 43995 -84 44029
rect 84 43995 100 44029
rect -100 43979 100 43995
rect -100 43921 100 43937
rect -100 43887 -84 43921
rect 84 43887 100 43921
rect -100 43849 100 43887
rect -100 42611 100 42649
rect -100 42577 -84 42611
rect 84 42577 100 42611
rect -100 42561 100 42577
rect -100 42503 100 42519
rect -100 42469 -84 42503
rect 84 42469 100 42503
rect -100 42431 100 42469
rect -100 41193 100 41231
rect -100 41159 -84 41193
rect 84 41159 100 41193
rect -100 41143 100 41159
rect -100 41085 100 41101
rect -100 41051 -84 41085
rect 84 41051 100 41085
rect -100 41013 100 41051
rect -100 39775 100 39813
rect -100 39741 -84 39775
rect 84 39741 100 39775
rect -100 39725 100 39741
rect -100 39667 100 39683
rect -100 39633 -84 39667
rect 84 39633 100 39667
rect -100 39595 100 39633
rect -100 38357 100 38395
rect -100 38323 -84 38357
rect 84 38323 100 38357
rect -100 38307 100 38323
rect -100 38249 100 38265
rect -100 38215 -84 38249
rect 84 38215 100 38249
rect -100 38177 100 38215
rect -100 36939 100 36977
rect -100 36905 -84 36939
rect 84 36905 100 36939
rect -100 36889 100 36905
rect -100 36831 100 36847
rect -100 36797 -84 36831
rect 84 36797 100 36831
rect -100 36759 100 36797
rect -100 35521 100 35559
rect -100 35487 -84 35521
rect 84 35487 100 35521
rect -100 35471 100 35487
rect -100 35413 100 35429
rect -100 35379 -84 35413
rect 84 35379 100 35413
rect -100 35341 100 35379
rect -100 34103 100 34141
rect -100 34069 -84 34103
rect 84 34069 100 34103
rect -100 34053 100 34069
rect -100 33995 100 34011
rect -100 33961 -84 33995
rect 84 33961 100 33995
rect -100 33923 100 33961
rect -100 32685 100 32723
rect -100 32651 -84 32685
rect 84 32651 100 32685
rect -100 32635 100 32651
rect -100 32577 100 32593
rect -100 32543 -84 32577
rect 84 32543 100 32577
rect -100 32505 100 32543
rect -100 31267 100 31305
rect -100 31233 -84 31267
rect 84 31233 100 31267
rect -100 31217 100 31233
rect -100 31159 100 31175
rect -100 31125 -84 31159
rect 84 31125 100 31159
rect -100 31087 100 31125
rect -100 29849 100 29887
rect -100 29815 -84 29849
rect 84 29815 100 29849
rect -100 29799 100 29815
rect -100 29741 100 29757
rect -100 29707 -84 29741
rect 84 29707 100 29741
rect -100 29669 100 29707
rect -100 28431 100 28469
rect -100 28397 -84 28431
rect 84 28397 100 28431
rect -100 28381 100 28397
rect -100 28323 100 28339
rect -100 28289 -84 28323
rect 84 28289 100 28323
rect -100 28251 100 28289
rect -100 27013 100 27051
rect -100 26979 -84 27013
rect 84 26979 100 27013
rect -100 26963 100 26979
rect -100 26905 100 26921
rect -100 26871 -84 26905
rect 84 26871 100 26905
rect -100 26833 100 26871
rect -100 25595 100 25633
rect -100 25561 -84 25595
rect 84 25561 100 25595
rect -100 25545 100 25561
rect -100 25487 100 25503
rect -100 25453 -84 25487
rect 84 25453 100 25487
rect -100 25415 100 25453
rect -100 24177 100 24215
rect -100 24143 -84 24177
rect 84 24143 100 24177
rect -100 24127 100 24143
rect -100 24069 100 24085
rect -100 24035 -84 24069
rect 84 24035 100 24069
rect -100 23997 100 24035
rect -100 22759 100 22797
rect -100 22725 -84 22759
rect 84 22725 100 22759
rect -100 22709 100 22725
rect -100 22651 100 22667
rect -100 22617 -84 22651
rect 84 22617 100 22651
rect -100 22579 100 22617
rect -100 21341 100 21379
rect -100 21307 -84 21341
rect 84 21307 100 21341
rect -100 21291 100 21307
rect -100 21233 100 21249
rect -100 21199 -84 21233
rect 84 21199 100 21233
rect -100 21161 100 21199
rect -100 19923 100 19961
rect -100 19889 -84 19923
rect 84 19889 100 19923
rect -100 19873 100 19889
rect -100 19815 100 19831
rect -100 19781 -84 19815
rect 84 19781 100 19815
rect -100 19743 100 19781
rect -100 18505 100 18543
rect -100 18471 -84 18505
rect 84 18471 100 18505
rect -100 18455 100 18471
rect -100 18397 100 18413
rect -100 18363 -84 18397
rect 84 18363 100 18397
rect -100 18325 100 18363
rect -100 17087 100 17125
rect -100 17053 -84 17087
rect 84 17053 100 17087
rect -100 17037 100 17053
rect -100 16979 100 16995
rect -100 16945 -84 16979
rect 84 16945 100 16979
rect -100 16907 100 16945
rect -100 15669 100 15707
rect -100 15635 -84 15669
rect 84 15635 100 15669
rect -100 15619 100 15635
rect -100 15561 100 15577
rect -100 15527 -84 15561
rect 84 15527 100 15561
rect -100 15489 100 15527
rect -100 14251 100 14289
rect -100 14217 -84 14251
rect 84 14217 100 14251
rect -100 14201 100 14217
rect -100 14143 100 14159
rect -100 14109 -84 14143
rect 84 14109 100 14143
rect -100 14071 100 14109
rect -100 12833 100 12871
rect -100 12799 -84 12833
rect 84 12799 100 12833
rect -100 12783 100 12799
rect -100 12725 100 12741
rect -100 12691 -84 12725
rect 84 12691 100 12725
rect -100 12653 100 12691
rect -100 11415 100 11453
rect -100 11381 -84 11415
rect 84 11381 100 11415
rect -100 11365 100 11381
rect -100 11307 100 11323
rect -100 11273 -84 11307
rect 84 11273 100 11307
rect -100 11235 100 11273
rect -100 9997 100 10035
rect -100 9963 -84 9997
rect 84 9963 100 9997
rect -100 9947 100 9963
rect -100 9889 100 9905
rect -100 9855 -84 9889
rect 84 9855 100 9889
rect -100 9817 100 9855
rect -100 8579 100 8617
rect -100 8545 -84 8579
rect 84 8545 100 8579
rect -100 8529 100 8545
rect -100 8471 100 8487
rect -100 8437 -84 8471
rect 84 8437 100 8471
rect -100 8399 100 8437
rect -100 7161 100 7199
rect -100 7127 -84 7161
rect 84 7127 100 7161
rect -100 7111 100 7127
rect -100 7053 100 7069
rect -100 7019 -84 7053
rect 84 7019 100 7053
rect -100 6981 100 7019
rect -100 5743 100 5781
rect -100 5709 -84 5743
rect 84 5709 100 5743
rect -100 5693 100 5709
rect -100 5635 100 5651
rect -100 5601 -84 5635
rect 84 5601 100 5635
rect -100 5563 100 5601
rect -100 4325 100 4363
rect -100 4291 -84 4325
rect 84 4291 100 4325
rect -100 4275 100 4291
rect -100 4217 100 4233
rect -100 4183 -84 4217
rect 84 4183 100 4217
rect -100 4145 100 4183
rect -100 2907 100 2945
rect -100 2873 -84 2907
rect 84 2873 100 2907
rect -100 2857 100 2873
rect -100 2799 100 2815
rect -100 2765 -84 2799
rect 84 2765 100 2799
rect -100 2727 100 2765
rect -100 1489 100 1527
rect -100 1455 -84 1489
rect 84 1455 100 1489
rect -100 1439 100 1455
rect -100 1381 100 1397
rect -100 1347 -84 1381
rect 84 1347 100 1381
rect -100 1309 100 1347
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -1347 100 -1309
rect -100 -1381 -84 -1347
rect 84 -1381 100 -1347
rect -100 -1397 100 -1381
rect -100 -1455 100 -1439
rect -100 -1489 -84 -1455
rect 84 -1489 100 -1455
rect -100 -1527 100 -1489
rect -100 -2765 100 -2727
rect -100 -2799 -84 -2765
rect 84 -2799 100 -2765
rect -100 -2815 100 -2799
rect -100 -2873 100 -2857
rect -100 -2907 -84 -2873
rect 84 -2907 100 -2873
rect -100 -2945 100 -2907
rect -100 -4183 100 -4145
rect -100 -4217 -84 -4183
rect 84 -4217 100 -4183
rect -100 -4233 100 -4217
rect -100 -4291 100 -4275
rect -100 -4325 -84 -4291
rect 84 -4325 100 -4291
rect -100 -4363 100 -4325
rect -100 -5601 100 -5563
rect -100 -5635 -84 -5601
rect 84 -5635 100 -5601
rect -100 -5651 100 -5635
rect -100 -5709 100 -5693
rect -100 -5743 -84 -5709
rect 84 -5743 100 -5709
rect -100 -5781 100 -5743
rect -100 -7019 100 -6981
rect -100 -7053 -84 -7019
rect 84 -7053 100 -7019
rect -100 -7069 100 -7053
rect -100 -7127 100 -7111
rect -100 -7161 -84 -7127
rect 84 -7161 100 -7127
rect -100 -7199 100 -7161
rect -100 -8437 100 -8399
rect -100 -8471 -84 -8437
rect 84 -8471 100 -8437
rect -100 -8487 100 -8471
rect -100 -8545 100 -8529
rect -100 -8579 -84 -8545
rect 84 -8579 100 -8545
rect -100 -8617 100 -8579
rect -100 -9855 100 -9817
rect -100 -9889 -84 -9855
rect 84 -9889 100 -9855
rect -100 -9905 100 -9889
rect -100 -9963 100 -9947
rect -100 -9997 -84 -9963
rect 84 -9997 100 -9963
rect -100 -10035 100 -9997
rect -100 -11273 100 -11235
rect -100 -11307 -84 -11273
rect 84 -11307 100 -11273
rect -100 -11323 100 -11307
rect -100 -11381 100 -11365
rect -100 -11415 -84 -11381
rect 84 -11415 100 -11381
rect -100 -11453 100 -11415
rect -100 -12691 100 -12653
rect -100 -12725 -84 -12691
rect 84 -12725 100 -12691
rect -100 -12741 100 -12725
rect -100 -12799 100 -12783
rect -100 -12833 -84 -12799
rect 84 -12833 100 -12799
rect -100 -12871 100 -12833
rect -100 -14109 100 -14071
rect -100 -14143 -84 -14109
rect 84 -14143 100 -14109
rect -100 -14159 100 -14143
rect -100 -14217 100 -14201
rect -100 -14251 -84 -14217
rect 84 -14251 100 -14217
rect -100 -14289 100 -14251
rect -100 -15527 100 -15489
rect -100 -15561 -84 -15527
rect 84 -15561 100 -15527
rect -100 -15577 100 -15561
rect -100 -15635 100 -15619
rect -100 -15669 -84 -15635
rect 84 -15669 100 -15635
rect -100 -15707 100 -15669
rect -100 -16945 100 -16907
rect -100 -16979 -84 -16945
rect 84 -16979 100 -16945
rect -100 -16995 100 -16979
rect -100 -17053 100 -17037
rect -100 -17087 -84 -17053
rect 84 -17087 100 -17053
rect -100 -17125 100 -17087
rect -100 -18363 100 -18325
rect -100 -18397 -84 -18363
rect 84 -18397 100 -18363
rect -100 -18413 100 -18397
rect -100 -18471 100 -18455
rect -100 -18505 -84 -18471
rect 84 -18505 100 -18471
rect -100 -18543 100 -18505
rect -100 -19781 100 -19743
rect -100 -19815 -84 -19781
rect 84 -19815 100 -19781
rect -100 -19831 100 -19815
rect -100 -19889 100 -19873
rect -100 -19923 -84 -19889
rect 84 -19923 100 -19889
rect -100 -19961 100 -19923
rect -100 -21199 100 -21161
rect -100 -21233 -84 -21199
rect 84 -21233 100 -21199
rect -100 -21249 100 -21233
rect -100 -21307 100 -21291
rect -100 -21341 -84 -21307
rect 84 -21341 100 -21307
rect -100 -21379 100 -21341
rect -100 -22617 100 -22579
rect -100 -22651 -84 -22617
rect 84 -22651 100 -22617
rect -100 -22667 100 -22651
rect -100 -22725 100 -22709
rect -100 -22759 -84 -22725
rect 84 -22759 100 -22725
rect -100 -22797 100 -22759
rect -100 -24035 100 -23997
rect -100 -24069 -84 -24035
rect 84 -24069 100 -24035
rect -100 -24085 100 -24069
rect -100 -24143 100 -24127
rect -100 -24177 -84 -24143
rect 84 -24177 100 -24143
rect -100 -24215 100 -24177
rect -100 -25453 100 -25415
rect -100 -25487 -84 -25453
rect 84 -25487 100 -25453
rect -100 -25503 100 -25487
rect -100 -25561 100 -25545
rect -100 -25595 -84 -25561
rect 84 -25595 100 -25561
rect -100 -25633 100 -25595
rect -100 -26871 100 -26833
rect -100 -26905 -84 -26871
rect 84 -26905 100 -26871
rect -100 -26921 100 -26905
rect -100 -26979 100 -26963
rect -100 -27013 -84 -26979
rect 84 -27013 100 -26979
rect -100 -27051 100 -27013
rect -100 -28289 100 -28251
rect -100 -28323 -84 -28289
rect 84 -28323 100 -28289
rect -100 -28339 100 -28323
rect -100 -28397 100 -28381
rect -100 -28431 -84 -28397
rect 84 -28431 100 -28397
rect -100 -28469 100 -28431
rect -100 -29707 100 -29669
rect -100 -29741 -84 -29707
rect 84 -29741 100 -29707
rect -100 -29757 100 -29741
rect -100 -29815 100 -29799
rect -100 -29849 -84 -29815
rect 84 -29849 100 -29815
rect -100 -29887 100 -29849
rect -100 -31125 100 -31087
rect -100 -31159 -84 -31125
rect 84 -31159 100 -31125
rect -100 -31175 100 -31159
rect -100 -31233 100 -31217
rect -100 -31267 -84 -31233
rect 84 -31267 100 -31233
rect -100 -31305 100 -31267
rect -100 -32543 100 -32505
rect -100 -32577 -84 -32543
rect 84 -32577 100 -32543
rect -100 -32593 100 -32577
rect -100 -32651 100 -32635
rect -100 -32685 -84 -32651
rect 84 -32685 100 -32651
rect -100 -32723 100 -32685
rect -100 -33961 100 -33923
rect -100 -33995 -84 -33961
rect 84 -33995 100 -33961
rect -100 -34011 100 -33995
rect -100 -34069 100 -34053
rect -100 -34103 -84 -34069
rect 84 -34103 100 -34069
rect -100 -34141 100 -34103
rect -100 -35379 100 -35341
rect -100 -35413 -84 -35379
rect 84 -35413 100 -35379
rect -100 -35429 100 -35413
rect -100 -35487 100 -35471
rect -100 -35521 -84 -35487
rect 84 -35521 100 -35487
rect -100 -35559 100 -35521
rect -100 -36797 100 -36759
rect -100 -36831 -84 -36797
rect 84 -36831 100 -36797
rect -100 -36847 100 -36831
rect -100 -36905 100 -36889
rect -100 -36939 -84 -36905
rect 84 -36939 100 -36905
rect -100 -36977 100 -36939
rect -100 -38215 100 -38177
rect -100 -38249 -84 -38215
rect 84 -38249 100 -38215
rect -100 -38265 100 -38249
rect -100 -38323 100 -38307
rect -100 -38357 -84 -38323
rect 84 -38357 100 -38323
rect -100 -38395 100 -38357
rect -100 -39633 100 -39595
rect -100 -39667 -84 -39633
rect 84 -39667 100 -39633
rect -100 -39683 100 -39667
rect -100 -39741 100 -39725
rect -100 -39775 -84 -39741
rect 84 -39775 100 -39741
rect -100 -39813 100 -39775
rect -100 -41051 100 -41013
rect -100 -41085 -84 -41051
rect 84 -41085 100 -41051
rect -100 -41101 100 -41085
rect -100 -41159 100 -41143
rect -100 -41193 -84 -41159
rect 84 -41193 100 -41159
rect -100 -41231 100 -41193
rect -100 -42469 100 -42431
rect -100 -42503 -84 -42469
rect 84 -42503 100 -42469
rect -100 -42519 100 -42503
rect -100 -42577 100 -42561
rect -100 -42611 -84 -42577
rect 84 -42611 100 -42577
rect -100 -42649 100 -42611
rect -100 -43887 100 -43849
rect -100 -43921 -84 -43887
rect 84 -43921 100 -43887
rect -100 -43937 100 -43921
rect -100 -43995 100 -43979
rect -100 -44029 -84 -43995
rect 84 -44029 100 -43995
rect -100 -44067 100 -44029
rect -100 -45305 100 -45267
rect -100 -45339 -84 -45305
rect 84 -45339 100 -45305
rect -100 -45355 100 -45339
rect -100 -45413 100 -45397
rect -100 -45447 -84 -45413
rect 84 -45447 100 -45413
rect -100 -45485 100 -45447
rect -100 -46723 100 -46685
rect -100 -46757 -84 -46723
rect 84 -46757 100 -46723
rect -100 -46773 100 -46757
rect -100 -46831 100 -46815
rect -100 -46865 -84 -46831
rect 84 -46865 100 -46831
rect -100 -46903 100 -46865
rect -100 -48141 100 -48103
rect -100 -48175 -84 -48141
rect 84 -48175 100 -48141
rect -100 -48191 100 -48175
rect -100 -48249 100 -48233
rect -100 -48283 -84 -48249
rect 84 -48283 100 -48249
rect -100 -48321 100 -48283
rect -100 -49559 100 -49521
rect -100 -49593 -84 -49559
rect 84 -49593 100 -49559
rect -100 -49609 100 -49593
rect -100 -49667 100 -49651
rect -100 -49701 -84 -49667
rect 84 -49701 100 -49667
rect -100 -49739 100 -49701
rect -100 -50977 100 -50939
rect -100 -51011 -84 -50977
rect 84 -51011 100 -50977
rect -100 -51027 100 -51011
rect -100 -51085 100 -51069
rect -100 -51119 -84 -51085
rect 84 -51119 100 -51085
rect -100 -51157 100 -51119
rect -100 -52395 100 -52357
rect -100 -52429 -84 -52395
rect 84 -52429 100 -52395
rect -100 -52445 100 -52429
rect -100 -52503 100 -52487
rect -100 -52537 -84 -52503
rect 84 -52537 100 -52503
rect -100 -52575 100 -52537
rect -100 -53813 100 -53775
rect -100 -53847 -84 -53813
rect 84 -53847 100 -53813
rect -100 -53863 100 -53847
rect -100 -53921 100 -53905
rect -100 -53955 -84 -53921
rect 84 -53955 100 -53921
rect -100 -53993 100 -53955
rect -100 -55231 100 -55193
rect -100 -55265 -84 -55231
rect 84 -55265 100 -55231
rect -100 -55281 100 -55265
rect -100 -55339 100 -55323
rect -100 -55373 -84 -55339
rect 84 -55373 100 -55339
rect -100 -55411 100 -55373
rect -100 -56649 100 -56611
rect -100 -56683 -84 -56649
rect 84 -56683 100 -56649
rect -100 -56699 100 -56683
rect -100 -56757 100 -56741
rect -100 -56791 -84 -56757
rect 84 -56791 100 -56757
rect -100 -56829 100 -56791
rect -100 -58067 100 -58029
rect -100 -58101 -84 -58067
rect 84 -58101 100 -58067
rect -100 -58117 100 -58101
rect -100 -58175 100 -58159
rect -100 -58209 -84 -58175
rect 84 -58209 100 -58175
rect -100 -58247 100 -58209
rect -100 -59485 100 -59447
rect -100 -59519 -84 -59485
rect 84 -59519 100 -59485
rect -100 -59535 100 -59519
rect -100 -59593 100 -59577
rect -100 -59627 -84 -59593
rect 84 -59627 100 -59593
rect -100 -59665 100 -59627
rect -100 -60903 100 -60865
rect -100 -60937 -84 -60903
rect 84 -60937 100 -60903
rect -100 -60953 100 -60937
rect -100 -61011 100 -60995
rect -100 -61045 -84 -61011
rect 84 -61045 100 -61011
rect -100 -61083 100 -61045
rect -100 -62321 100 -62283
rect -100 -62355 -84 -62321
rect 84 -62355 100 -62321
rect -100 -62371 100 -62355
rect -100 -62429 100 -62413
rect -100 -62463 -84 -62429
rect 84 -62463 100 -62429
rect -100 -62501 100 -62463
rect -100 -63739 100 -63701
rect -100 -63773 -84 -63739
rect 84 -63773 100 -63739
rect -100 -63789 100 -63773
rect -100 -63847 100 -63831
rect -100 -63881 -84 -63847
rect 84 -63881 100 -63847
rect -100 -63919 100 -63881
rect -100 -65157 100 -65119
rect -100 -65191 -84 -65157
rect 84 -65191 100 -65157
rect -100 -65207 100 -65191
rect -100 -65265 100 -65249
rect -100 -65299 -84 -65265
rect 84 -65299 100 -65265
rect -100 -65337 100 -65299
rect -100 -66575 100 -66537
rect -100 -66609 -84 -66575
rect 84 -66609 100 -66575
rect -100 -66625 100 -66609
rect -100 -66683 100 -66667
rect -100 -66717 -84 -66683
rect 84 -66717 100 -66683
rect -100 -66755 100 -66717
rect -100 -67993 100 -67955
rect -100 -68027 -84 -67993
rect 84 -68027 100 -67993
rect -100 -68043 100 -68027
rect -100 -68101 100 -68085
rect -100 -68135 -84 -68101
rect 84 -68135 100 -68101
rect -100 -68173 100 -68135
rect -100 -69411 100 -69373
rect -100 -69445 -84 -69411
rect 84 -69445 100 -69411
rect -100 -69461 100 -69445
rect -100 -69519 100 -69503
rect -100 -69553 -84 -69519
rect 84 -69553 100 -69519
rect -100 -69591 100 -69553
rect -100 -70829 100 -70791
rect -100 -70863 -84 -70829
rect 84 -70863 100 -70829
rect -100 -70879 100 -70863
rect -100 -70937 100 -70921
rect -100 -70971 -84 -70937
rect 84 -70971 100 -70937
rect -100 -71009 100 -70971
rect -100 -72247 100 -72209
rect -100 -72281 -84 -72247
rect 84 -72281 100 -72247
rect -100 -72297 100 -72281
rect -100 -72355 100 -72339
rect -100 -72389 -84 -72355
rect 84 -72389 100 -72355
rect -100 -72427 100 -72389
rect -100 -73665 100 -73627
rect -100 -73699 -84 -73665
rect 84 -73699 100 -73665
rect -100 -73715 100 -73699
rect -100 -73773 100 -73757
rect -100 -73807 -84 -73773
rect 84 -73807 100 -73773
rect -100 -73845 100 -73807
rect -100 -75083 100 -75045
rect -100 -75117 -84 -75083
rect 84 -75117 100 -75083
rect -100 -75133 100 -75117
rect -100 -75191 100 -75175
rect -100 -75225 -84 -75191
rect 84 -75225 100 -75191
rect -100 -75263 100 -75225
rect -100 -76501 100 -76463
rect -100 -76535 -84 -76501
rect 84 -76535 100 -76501
rect -100 -76551 100 -76535
rect -100 -76609 100 -76593
rect -100 -76643 -84 -76609
rect 84 -76643 100 -76609
rect -100 -76681 100 -76643
rect -100 -77919 100 -77881
rect -100 -77953 -84 -77919
rect 84 -77953 100 -77919
rect -100 -77969 100 -77953
rect -100 -78027 100 -78011
rect -100 -78061 -84 -78027
rect 84 -78061 100 -78027
rect -100 -78099 100 -78061
rect -100 -79337 100 -79299
rect -100 -79371 -84 -79337
rect 84 -79371 100 -79337
rect -100 -79387 100 -79371
rect -100 -79445 100 -79429
rect -100 -79479 -84 -79445
rect 84 -79479 100 -79445
rect -100 -79517 100 -79479
rect -100 -80755 100 -80717
rect -100 -80789 -84 -80755
rect 84 -80789 100 -80755
rect -100 -80805 100 -80789
rect -100 -80863 100 -80847
rect -100 -80897 -84 -80863
rect 84 -80897 100 -80863
rect -100 -80935 100 -80897
rect -100 -82173 100 -82135
rect -100 -82207 -84 -82173
rect 84 -82207 100 -82173
rect -100 -82223 100 -82207
rect -100 -82281 100 -82265
rect -100 -82315 -84 -82281
rect 84 -82315 100 -82281
rect -100 -82353 100 -82315
rect -100 -83591 100 -83553
rect -100 -83625 -84 -83591
rect 84 -83625 100 -83591
rect -100 -83641 100 -83625
rect -100 -83699 100 -83683
rect -100 -83733 -84 -83699
rect 84 -83733 100 -83699
rect -100 -83771 100 -83733
rect -100 -85009 100 -84971
rect -100 -85043 -84 -85009
rect 84 -85043 100 -85009
rect -100 -85059 100 -85043
rect -100 -85117 100 -85101
rect -100 -85151 -84 -85117
rect 84 -85151 100 -85117
rect -100 -85189 100 -85151
rect -100 -86427 100 -86389
rect -100 -86461 -84 -86427
rect 84 -86461 100 -86427
rect -100 -86477 100 -86461
rect -100 -86535 100 -86519
rect -100 -86569 -84 -86535
rect 84 -86569 100 -86535
rect -100 -86607 100 -86569
rect -100 -87845 100 -87807
rect -100 -87879 -84 -87845
rect 84 -87879 100 -87845
rect -100 -87895 100 -87879
rect -100 -87953 100 -87937
rect -100 -87987 -84 -87953
rect 84 -87987 100 -87953
rect -100 -88025 100 -87987
rect -100 -89263 100 -89225
rect -100 -89297 -84 -89263
rect 84 -89297 100 -89263
rect -100 -89313 100 -89297
rect -100 -89371 100 -89355
rect -100 -89405 -84 -89371
rect 84 -89405 100 -89371
rect -100 -89443 100 -89405
rect -100 -90681 100 -90643
rect -100 -90715 -84 -90681
rect 84 -90715 100 -90681
rect -100 -90731 100 -90715
rect -100 -90789 100 -90773
rect -100 -90823 -84 -90789
rect 84 -90823 100 -90789
rect -100 -90861 100 -90823
rect -100 -92099 100 -92061
rect -100 -92133 -84 -92099
rect 84 -92133 100 -92099
rect -100 -92149 100 -92133
rect -100 -92207 100 -92191
rect -100 -92241 -84 -92207
rect 84 -92241 100 -92207
rect -100 -92279 100 -92241
rect -100 -93517 100 -93479
rect -100 -93551 -84 -93517
rect 84 -93551 100 -93517
rect -100 -93567 100 -93551
rect -100 -93625 100 -93609
rect -100 -93659 -84 -93625
rect 84 -93659 100 -93625
rect -100 -93697 100 -93659
rect -100 -94935 100 -94897
rect -100 -94969 -84 -94935
rect 84 -94969 100 -94935
rect -100 -94985 100 -94969
rect -100 -95043 100 -95027
rect -100 -95077 -84 -95043
rect 84 -95077 100 -95043
rect -100 -95115 100 -95077
rect -100 -96353 100 -96315
rect -100 -96387 -84 -96353
rect 84 -96387 100 -96353
rect -100 -96403 100 -96387
rect -100 -96461 100 -96445
rect -100 -96495 -84 -96461
rect 84 -96495 100 -96461
rect -100 -96533 100 -96495
rect -100 -97771 100 -97733
rect -100 -97805 -84 -97771
rect 84 -97805 100 -97771
rect -100 -97821 100 -97805
rect -100 -97879 100 -97863
rect -100 -97913 -84 -97879
rect 84 -97913 100 -97879
rect -100 -97951 100 -97913
rect -100 -99189 100 -99151
rect -100 -99223 -84 -99189
rect 84 -99223 100 -99189
rect -100 -99239 100 -99223
rect -100 -99297 100 -99281
rect -100 -99331 -84 -99297
rect 84 -99331 100 -99297
rect -100 -99369 100 -99331
rect -100 -100607 100 -100569
rect -100 -100641 -84 -100607
rect 84 -100641 100 -100607
rect -100 -100657 100 -100641
rect -100 -100715 100 -100699
rect -100 -100749 -84 -100715
rect 84 -100749 100 -100715
rect -100 -100787 100 -100749
rect -100 -102025 100 -101987
rect -100 -102059 -84 -102025
rect 84 -102059 100 -102025
rect -100 -102075 100 -102059
rect -100 -102133 100 -102117
rect -100 -102167 -84 -102133
rect 84 -102167 100 -102133
rect -100 -102205 100 -102167
rect -100 -103443 100 -103405
rect -100 -103477 -84 -103443
rect 84 -103477 100 -103443
rect -100 -103493 100 -103477
rect -100 -103551 100 -103535
rect -100 -103585 -84 -103551
rect 84 -103585 100 -103551
rect -100 -103623 100 -103585
rect -100 -104861 100 -104823
rect -100 -104895 -84 -104861
rect 84 -104895 100 -104861
rect -100 -104911 100 -104895
rect -100 -104969 100 -104953
rect -100 -105003 -84 -104969
rect 84 -105003 100 -104969
rect -100 -105041 100 -105003
rect -100 -106279 100 -106241
rect -100 -106313 -84 -106279
rect 84 -106313 100 -106279
rect -100 -106329 100 -106313
rect -100 -106387 100 -106371
rect -100 -106421 -84 -106387
rect 84 -106421 100 -106387
rect -100 -106459 100 -106421
rect -100 -107697 100 -107659
rect -100 -107731 -84 -107697
rect 84 -107731 100 -107697
rect -100 -107747 100 -107731
rect -100 -107805 100 -107789
rect -100 -107839 -84 -107805
rect 84 -107839 100 -107805
rect -100 -107877 100 -107839
rect -100 -109115 100 -109077
rect -100 -109149 -84 -109115
rect 84 -109149 100 -109115
rect -100 -109165 100 -109149
rect -100 -109223 100 -109207
rect -100 -109257 -84 -109223
rect 84 -109257 100 -109223
rect -100 -109295 100 -109257
rect -100 -110533 100 -110495
rect -100 -110567 -84 -110533
rect 84 -110567 100 -110533
rect -100 -110583 100 -110567
rect -100 -110641 100 -110625
rect -100 -110675 -84 -110641
rect 84 -110675 100 -110641
rect -100 -110713 100 -110675
rect -100 -111951 100 -111913
rect -100 -111985 -84 -111951
rect 84 -111985 100 -111951
rect -100 -112001 100 -111985
rect -100 -112059 100 -112043
rect -100 -112093 -84 -112059
rect 84 -112093 100 -112059
rect -100 -112131 100 -112093
rect -100 -113369 100 -113331
rect -100 -113403 -84 -113369
rect 84 -113403 100 -113369
rect -100 -113419 100 -113403
rect -100 -113477 100 -113461
rect -100 -113511 -84 -113477
rect 84 -113511 100 -113477
rect -100 -113549 100 -113511
rect -100 -114787 100 -114749
rect -100 -114821 -84 -114787
rect 84 -114821 100 -114787
rect -100 -114837 100 -114821
rect -100 -114895 100 -114879
rect -100 -114929 -84 -114895
rect 84 -114929 100 -114895
rect -100 -114967 100 -114929
rect -100 -116205 100 -116167
rect -100 -116239 -84 -116205
rect 84 -116239 100 -116205
rect -100 -116255 100 -116239
rect -100 -116313 100 -116297
rect -100 -116347 -84 -116313
rect 84 -116347 100 -116313
rect -100 -116385 100 -116347
rect -100 -117623 100 -117585
rect -100 -117657 -84 -117623
rect 84 -117657 100 -117623
rect -100 -117673 100 -117657
rect -100 -117731 100 -117715
rect -100 -117765 -84 -117731
rect 84 -117765 100 -117731
rect -100 -117803 100 -117765
rect -100 -119041 100 -119003
rect -100 -119075 -84 -119041
rect 84 -119075 100 -119041
rect -100 -119091 100 -119075
rect -100 -119149 100 -119133
rect -100 -119183 -84 -119149
rect 84 -119183 100 -119149
rect -100 -119221 100 -119183
rect -100 -120459 100 -120421
rect -100 -120493 -84 -120459
rect 84 -120493 100 -120459
rect -100 -120509 100 -120493
rect -100 -120567 100 -120551
rect -100 -120601 -84 -120567
rect 84 -120601 100 -120567
rect -100 -120639 100 -120601
rect -100 -121877 100 -121839
rect -100 -121911 -84 -121877
rect 84 -121911 100 -121877
rect -100 -121927 100 -121911
rect -100 -121985 100 -121969
rect -100 -122019 -84 -121985
rect 84 -122019 100 -121985
rect -100 -122057 100 -122019
rect -100 -123295 100 -123257
rect -100 -123329 -84 -123295
rect 84 -123329 100 -123295
rect -100 -123345 100 -123329
rect -100 -123403 100 -123387
rect -100 -123437 -84 -123403
rect 84 -123437 100 -123403
rect -100 -123475 100 -123437
rect -100 -124713 100 -124675
rect -100 -124747 -84 -124713
rect 84 -124747 100 -124713
rect -100 -124763 100 -124747
rect -100 -124821 100 -124805
rect -100 -124855 -84 -124821
rect 84 -124855 100 -124821
rect -100 -124893 100 -124855
rect -100 -126131 100 -126093
rect -100 -126165 -84 -126131
rect 84 -126165 100 -126131
rect -100 -126181 100 -126165
rect -100 -126239 100 -126223
rect -100 -126273 -84 -126239
rect 84 -126273 100 -126239
rect -100 -126311 100 -126273
rect -100 -127549 100 -127511
rect -100 -127583 -84 -127549
rect 84 -127583 100 -127549
rect -100 -127599 100 -127583
rect -100 -127657 100 -127641
rect -100 -127691 -84 -127657
rect 84 -127691 100 -127657
rect -100 -127729 100 -127691
rect -100 -128967 100 -128929
rect -100 -129001 -84 -128967
rect 84 -129001 100 -128967
rect -100 -129017 100 -129001
rect -100 -129075 100 -129059
rect -100 -129109 -84 -129075
rect 84 -129109 100 -129075
rect -100 -129147 100 -129109
rect -100 -130385 100 -130347
rect -100 -130419 -84 -130385
rect 84 -130419 100 -130385
rect -100 -130435 100 -130419
rect -100 -130493 100 -130477
rect -100 -130527 -84 -130493
rect 84 -130527 100 -130493
rect -100 -130565 100 -130527
rect -100 -131803 100 -131765
rect -100 -131837 -84 -131803
rect 84 -131837 100 -131803
rect -100 -131853 100 -131837
rect -100 -131911 100 -131895
rect -100 -131945 -84 -131911
rect 84 -131945 100 -131911
rect -100 -131983 100 -131945
rect -100 -133221 100 -133183
rect -100 -133255 -84 -133221
rect 84 -133255 100 -133221
rect -100 -133271 100 -133255
rect -100 -133329 100 -133313
rect -100 -133363 -84 -133329
rect 84 -133363 100 -133329
rect -100 -133401 100 -133363
rect -100 -134639 100 -134601
rect -100 -134673 -84 -134639
rect 84 -134673 100 -134639
rect -100 -134689 100 -134673
rect -100 -134747 100 -134731
rect -100 -134781 -84 -134747
rect 84 -134781 100 -134747
rect -100 -134819 100 -134781
rect -100 -136057 100 -136019
rect -100 -136091 -84 -136057
rect 84 -136091 100 -136057
rect -100 -136107 100 -136091
rect -100 -136165 100 -136149
rect -100 -136199 -84 -136165
rect 84 -136199 100 -136165
rect -100 -136237 100 -136199
rect -100 -137475 100 -137437
rect -100 -137509 -84 -137475
rect 84 -137509 100 -137475
rect -100 -137525 100 -137509
rect -100 -137583 100 -137567
rect -100 -137617 -84 -137583
rect 84 -137617 100 -137583
rect -100 -137655 100 -137617
rect -100 -138893 100 -138855
rect -100 -138927 -84 -138893
rect 84 -138927 100 -138893
rect -100 -138943 100 -138927
rect -100 -139001 100 -138985
rect -100 -139035 -84 -139001
rect 84 -139035 100 -139001
rect -100 -139073 100 -139035
rect -100 -140311 100 -140273
rect -100 -140345 -84 -140311
rect 84 -140345 100 -140311
rect -100 -140361 100 -140345
rect -100 -140419 100 -140403
rect -100 -140453 -84 -140419
rect 84 -140453 100 -140419
rect -100 -140491 100 -140453
rect -100 -141729 100 -141691
rect -100 -141763 -84 -141729
rect 84 -141763 100 -141729
rect -100 -141779 100 -141763
rect -100 -141837 100 -141821
rect -100 -141871 -84 -141837
rect 84 -141871 100 -141837
rect -100 -141909 100 -141871
rect -100 -143147 100 -143109
rect -100 -143181 -84 -143147
rect 84 -143181 100 -143147
rect -100 -143197 100 -143181
rect -100 -143255 100 -143239
rect -100 -143289 -84 -143255
rect 84 -143289 100 -143255
rect -100 -143327 100 -143289
rect -100 -144565 100 -144527
rect -100 -144599 -84 -144565
rect 84 -144599 100 -144565
rect -100 -144615 100 -144599
rect -100 -144673 100 -144657
rect -100 -144707 -84 -144673
rect 84 -144707 100 -144673
rect -100 -144745 100 -144707
rect -100 -145983 100 -145945
rect -100 -146017 -84 -145983
rect 84 -146017 100 -145983
rect -100 -146033 100 -146017
rect -100 -146091 100 -146075
rect -100 -146125 -84 -146091
rect 84 -146125 100 -146091
rect -100 -146163 100 -146125
rect -100 -147401 100 -147363
rect -100 -147435 -84 -147401
rect 84 -147435 100 -147401
rect -100 -147451 100 -147435
rect -100 -147509 100 -147493
rect -100 -147543 -84 -147509
rect 84 -147543 100 -147509
rect -100 -147581 100 -147543
rect -100 -148819 100 -148781
rect -100 -148853 -84 -148819
rect 84 -148853 100 -148819
rect -100 -148869 100 -148853
rect -100 -148927 100 -148911
rect -100 -148961 -84 -148927
rect 84 -148961 100 -148927
rect -100 -148999 100 -148961
rect -100 -150237 100 -150199
rect -100 -150271 -84 -150237
rect 84 -150271 100 -150237
rect -100 -150287 100 -150271
rect -100 -150345 100 -150329
rect -100 -150379 -84 -150345
rect 84 -150379 100 -150345
rect -100 -150417 100 -150379
rect -100 -151655 100 -151617
rect -100 -151689 -84 -151655
rect 84 -151689 100 -151655
rect -100 -151705 100 -151689
rect -100 -151763 100 -151747
rect -100 -151797 -84 -151763
rect 84 -151797 100 -151763
rect -100 -151835 100 -151797
rect -100 -153073 100 -153035
rect -100 -153107 -84 -153073
rect 84 -153107 100 -153073
rect -100 -153123 100 -153107
rect -100 -153181 100 -153165
rect -100 -153215 -84 -153181
rect 84 -153215 100 -153181
rect -100 -153253 100 -153215
rect -100 -154491 100 -154453
rect -100 -154525 -84 -154491
rect 84 -154525 100 -154491
rect -100 -154541 100 -154525
rect -100 -154599 100 -154583
rect -100 -154633 -84 -154599
rect 84 -154633 100 -154599
rect -100 -154671 100 -154633
rect -100 -155909 100 -155871
rect -100 -155943 -84 -155909
rect 84 -155943 100 -155909
rect -100 -155959 100 -155943
rect -100 -156017 100 -156001
rect -100 -156051 -84 -156017
rect 84 -156051 100 -156017
rect -100 -156089 100 -156051
rect -100 -157327 100 -157289
rect -100 -157361 -84 -157327
rect 84 -157361 100 -157327
rect -100 -157377 100 -157361
rect -100 -157435 100 -157419
rect -100 -157469 -84 -157435
rect 84 -157469 100 -157435
rect -100 -157507 100 -157469
rect -100 -158745 100 -158707
rect -100 -158779 -84 -158745
rect 84 -158779 100 -158745
rect -100 -158795 100 -158779
rect -100 -158853 100 -158837
rect -100 -158887 -84 -158853
rect 84 -158887 100 -158853
rect -100 -158925 100 -158887
rect -100 -160163 100 -160125
rect -100 -160197 -84 -160163
rect 84 -160197 100 -160163
rect -100 -160213 100 -160197
rect -100 -160271 100 -160255
rect -100 -160305 -84 -160271
rect 84 -160305 100 -160271
rect -100 -160343 100 -160305
rect -100 -161581 100 -161543
rect -100 -161615 -84 -161581
rect 84 -161615 100 -161581
rect -100 -161631 100 -161615
rect -100 -161689 100 -161673
rect -100 -161723 -84 -161689
rect 84 -161723 100 -161689
rect -100 -161761 100 -161723
rect -100 -162999 100 -162961
rect -100 -163033 -84 -162999
rect 84 -163033 100 -162999
rect -100 -163049 100 -163033
rect -100 -163107 100 -163091
rect -100 -163141 -84 -163107
rect 84 -163141 100 -163107
rect -100 -163179 100 -163141
rect -100 -164417 100 -164379
rect -100 -164451 -84 -164417
rect 84 -164451 100 -164417
rect -100 -164467 100 -164451
rect -100 -164525 100 -164509
rect -100 -164559 -84 -164525
rect 84 -164559 100 -164525
rect -100 -164597 100 -164559
rect -100 -165835 100 -165797
rect -100 -165869 -84 -165835
rect 84 -165869 100 -165835
rect -100 -165885 100 -165869
rect -100 -165943 100 -165927
rect -100 -165977 -84 -165943
rect 84 -165977 100 -165943
rect -100 -166015 100 -165977
rect -100 -167253 100 -167215
rect -100 -167287 -84 -167253
rect 84 -167287 100 -167253
rect -100 -167303 100 -167287
rect -100 -167361 100 -167345
rect -100 -167395 -84 -167361
rect 84 -167395 100 -167361
rect -100 -167433 100 -167395
rect -100 -168671 100 -168633
rect -100 -168705 -84 -168671
rect 84 -168705 100 -168671
rect -100 -168721 100 -168705
rect -100 -168779 100 -168763
rect -100 -168813 -84 -168779
rect 84 -168813 100 -168779
rect -100 -168851 100 -168813
rect -100 -170089 100 -170051
rect -100 -170123 -84 -170089
rect 84 -170123 100 -170089
rect -100 -170139 100 -170123
rect -100 -170197 100 -170181
rect -100 -170231 -84 -170197
rect 84 -170231 100 -170197
rect -100 -170269 100 -170231
rect -100 -171507 100 -171469
rect -100 -171541 -84 -171507
rect 84 -171541 100 -171507
rect -100 -171557 100 -171541
rect -100 -171615 100 -171599
rect -100 -171649 -84 -171615
rect 84 -171649 100 -171615
rect -100 -171687 100 -171649
rect -100 -172925 100 -172887
rect -100 -172959 -84 -172925
rect 84 -172959 100 -172925
rect -100 -172975 100 -172959
rect -100 -173033 100 -173017
rect -100 -173067 -84 -173033
rect 84 -173067 100 -173033
rect -100 -173105 100 -173067
rect -100 -174343 100 -174305
rect -100 -174377 -84 -174343
rect 84 -174377 100 -174343
rect -100 -174393 100 -174377
rect -100 -174451 100 -174435
rect -100 -174485 -84 -174451
rect 84 -174485 100 -174451
rect -100 -174523 100 -174485
rect -100 -175761 100 -175723
rect -100 -175795 -84 -175761
rect 84 -175795 100 -175761
rect -100 -175811 100 -175795
rect -100 -175869 100 -175853
rect -100 -175903 -84 -175869
rect 84 -175903 100 -175869
rect -100 -175941 100 -175903
rect -100 -177179 100 -177141
rect -100 -177213 -84 -177179
rect 84 -177213 100 -177179
rect -100 -177229 100 -177213
rect -100 -177287 100 -177271
rect -100 -177321 -84 -177287
rect 84 -177321 100 -177287
rect -100 -177359 100 -177321
rect -100 -178597 100 -178559
rect -100 -178631 -84 -178597
rect 84 -178631 100 -178597
rect -100 -178647 100 -178631
rect -100 -178705 100 -178689
rect -100 -178739 -84 -178705
rect 84 -178739 100 -178705
rect -100 -178777 100 -178739
rect -100 -180015 100 -179977
rect -100 -180049 -84 -180015
rect 84 -180049 100 -180015
rect -100 -180065 100 -180049
rect -100 -180123 100 -180107
rect -100 -180157 -84 -180123
rect 84 -180157 100 -180123
rect -100 -180195 100 -180157
rect -100 -181433 100 -181395
rect -100 -181467 -84 -181433
rect 84 -181467 100 -181433
rect -100 -181483 100 -181467
<< polycont >>
rect -84 181433 84 181467
rect -84 180123 84 180157
rect -84 180015 84 180049
rect -84 178705 84 178739
rect -84 178597 84 178631
rect -84 177287 84 177321
rect -84 177179 84 177213
rect -84 175869 84 175903
rect -84 175761 84 175795
rect -84 174451 84 174485
rect -84 174343 84 174377
rect -84 173033 84 173067
rect -84 172925 84 172959
rect -84 171615 84 171649
rect -84 171507 84 171541
rect -84 170197 84 170231
rect -84 170089 84 170123
rect -84 168779 84 168813
rect -84 168671 84 168705
rect -84 167361 84 167395
rect -84 167253 84 167287
rect -84 165943 84 165977
rect -84 165835 84 165869
rect -84 164525 84 164559
rect -84 164417 84 164451
rect -84 163107 84 163141
rect -84 162999 84 163033
rect -84 161689 84 161723
rect -84 161581 84 161615
rect -84 160271 84 160305
rect -84 160163 84 160197
rect -84 158853 84 158887
rect -84 158745 84 158779
rect -84 157435 84 157469
rect -84 157327 84 157361
rect -84 156017 84 156051
rect -84 155909 84 155943
rect -84 154599 84 154633
rect -84 154491 84 154525
rect -84 153181 84 153215
rect -84 153073 84 153107
rect -84 151763 84 151797
rect -84 151655 84 151689
rect -84 150345 84 150379
rect -84 150237 84 150271
rect -84 148927 84 148961
rect -84 148819 84 148853
rect -84 147509 84 147543
rect -84 147401 84 147435
rect -84 146091 84 146125
rect -84 145983 84 146017
rect -84 144673 84 144707
rect -84 144565 84 144599
rect -84 143255 84 143289
rect -84 143147 84 143181
rect -84 141837 84 141871
rect -84 141729 84 141763
rect -84 140419 84 140453
rect -84 140311 84 140345
rect -84 139001 84 139035
rect -84 138893 84 138927
rect -84 137583 84 137617
rect -84 137475 84 137509
rect -84 136165 84 136199
rect -84 136057 84 136091
rect -84 134747 84 134781
rect -84 134639 84 134673
rect -84 133329 84 133363
rect -84 133221 84 133255
rect -84 131911 84 131945
rect -84 131803 84 131837
rect -84 130493 84 130527
rect -84 130385 84 130419
rect -84 129075 84 129109
rect -84 128967 84 129001
rect -84 127657 84 127691
rect -84 127549 84 127583
rect -84 126239 84 126273
rect -84 126131 84 126165
rect -84 124821 84 124855
rect -84 124713 84 124747
rect -84 123403 84 123437
rect -84 123295 84 123329
rect -84 121985 84 122019
rect -84 121877 84 121911
rect -84 120567 84 120601
rect -84 120459 84 120493
rect -84 119149 84 119183
rect -84 119041 84 119075
rect -84 117731 84 117765
rect -84 117623 84 117657
rect -84 116313 84 116347
rect -84 116205 84 116239
rect -84 114895 84 114929
rect -84 114787 84 114821
rect -84 113477 84 113511
rect -84 113369 84 113403
rect -84 112059 84 112093
rect -84 111951 84 111985
rect -84 110641 84 110675
rect -84 110533 84 110567
rect -84 109223 84 109257
rect -84 109115 84 109149
rect -84 107805 84 107839
rect -84 107697 84 107731
rect -84 106387 84 106421
rect -84 106279 84 106313
rect -84 104969 84 105003
rect -84 104861 84 104895
rect -84 103551 84 103585
rect -84 103443 84 103477
rect -84 102133 84 102167
rect -84 102025 84 102059
rect -84 100715 84 100749
rect -84 100607 84 100641
rect -84 99297 84 99331
rect -84 99189 84 99223
rect -84 97879 84 97913
rect -84 97771 84 97805
rect -84 96461 84 96495
rect -84 96353 84 96387
rect -84 95043 84 95077
rect -84 94935 84 94969
rect -84 93625 84 93659
rect -84 93517 84 93551
rect -84 92207 84 92241
rect -84 92099 84 92133
rect -84 90789 84 90823
rect -84 90681 84 90715
rect -84 89371 84 89405
rect -84 89263 84 89297
rect -84 87953 84 87987
rect -84 87845 84 87879
rect -84 86535 84 86569
rect -84 86427 84 86461
rect -84 85117 84 85151
rect -84 85009 84 85043
rect -84 83699 84 83733
rect -84 83591 84 83625
rect -84 82281 84 82315
rect -84 82173 84 82207
rect -84 80863 84 80897
rect -84 80755 84 80789
rect -84 79445 84 79479
rect -84 79337 84 79371
rect -84 78027 84 78061
rect -84 77919 84 77953
rect -84 76609 84 76643
rect -84 76501 84 76535
rect -84 75191 84 75225
rect -84 75083 84 75117
rect -84 73773 84 73807
rect -84 73665 84 73699
rect -84 72355 84 72389
rect -84 72247 84 72281
rect -84 70937 84 70971
rect -84 70829 84 70863
rect -84 69519 84 69553
rect -84 69411 84 69445
rect -84 68101 84 68135
rect -84 67993 84 68027
rect -84 66683 84 66717
rect -84 66575 84 66609
rect -84 65265 84 65299
rect -84 65157 84 65191
rect -84 63847 84 63881
rect -84 63739 84 63773
rect -84 62429 84 62463
rect -84 62321 84 62355
rect -84 61011 84 61045
rect -84 60903 84 60937
rect -84 59593 84 59627
rect -84 59485 84 59519
rect -84 58175 84 58209
rect -84 58067 84 58101
rect -84 56757 84 56791
rect -84 56649 84 56683
rect -84 55339 84 55373
rect -84 55231 84 55265
rect -84 53921 84 53955
rect -84 53813 84 53847
rect -84 52503 84 52537
rect -84 52395 84 52429
rect -84 51085 84 51119
rect -84 50977 84 51011
rect -84 49667 84 49701
rect -84 49559 84 49593
rect -84 48249 84 48283
rect -84 48141 84 48175
rect -84 46831 84 46865
rect -84 46723 84 46757
rect -84 45413 84 45447
rect -84 45305 84 45339
rect -84 43995 84 44029
rect -84 43887 84 43921
rect -84 42577 84 42611
rect -84 42469 84 42503
rect -84 41159 84 41193
rect -84 41051 84 41085
rect -84 39741 84 39775
rect -84 39633 84 39667
rect -84 38323 84 38357
rect -84 38215 84 38249
rect -84 36905 84 36939
rect -84 36797 84 36831
rect -84 35487 84 35521
rect -84 35379 84 35413
rect -84 34069 84 34103
rect -84 33961 84 33995
rect -84 32651 84 32685
rect -84 32543 84 32577
rect -84 31233 84 31267
rect -84 31125 84 31159
rect -84 29815 84 29849
rect -84 29707 84 29741
rect -84 28397 84 28431
rect -84 28289 84 28323
rect -84 26979 84 27013
rect -84 26871 84 26905
rect -84 25561 84 25595
rect -84 25453 84 25487
rect -84 24143 84 24177
rect -84 24035 84 24069
rect -84 22725 84 22759
rect -84 22617 84 22651
rect -84 21307 84 21341
rect -84 21199 84 21233
rect -84 19889 84 19923
rect -84 19781 84 19815
rect -84 18471 84 18505
rect -84 18363 84 18397
rect -84 17053 84 17087
rect -84 16945 84 16979
rect -84 15635 84 15669
rect -84 15527 84 15561
rect -84 14217 84 14251
rect -84 14109 84 14143
rect -84 12799 84 12833
rect -84 12691 84 12725
rect -84 11381 84 11415
rect -84 11273 84 11307
rect -84 9963 84 9997
rect -84 9855 84 9889
rect -84 8545 84 8579
rect -84 8437 84 8471
rect -84 7127 84 7161
rect -84 7019 84 7053
rect -84 5709 84 5743
rect -84 5601 84 5635
rect -84 4291 84 4325
rect -84 4183 84 4217
rect -84 2873 84 2907
rect -84 2765 84 2799
rect -84 1455 84 1489
rect -84 1347 84 1381
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -1381 84 -1347
rect -84 -1489 84 -1455
rect -84 -2799 84 -2765
rect -84 -2907 84 -2873
rect -84 -4217 84 -4183
rect -84 -4325 84 -4291
rect -84 -5635 84 -5601
rect -84 -5743 84 -5709
rect -84 -7053 84 -7019
rect -84 -7161 84 -7127
rect -84 -8471 84 -8437
rect -84 -8579 84 -8545
rect -84 -9889 84 -9855
rect -84 -9997 84 -9963
rect -84 -11307 84 -11273
rect -84 -11415 84 -11381
rect -84 -12725 84 -12691
rect -84 -12833 84 -12799
rect -84 -14143 84 -14109
rect -84 -14251 84 -14217
rect -84 -15561 84 -15527
rect -84 -15669 84 -15635
rect -84 -16979 84 -16945
rect -84 -17087 84 -17053
rect -84 -18397 84 -18363
rect -84 -18505 84 -18471
rect -84 -19815 84 -19781
rect -84 -19923 84 -19889
rect -84 -21233 84 -21199
rect -84 -21341 84 -21307
rect -84 -22651 84 -22617
rect -84 -22759 84 -22725
rect -84 -24069 84 -24035
rect -84 -24177 84 -24143
rect -84 -25487 84 -25453
rect -84 -25595 84 -25561
rect -84 -26905 84 -26871
rect -84 -27013 84 -26979
rect -84 -28323 84 -28289
rect -84 -28431 84 -28397
rect -84 -29741 84 -29707
rect -84 -29849 84 -29815
rect -84 -31159 84 -31125
rect -84 -31267 84 -31233
rect -84 -32577 84 -32543
rect -84 -32685 84 -32651
rect -84 -33995 84 -33961
rect -84 -34103 84 -34069
rect -84 -35413 84 -35379
rect -84 -35521 84 -35487
rect -84 -36831 84 -36797
rect -84 -36939 84 -36905
rect -84 -38249 84 -38215
rect -84 -38357 84 -38323
rect -84 -39667 84 -39633
rect -84 -39775 84 -39741
rect -84 -41085 84 -41051
rect -84 -41193 84 -41159
rect -84 -42503 84 -42469
rect -84 -42611 84 -42577
rect -84 -43921 84 -43887
rect -84 -44029 84 -43995
rect -84 -45339 84 -45305
rect -84 -45447 84 -45413
rect -84 -46757 84 -46723
rect -84 -46865 84 -46831
rect -84 -48175 84 -48141
rect -84 -48283 84 -48249
rect -84 -49593 84 -49559
rect -84 -49701 84 -49667
rect -84 -51011 84 -50977
rect -84 -51119 84 -51085
rect -84 -52429 84 -52395
rect -84 -52537 84 -52503
rect -84 -53847 84 -53813
rect -84 -53955 84 -53921
rect -84 -55265 84 -55231
rect -84 -55373 84 -55339
rect -84 -56683 84 -56649
rect -84 -56791 84 -56757
rect -84 -58101 84 -58067
rect -84 -58209 84 -58175
rect -84 -59519 84 -59485
rect -84 -59627 84 -59593
rect -84 -60937 84 -60903
rect -84 -61045 84 -61011
rect -84 -62355 84 -62321
rect -84 -62463 84 -62429
rect -84 -63773 84 -63739
rect -84 -63881 84 -63847
rect -84 -65191 84 -65157
rect -84 -65299 84 -65265
rect -84 -66609 84 -66575
rect -84 -66717 84 -66683
rect -84 -68027 84 -67993
rect -84 -68135 84 -68101
rect -84 -69445 84 -69411
rect -84 -69553 84 -69519
rect -84 -70863 84 -70829
rect -84 -70971 84 -70937
rect -84 -72281 84 -72247
rect -84 -72389 84 -72355
rect -84 -73699 84 -73665
rect -84 -73807 84 -73773
rect -84 -75117 84 -75083
rect -84 -75225 84 -75191
rect -84 -76535 84 -76501
rect -84 -76643 84 -76609
rect -84 -77953 84 -77919
rect -84 -78061 84 -78027
rect -84 -79371 84 -79337
rect -84 -79479 84 -79445
rect -84 -80789 84 -80755
rect -84 -80897 84 -80863
rect -84 -82207 84 -82173
rect -84 -82315 84 -82281
rect -84 -83625 84 -83591
rect -84 -83733 84 -83699
rect -84 -85043 84 -85009
rect -84 -85151 84 -85117
rect -84 -86461 84 -86427
rect -84 -86569 84 -86535
rect -84 -87879 84 -87845
rect -84 -87987 84 -87953
rect -84 -89297 84 -89263
rect -84 -89405 84 -89371
rect -84 -90715 84 -90681
rect -84 -90823 84 -90789
rect -84 -92133 84 -92099
rect -84 -92241 84 -92207
rect -84 -93551 84 -93517
rect -84 -93659 84 -93625
rect -84 -94969 84 -94935
rect -84 -95077 84 -95043
rect -84 -96387 84 -96353
rect -84 -96495 84 -96461
rect -84 -97805 84 -97771
rect -84 -97913 84 -97879
rect -84 -99223 84 -99189
rect -84 -99331 84 -99297
rect -84 -100641 84 -100607
rect -84 -100749 84 -100715
rect -84 -102059 84 -102025
rect -84 -102167 84 -102133
rect -84 -103477 84 -103443
rect -84 -103585 84 -103551
rect -84 -104895 84 -104861
rect -84 -105003 84 -104969
rect -84 -106313 84 -106279
rect -84 -106421 84 -106387
rect -84 -107731 84 -107697
rect -84 -107839 84 -107805
rect -84 -109149 84 -109115
rect -84 -109257 84 -109223
rect -84 -110567 84 -110533
rect -84 -110675 84 -110641
rect -84 -111985 84 -111951
rect -84 -112093 84 -112059
rect -84 -113403 84 -113369
rect -84 -113511 84 -113477
rect -84 -114821 84 -114787
rect -84 -114929 84 -114895
rect -84 -116239 84 -116205
rect -84 -116347 84 -116313
rect -84 -117657 84 -117623
rect -84 -117765 84 -117731
rect -84 -119075 84 -119041
rect -84 -119183 84 -119149
rect -84 -120493 84 -120459
rect -84 -120601 84 -120567
rect -84 -121911 84 -121877
rect -84 -122019 84 -121985
rect -84 -123329 84 -123295
rect -84 -123437 84 -123403
rect -84 -124747 84 -124713
rect -84 -124855 84 -124821
rect -84 -126165 84 -126131
rect -84 -126273 84 -126239
rect -84 -127583 84 -127549
rect -84 -127691 84 -127657
rect -84 -129001 84 -128967
rect -84 -129109 84 -129075
rect -84 -130419 84 -130385
rect -84 -130527 84 -130493
rect -84 -131837 84 -131803
rect -84 -131945 84 -131911
rect -84 -133255 84 -133221
rect -84 -133363 84 -133329
rect -84 -134673 84 -134639
rect -84 -134781 84 -134747
rect -84 -136091 84 -136057
rect -84 -136199 84 -136165
rect -84 -137509 84 -137475
rect -84 -137617 84 -137583
rect -84 -138927 84 -138893
rect -84 -139035 84 -139001
rect -84 -140345 84 -140311
rect -84 -140453 84 -140419
rect -84 -141763 84 -141729
rect -84 -141871 84 -141837
rect -84 -143181 84 -143147
rect -84 -143289 84 -143255
rect -84 -144599 84 -144565
rect -84 -144707 84 -144673
rect -84 -146017 84 -145983
rect -84 -146125 84 -146091
rect -84 -147435 84 -147401
rect -84 -147543 84 -147509
rect -84 -148853 84 -148819
rect -84 -148961 84 -148927
rect -84 -150271 84 -150237
rect -84 -150379 84 -150345
rect -84 -151689 84 -151655
rect -84 -151797 84 -151763
rect -84 -153107 84 -153073
rect -84 -153215 84 -153181
rect -84 -154525 84 -154491
rect -84 -154633 84 -154599
rect -84 -155943 84 -155909
rect -84 -156051 84 -156017
rect -84 -157361 84 -157327
rect -84 -157469 84 -157435
rect -84 -158779 84 -158745
rect -84 -158887 84 -158853
rect -84 -160197 84 -160163
rect -84 -160305 84 -160271
rect -84 -161615 84 -161581
rect -84 -161723 84 -161689
rect -84 -163033 84 -162999
rect -84 -163141 84 -163107
rect -84 -164451 84 -164417
rect -84 -164559 84 -164525
rect -84 -165869 84 -165835
rect -84 -165977 84 -165943
rect -84 -167287 84 -167253
rect -84 -167395 84 -167361
rect -84 -168705 84 -168671
rect -84 -168813 84 -168779
rect -84 -170123 84 -170089
rect -84 -170231 84 -170197
rect -84 -171541 84 -171507
rect -84 -171649 84 -171615
rect -84 -172959 84 -172925
rect -84 -173067 84 -173033
rect -84 -174377 84 -174343
rect -84 -174485 84 -174451
rect -84 -175795 84 -175761
rect -84 -175903 84 -175869
rect -84 -177213 84 -177179
rect -84 -177321 84 -177287
rect -84 -178631 84 -178597
rect -84 -178739 84 -178705
rect -84 -180049 84 -180015
rect -84 -180157 84 -180123
rect -84 -181467 84 -181433
<< locali >>
rect -280 181571 -184 181605
rect 184 181571 280 181605
rect -280 181509 -246 181571
rect 246 181509 280 181571
rect -100 181433 -84 181467
rect 84 181433 100 181467
rect -146 181383 -112 181399
rect -146 180191 -112 180207
rect 112 181383 146 181399
rect 112 180191 146 180207
rect -100 180123 -84 180157
rect 84 180123 100 180157
rect -100 180015 -84 180049
rect 84 180015 100 180049
rect -146 179965 -112 179981
rect -146 178773 -112 178789
rect 112 179965 146 179981
rect 112 178773 146 178789
rect -100 178705 -84 178739
rect 84 178705 100 178739
rect -100 178597 -84 178631
rect 84 178597 100 178631
rect -146 178547 -112 178563
rect -146 177355 -112 177371
rect 112 178547 146 178563
rect 112 177355 146 177371
rect -100 177287 -84 177321
rect 84 177287 100 177321
rect -100 177179 -84 177213
rect 84 177179 100 177213
rect -146 177129 -112 177145
rect -146 175937 -112 175953
rect 112 177129 146 177145
rect 112 175937 146 175953
rect -100 175869 -84 175903
rect 84 175869 100 175903
rect -100 175761 -84 175795
rect 84 175761 100 175795
rect -146 175711 -112 175727
rect -146 174519 -112 174535
rect 112 175711 146 175727
rect 112 174519 146 174535
rect -100 174451 -84 174485
rect 84 174451 100 174485
rect -100 174343 -84 174377
rect 84 174343 100 174377
rect -146 174293 -112 174309
rect -146 173101 -112 173117
rect 112 174293 146 174309
rect 112 173101 146 173117
rect -100 173033 -84 173067
rect 84 173033 100 173067
rect -100 172925 -84 172959
rect 84 172925 100 172959
rect -146 172875 -112 172891
rect -146 171683 -112 171699
rect 112 172875 146 172891
rect 112 171683 146 171699
rect -100 171615 -84 171649
rect 84 171615 100 171649
rect -100 171507 -84 171541
rect 84 171507 100 171541
rect -146 171457 -112 171473
rect -146 170265 -112 170281
rect 112 171457 146 171473
rect 112 170265 146 170281
rect -100 170197 -84 170231
rect 84 170197 100 170231
rect -100 170089 -84 170123
rect 84 170089 100 170123
rect -146 170039 -112 170055
rect -146 168847 -112 168863
rect 112 170039 146 170055
rect 112 168847 146 168863
rect -100 168779 -84 168813
rect 84 168779 100 168813
rect -100 168671 -84 168705
rect 84 168671 100 168705
rect -146 168621 -112 168637
rect -146 167429 -112 167445
rect 112 168621 146 168637
rect 112 167429 146 167445
rect -100 167361 -84 167395
rect 84 167361 100 167395
rect -100 167253 -84 167287
rect 84 167253 100 167287
rect -146 167203 -112 167219
rect -146 166011 -112 166027
rect 112 167203 146 167219
rect 112 166011 146 166027
rect -100 165943 -84 165977
rect 84 165943 100 165977
rect -100 165835 -84 165869
rect 84 165835 100 165869
rect -146 165785 -112 165801
rect -146 164593 -112 164609
rect 112 165785 146 165801
rect 112 164593 146 164609
rect -100 164525 -84 164559
rect 84 164525 100 164559
rect -100 164417 -84 164451
rect 84 164417 100 164451
rect -146 164367 -112 164383
rect -146 163175 -112 163191
rect 112 164367 146 164383
rect 112 163175 146 163191
rect -100 163107 -84 163141
rect 84 163107 100 163141
rect -100 162999 -84 163033
rect 84 162999 100 163033
rect -146 162949 -112 162965
rect -146 161757 -112 161773
rect 112 162949 146 162965
rect 112 161757 146 161773
rect -100 161689 -84 161723
rect 84 161689 100 161723
rect -100 161581 -84 161615
rect 84 161581 100 161615
rect -146 161531 -112 161547
rect -146 160339 -112 160355
rect 112 161531 146 161547
rect 112 160339 146 160355
rect -100 160271 -84 160305
rect 84 160271 100 160305
rect -100 160163 -84 160197
rect 84 160163 100 160197
rect -146 160113 -112 160129
rect -146 158921 -112 158937
rect 112 160113 146 160129
rect 112 158921 146 158937
rect -100 158853 -84 158887
rect 84 158853 100 158887
rect -100 158745 -84 158779
rect 84 158745 100 158779
rect -146 158695 -112 158711
rect -146 157503 -112 157519
rect 112 158695 146 158711
rect 112 157503 146 157519
rect -100 157435 -84 157469
rect 84 157435 100 157469
rect -100 157327 -84 157361
rect 84 157327 100 157361
rect -146 157277 -112 157293
rect -146 156085 -112 156101
rect 112 157277 146 157293
rect 112 156085 146 156101
rect -100 156017 -84 156051
rect 84 156017 100 156051
rect -100 155909 -84 155943
rect 84 155909 100 155943
rect -146 155859 -112 155875
rect -146 154667 -112 154683
rect 112 155859 146 155875
rect 112 154667 146 154683
rect -100 154599 -84 154633
rect 84 154599 100 154633
rect -100 154491 -84 154525
rect 84 154491 100 154525
rect -146 154441 -112 154457
rect -146 153249 -112 153265
rect 112 154441 146 154457
rect 112 153249 146 153265
rect -100 153181 -84 153215
rect 84 153181 100 153215
rect -100 153073 -84 153107
rect 84 153073 100 153107
rect -146 153023 -112 153039
rect -146 151831 -112 151847
rect 112 153023 146 153039
rect 112 151831 146 151847
rect -100 151763 -84 151797
rect 84 151763 100 151797
rect -100 151655 -84 151689
rect 84 151655 100 151689
rect -146 151605 -112 151621
rect -146 150413 -112 150429
rect 112 151605 146 151621
rect 112 150413 146 150429
rect -100 150345 -84 150379
rect 84 150345 100 150379
rect -100 150237 -84 150271
rect 84 150237 100 150271
rect -146 150187 -112 150203
rect -146 148995 -112 149011
rect 112 150187 146 150203
rect 112 148995 146 149011
rect -100 148927 -84 148961
rect 84 148927 100 148961
rect -100 148819 -84 148853
rect 84 148819 100 148853
rect -146 148769 -112 148785
rect -146 147577 -112 147593
rect 112 148769 146 148785
rect 112 147577 146 147593
rect -100 147509 -84 147543
rect 84 147509 100 147543
rect -100 147401 -84 147435
rect 84 147401 100 147435
rect -146 147351 -112 147367
rect -146 146159 -112 146175
rect 112 147351 146 147367
rect 112 146159 146 146175
rect -100 146091 -84 146125
rect 84 146091 100 146125
rect -100 145983 -84 146017
rect 84 145983 100 146017
rect -146 145933 -112 145949
rect -146 144741 -112 144757
rect 112 145933 146 145949
rect 112 144741 146 144757
rect -100 144673 -84 144707
rect 84 144673 100 144707
rect -100 144565 -84 144599
rect 84 144565 100 144599
rect -146 144515 -112 144531
rect -146 143323 -112 143339
rect 112 144515 146 144531
rect 112 143323 146 143339
rect -100 143255 -84 143289
rect 84 143255 100 143289
rect -100 143147 -84 143181
rect 84 143147 100 143181
rect -146 143097 -112 143113
rect -146 141905 -112 141921
rect 112 143097 146 143113
rect 112 141905 146 141921
rect -100 141837 -84 141871
rect 84 141837 100 141871
rect -100 141729 -84 141763
rect 84 141729 100 141763
rect -146 141679 -112 141695
rect -146 140487 -112 140503
rect 112 141679 146 141695
rect 112 140487 146 140503
rect -100 140419 -84 140453
rect 84 140419 100 140453
rect -100 140311 -84 140345
rect 84 140311 100 140345
rect -146 140261 -112 140277
rect -146 139069 -112 139085
rect 112 140261 146 140277
rect 112 139069 146 139085
rect -100 139001 -84 139035
rect 84 139001 100 139035
rect -100 138893 -84 138927
rect 84 138893 100 138927
rect -146 138843 -112 138859
rect -146 137651 -112 137667
rect 112 138843 146 138859
rect 112 137651 146 137667
rect -100 137583 -84 137617
rect 84 137583 100 137617
rect -100 137475 -84 137509
rect 84 137475 100 137509
rect -146 137425 -112 137441
rect -146 136233 -112 136249
rect 112 137425 146 137441
rect 112 136233 146 136249
rect -100 136165 -84 136199
rect 84 136165 100 136199
rect -100 136057 -84 136091
rect 84 136057 100 136091
rect -146 136007 -112 136023
rect -146 134815 -112 134831
rect 112 136007 146 136023
rect 112 134815 146 134831
rect -100 134747 -84 134781
rect 84 134747 100 134781
rect -100 134639 -84 134673
rect 84 134639 100 134673
rect -146 134589 -112 134605
rect -146 133397 -112 133413
rect 112 134589 146 134605
rect 112 133397 146 133413
rect -100 133329 -84 133363
rect 84 133329 100 133363
rect -100 133221 -84 133255
rect 84 133221 100 133255
rect -146 133171 -112 133187
rect -146 131979 -112 131995
rect 112 133171 146 133187
rect 112 131979 146 131995
rect -100 131911 -84 131945
rect 84 131911 100 131945
rect -100 131803 -84 131837
rect 84 131803 100 131837
rect -146 131753 -112 131769
rect -146 130561 -112 130577
rect 112 131753 146 131769
rect 112 130561 146 130577
rect -100 130493 -84 130527
rect 84 130493 100 130527
rect -100 130385 -84 130419
rect 84 130385 100 130419
rect -146 130335 -112 130351
rect -146 129143 -112 129159
rect 112 130335 146 130351
rect 112 129143 146 129159
rect -100 129075 -84 129109
rect 84 129075 100 129109
rect -100 128967 -84 129001
rect 84 128967 100 129001
rect -146 128917 -112 128933
rect -146 127725 -112 127741
rect 112 128917 146 128933
rect 112 127725 146 127741
rect -100 127657 -84 127691
rect 84 127657 100 127691
rect -100 127549 -84 127583
rect 84 127549 100 127583
rect -146 127499 -112 127515
rect -146 126307 -112 126323
rect 112 127499 146 127515
rect 112 126307 146 126323
rect -100 126239 -84 126273
rect 84 126239 100 126273
rect -100 126131 -84 126165
rect 84 126131 100 126165
rect -146 126081 -112 126097
rect -146 124889 -112 124905
rect 112 126081 146 126097
rect 112 124889 146 124905
rect -100 124821 -84 124855
rect 84 124821 100 124855
rect -100 124713 -84 124747
rect 84 124713 100 124747
rect -146 124663 -112 124679
rect -146 123471 -112 123487
rect 112 124663 146 124679
rect 112 123471 146 123487
rect -100 123403 -84 123437
rect 84 123403 100 123437
rect -100 123295 -84 123329
rect 84 123295 100 123329
rect -146 123245 -112 123261
rect -146 122053 -112 122069
rect 112 123245 146 123261
rect 112 122053 146 122069
rect -100 121985 -84 122019
rect 84 121985 100 122019
rect -100 121877 -84 121911
rect 84 121877 100 121911
rect -146 121827 -112 121843
rect -146 120635 -112 120651
rect 112 121827 146 121843
rect 112 120635 146 120651
rect -100 120567 -84 120601
rect 84 120567 100 120601
rect -100 120459 -84 120493
rect 84 120459 100 120493
rect -146 120409 -112 120425
rect -146 119217 -112 119233
rect 112 120409 146 120425
rect 112 119217 146 119233
rect -100 119149 -84 119183
rect 84 119149 100 119183
rect -100 119041 -84 119075
rect 84 119041 100 119075
rect -146 118991 -112 119007
rect -146 117799 -112 117815
rect 112 118991 146 119007
rect 112 117799 146 117815
rect -100 117731 -84 117765
rect 84 117731 100 117765
rect -100 117623 -84 117657
rect 84 117623 100 117657
rect -146 117573 -112 117589
rect -146 116381 -112 116397
rect 112 117573 146 117589
rect 112 116381 146 116397
rect -100 116313 -84 116347
rect 84 116313 100 116347
rect -100 116205 -84 116239
rect 84 116205 100 116239
rect -146 116155 -112 116171
rect -146 114963 -112 114979
rect 112 116155 146 116171
rect 112 114963 146 114979
rect -100 114895 -84 114929
rect 84 114895 100 114929
rect -100 114787 -84 114821
rect 84 114787 100 114821
rect -146 114737 -112 114753
rect -146 113545 -112 113561
rect 112 114737 146 114753
rect 112 113545 146 113561
rect -100 113477 -84 113511
rect 84 113477 100 113511
rect -100 113369 -84 113403
rect 84 113369 100 113403
rect -146 113319 -112 113335
rect -146 112127 -112 112143
rect 112 113319 146 113335
rect 112 112127 146 112143
rect -100 112059 -84 112093
rect 84 112059 100 112093
rect -100 111951 -84 111985
rect 84 111951 100 111985
rect -146 111901 -112 111917
rect -146 110709 -112 110725
rect 112 111901 146 111917
rect 112 110709 146 110725
rect -100 110641 -84 110675
rect 84 110641 100 110675
rect -100 110533 -84 110567
rect 84 110533 100 110567
rect -146 110483 -112 110499
rect -146 109291 -112 109307
rect 112 110483 146 110499
rect 112 109291 146 109307
rect -100 109223 -84 109257
rect 84 109223 100 109257
rect -100 109115 -84 109149
rect 84 109115 100 109149
rect -146 109065 -112 109081
rect -146 107873 -112 107889
rect 112 109065 146 109081
rect 112 107873 146 107889
rect -100 107805 -84 107839
rect 84 107805 100 107839
rect -100 107697 -84 107731
rect 84 107697 100 107731
rect -146 107647 -112 107663
rect -146 106455 -112 106471
rect 112 107647 146 107663
rect 112 106455 146 106471
rect -100 106387 -84 106421
rect 84 106387 100 106421
rect -100 106279 -84 106313
rect 84 106279 100 106313
rect -146 106229 -112 106245
rect -146 105037 -112 105053
rect 112 106229 146 106245
rect 112 105037 146 105053
rect -100 104969 -84 105003
rect 84 104969 100 105003
rect -100 104861 -84 104895
rect 84 104861 100 104895
rect -146 104811 -112 104827
rect -146 103619 -112 103635
rect 112 104811 146 104827
rect 112 103619 146 103635
rect -100 103551 -84 103585
rect 84 103551 100 103585
rect -100 103443 -84 103477
rect 84 103443 100 103477
rect -146 103393 -112 103409
rect -146 102201 -112 102217
rect 112 103393 146 103409
rect 112 102201 146 102217
rect -100 102133 -84 102167
rect 84 102133 100 102167
rect -100 102025 -84 102059
rect 84 102025 100 102059
rect -146 101975 -112 101991
rect -146 100783 -112 100799
rect 112 101975 146 101991
rect 112 100783 146 100799
rect -100 100715 -84 100749
rect 84 100715 100 100749
rect -100 100607 -84 100641
rect 84 100607 100 100641
rect -146 100557 -112 100573
rect -146 99365 -112 99381
rect 112 100557 146 100573
rect 112 99365 146 99381
rect -100 99297 -84 99331
rect 84 99297 100 99331
rect -100 99189 -84 99223
rect 84 99189 100 99223
rect -146 99139 -112 99155
rect -146 97947 -112 97963
rect 112 99139 146 99155
rect 112 97947 146 97963
rect -100 97879 -84 97913
rect 84 97879 100 97913
rect -100 97771 -84 97805
rect 84 97771 100 97805
rect -146 97721 -112 97737
rect -146 96529 -112 96545
rect 112 97721 146 97737
rect 112 96529 146 96545
rect -100 96461 -84 96495
rect 84 96461 100 96495
rect -100 96353 -84 96387
rect 84 96353 100 96387
rect -146 96303 -112 96319
rect -146 95111 -112 95127
rect 112 96303 146 96319
rect 112 95111 146 95127
rect -100 95043 -84 95077
rect 84 95043 100 95077
rect -100 94935 -84 94969
rect 84 94935 100 94969
rect -146 94885 -112 94901
rect -146 93693 -112 93709
rect 112 94885 146 94901
rect 112 93693 146 93709
rect -100 93625 -84 93659
rect 84 93625 100 93659
rect -100 93517 -84 93551
rect 84 93517 100 93551
rect -146 93467 -112 93483
rect -146 92275 -112 92291
rect 112 93467 146 93483
rect 112 92275 146 92291
rect -100 92207 -84 92241
rect 84 92207 100 92241
rect -100 92099 -84 92133
rect 84 92099 100 92133
rect -146 92049 -112 92065
rect -146 90857 -112 90873
rect 112 92049 146 92065
rect 112 90857 146 90873
rect -100 90789 -84 90823
rect 84 90789 100 90823
rect -100 90681 -84 90715
rect 84 90681 100 90715
rect -146 90631 -112 90647
rect -146 89439 -112 89455
rect 112 90631 146 90647
rect 112 89439 146 89455
rect -100 89371 -84 89405
rect 84 89371 100 89405
rect -100 89263 -84 89297
rect 84 89263 100 89297
rect -146 89213 -112 89229
rect -146 88021 -112 88037
rect 112 89213 146 89229
rect 112 88021 146 88037
rect -100 87953 -84 87987
rect 84 87953 100 87987
rect -100 87845 -84 87879
rect 84 87845 100 87879
rect -146 87795 -112 87811
rect -146 86603 -112 86619
rect 112 87795 146 87811
rect 112 86603 146 86619
rect -100 86535 -84 86569
rect 84 86535 100 86569
rect -100 86427 -84 86461
rect 84 86427 100 86461
rect -146 86377 -112 86393
rect -146 85185 -112 85201
rect 112 86377 146 86393
rect 112 85185 146 85201
rect -100 85117 -84 85151
rect 84 85117 100 85151
rect -100 85009 -84 85043
rect 84 85009 100 85043
rect -146 84959 -112 84975
rect -146 83767 -112 83783
rect 112 84959 146 84975
rect 112 83767 146 83783
rect -100 83699 -84 83733
rect 84 83699 100 83733
rect -100 83591 -84 83625
rect 84 83591 100 83625
rect -146 83541 -112 83557
rect -146 82349 -112 82365
rect 112 83541 146 83557
rect 112 82349 146 82365
rect -100 82281 -84 82315
rect 84 82281 100 82315
rect -100 82173 -84 82207
rect 84 82173 100 82207
rect -146 82123 -112 82139
rect -146 80931 -112 80947
rect 112 82123 146 82139
rect 112 80931 146 80947
rect -100 80863 -84 80897
rect 84 80863 100 80897
rect -100 80755 -84 80789
rect 84 80755 100 80789
rect -146 80705 -112 80721
rect -146 79513 -112 79529
rect 112 80705 146 80721
rect 112 79513 146 79529
rect -100 79445 -84 79479
rect 84 79445 100 79479
rect -100 79337 -84 79371
rect 84 79337 100 79371
rect -146 79287 -112 79303
rect -146 78095 -112 78111
rect 112 79287 146 79303
rect 112 78095 146 78111
rect -100 78027 -84 78061
rect 84 78027 100 78061
rect -100 77919 -84 77953
rect 84 77919 100 77953
rect -146 77869 -112 77885
rect -146 76677 -112 76693
rect 112 77869 146 77885
rect 112 76677 146 76693
rect -100 76609 -84 76643
rect 84 76609 100 76643
rect -100 76501 -84 76535
rect 84 76501 100 76535
rect -146 76451 -112 76467
rect -146 75259 -112 75275
rect 112 76451 146 76467
rect 112 75259 146 75275
rect -100 75191 -84 75225
rect 84 75191 100 75225
rect -100 75083 -84 75117
rect 84 75083 100 75117
rect -146 75033 -112 75049
rect -146 73841 -112 73857
rect 112 75033 146 75049
rect 112 73841 146 73857
rect -100 73773 -84 73807
rect 84 73773 100 73807
rect -100 73665 -84 73699
rect 84 73665 100 73699
rect -146 73615 -112 73631
rect -146 72423 -112 72439
rect 112 73615 146 73631
rect 112 72423 146 72439
rect -100 72355 -84 72389
rect 84 72355 100 72389
rect -100 72247 -84 72281
rect 84 72247 100 72281
rect -146 72197 -112 72213
rect -146 71005 -112 71021
rect 112 72197 146 72213
rect 112 71005 146 71021
rect -100 70937 -84 70971
rect 84 70937 100 70971
rect -100 70829 -84 70863
rect 84 70829 100 70863
rect -146 70779 -112 70795
rect -146 69587 -112 69603
rect 112 70779 146 70795
rect 112 69587 146 69603
rect -100 69519 -84 69553
rect 84 69519 100 69553
rect -100 69411 -84 69445
rect 84 69411 100 69445
rect -146 69361 -112 69377
rect -146 68169 -112 68185
rect 112 69361 146 69377
rect 112 68169 146 68185
rect -100 68101 -84 68135
rect 84 68101 100 68135
rect -100 67993 -84 68027
rect 84 67993 100 68027
rect -146 67943 -112 67959
rect -146 66751 -112 66767
rect 112 67943 146 67959
rect 112 66751 146 66767
rect -100 66683 -84 66717
rect 84 66683 100 66717
rect -100 66575 -84 66609
rect 84 66575 100 66609
rect -146 66525 -112 66541
rect -146 65333 -112 65349
rect 112 66525 146 66541
rect 112 65333 146 65349
rect -100 65265 -84 65299
rect 84 65265 100 65299
rect -100 65157 -84 65191
rect 84 65157 100 65191
rect -146 65107 -112 65123
rect -146 63915 -112 63931
rect 112 65107 146 65123
rect 112 63915 146 63931
rect -100 63847 -84 63881
rect 84 63847 100 63881
rect -100 63739 -84 63773
rect 84 63739 100 63773
rect -146 63689 -112 63705
rect -146 62497 -112 62513
rect 112 63689 146 63705
rect 112 62497 146 62513
rect -100 62429 -84 62463
rect 84 62429 100 62463
rect -100 62321 -84 62355
rect 84 62321 100 62355
rect -146 62271 -112 62287
rect -146 61079 -112 61095
rect 112 62271 146 62287
rect 112 61079 146 61095
rect -100 61011 -84 61045
rect 84 61011 100 61045
rect -100 60903 -84 60937
rect 84 60903 100 60937
rect -146 60853 -112 60869
rect -146 59661 -112 59677
rect 112 60853 146 60869
rect 112 59661 146 59677
rect -100 59593 -84 59627
rect 84 59593 100 59627
rect -100 59485 -84 59519
rect 84 59485 100 59519
rect -146 59435 -112 59451
rect -146 58243 -112 58259
rect 112 59435 146 59451
rect 112 58243 146 58259
rect -100 58175 -84 58209
rect 84 58175 100 58209
rect -100 58067 -84 58101
rect 84 58067 100 58101
rect -146 58017 -112 58033
rect -146 56825 -112 56841
rect 112 58017 146 58033
rect 112 56825 146 56841
rect -100 56757 -84 56791
rect 84 56757 100 56791
rect -100 56649 -84 56683
rect 84 56649 100 56683
rect -146 56599 -112 56615
rect -146 55407 -112 55423
rect 112 56599 146 56615
rect 112 55407 146 55423
rect -100 55339 -84 55373
rect 84 55339 100 55373
rect -100 55231 -84 55265
rect 84 55231 100 55265
rect -146 55181 -112 55197
rect -146 53989 -112 54005
rect 112 55181 146 55197
rect 112 53989 146 54005
rect -100 53921 -84 53955
rect 84 53921 100 53955
rect -100 53813 -84 53847
rect 84 53813 100 53847
rect -146 53763 -112 53779
rect -146 52571 -112 52587
rect 112 53763 146 53779
rect 112 52571 146 52587
rect -100 52503 -84 52537
rect 84 52503 100 52537
rect -100 52395 -84 52429
rect 84 52395 100 52429
rect -146 52345 -112 52361
rect -146 51153 -112 51169
rect 112 52345 146 52361
rect 112 51153 146 51169
rect -100 51085 -84 51119
rect 84 51085 100 51119
rect -100 50977 -84 51011
rect 84 50977 100 51011
rect -146 50927 -112 50943
rect -146 49735 -112 49751
rect 112 50927 146 50943
rect 112 49735 146 49751
rect -100 49667 -84 49701
rect 84 49667 100 49701
rect -100 49559 -84 49593
rect 84 49559 100 49593
rect -146 49509 -112 49525
rect -146 48317 -112 48333
rect 112 49509 146 49525
rect 112 48317 146 48333
rect -100 48249 -84 48283
rect 84 48249 100 48283
rect -100 48141 -84 48175
rect 84 48141 100 48175
rect -146 48091 -112 48107
rect -146 46899 -112 46915
rect 112 48091 146 48107
rect 112 46899 146 46915
rect -100 46831 -84 46865
rect 84 46831 100 46865
rect -100 46723 -84 46757
rect 84 46723 100 46757
rect -146 46673 -112 46689
rect -146 45481 -112 45497
rect 112 46673 146 46689
rect 112 45481 146 45497
rect -100 45413 -84 45447
rect 84 45413 100 45447
rect -100 45305 -84 45339
rect 84 45305 100 45339
rect -146 45255 -112 45271
rect -146 44063 -112 44079
rect 112 45255 146 45271
rect 112 44063 146 44079
rect -100 43995 -84 44029
rect 84 43995 100 44029
rect -100 43887 -84 43921
rect 84 43887 100 43921
rect -146 43837 -112 43853
rect -146 42645 -112 42661
rect 112 43837 146 43853
rect 112 42645 146 42661
rect -100 42577 -84 42611
rect 84 42577 100 42611
rect -100 42469 -84 42503
rect 84 42469 100 42503
rect -146 42419 -112 42435
rect -146 41227 -112 41243
rect 112 42419 146 42435
rect 112 41227 146 41243
rect -100 41159 -84 41193
rect 84 41159 100 41193
rect -100 41051 -84 41085
rect 84 41051 100 41085
rect -146 41001 -112 41017
rect -146 39809 -112 39825
rect 112 41001 146 41017
rect 112 39809 146 39825
rect -100 39741 -84 39775
rect 84 39741 100 39775
rect -100 39633 -84 39667
rect 84 39633 100 39667
rect -146 39583 -112 39599
rect -146 38391 -112 38407
rect 112 39583 146 39599
rect 112 38391 146 38407
rect -100 38323 -84 38357
rect 84 38323 100 38357
rect -100 38215 -84 38249
rect 84 38215 100 38249
rect -146 38165 -112 38181
rect -146 36973 -112 36989
rect 112 38165 146 38181
rect 112 36973 146 36989
rect -100 36905 -84 36939
rect 84 36905 100 36939
rect -100 36797 -84 36831
rect 84 36797 100 36831
rect -146 36747 -112 36763
rect -146 35555 -112 35571
rect 112 36747 146 36763
rect 112 35555 146 35571
rect -100 35487 -84 35521
rect 84 35487 100 35521
rect -100 35379 -84 35413
rect 84 35379 100 35413
rect -146 35329 -112 35345
rect -146 34137 -112 34153
rect 112 35329 146 35345
rect 112 34137 146 34153
rect -100 34069 -84 34103
rect 84 34069 100 34103
rect -100 33961 -84 33995
rect 84 33961 100 33995
rect -146 33911 -112 33927
rect -146 32719 -112 32735
rect 112 33911 146 33927
rect 112 32719 146 32735
rect -100 32651 -84 32685
rect 84 32651 100 32685
rect -100 32543 -84 32577
rect 84 32543 100 32577
rect -146 32493 -112 32509
rect -146 31301 -112 31317
rect 112 32493 146 32509
rect 112 31301 146 31317
rect -100 31233 -84 31267
rect 84 31233 100 31267
rect -100 31125 -84 31159
rect 84 31125 100 31159
rect -146 31075 -112 31091
rect -146 29883 -112 29899
rect 112 31075 146 31091
rect 112 29883 146 29899
rect -100 29815 -84 29849
rect 84 29815 100 29849
rect -100 29707 -84 29741
rect 84 29707 100 29741
rect -146 29657 -112 29673
rect -146 28465 -112 28481
rect 112 29657 146 29673
rect 112 28465 146 28481
rect -100 28397 -84 28431
rect 84 28397 100 28431
rect -100 28289 -84 28323
rect 84 28289 100 28323
rect -146 28239 -112 28255
rect -146 27047 -112 27063
rect 112 28239 146 28255
rect 112 27047 146 27063
rect -100 26979 -84 27013
rect 84 26979 100 27013
rect -100 26871 -84 26905
rect 84 26871 100 26905
rect -146 26821 -112 26837
rect -146 25629 -112 25645
rect 112 26821 146 26837
rect 112 25629 146 25645
rect -100 25561 -84 25595
rect 84 25561 100 25595
rect -100 25453 -84 25487
rect 84 25453 100 25487
rect -146 25403 -112 25419
rect -146 24211 -112 24227
rect 112 25403 146 25419
rect 112 24211 146 24227
rect -100 24143 -84 24177
rect 84 24143 100 24177
rect -100 24035 -84 24069
rect 84 24035 100 24069
rect -146 23985 -112 24001
rect -146 22793 -112 22809
rect 112 23985 146 24001
rect 112 22793 146 22809
rect -100 22725 -84 22759
rect 84 22725 100 22759
rect -100 22617 -84 22651
rect 84 22617 100 22651
rect -146 22567 -112 22583
rect -146 21375 -112 21391
rect 112 22567 146 22583
rect 112 21375 146 21391
rect -100 21307 -84 21341
rect 84 21307 100 21341
rect -100 21199 -84 21233
rect 84 21199 100 21233
rect -146 21149 -112 21165
rect -146 19957 -112 19973
rect 112 21149 146 21165
rect 112 19957 146 19973
rect -100 19889 -84 19923
rect 84 19889 100 19923
rect -100 19781 -84 19815
rect 84 19781 100 19815
rect -146 19731 -112 19747
rect -146 18539 -112 18555
rect 112 19731 146 19747
rect 112 18539 146 18555
rect -100 18471 -84 18505
rect 84 18471 100 18505
rect -100 18363 -84 18397
rect 84 18363 100 18397
rect -146 18313 -112 18329
rect -146 17121 -112 17137
rect 112 18313 146 18329
rect 112 17121 146 17137
rect -100 17053 -84 17087
rect 84 17053 100 17087
rect -100 16945 -84 16979
rect 84 16945 100 16979
rect -146 16895 -112 16911
rect -146 15703 -112 15719
rect 112 16895 146 16911
rect 112 15703 146 15719
rect -100 15635 -84 15669
rect 84 15635 100 15669
rect -100 15527 -84 15561
rect 84 15527 100 15561
rect -146 15477 -112 15493
rect -146 14285 -112 14301
rect 112 15477 146 15493
rect 112 14285 146 14301
rect -100 14217 -84 14251
rect 84 14217 100 14251
rect -100 14109 -84 14143
rect 84 14109 100 14143
rect -146 14059 -112 14075
rect -146 12867 -112 12883
rect 112 14059 146 14075
rect 112 12867 146 12883
rect -100 12799 -84 12833
rect 84 12799 100 12833
rect -100 12691 -84 12725
rect 84 12691 100 12725
rect -146 12641 -112 12657
rect -146 11449 -112 11465
rect 112 12641 146 12657
rect 112 11449 146 11465
rect -100 11381 -84 11415
rect 84 11381 100 11415
rect -100 11273 -84 11307
rect 84 11273 100 11307
rect -146 11223 -112 11239
rect -146 10031 -112 10047
rect 112 11223 146 11239
rect 112 10031 146 10047
rect -100 9963 -84 9997
rect 84 9963 100 9997
rect -100 9855 -84 9889
rect 84 9855 100 9889
rect -146 9805 -112 9821
rect -146 8613 -112 8629
rect 112 9805 146 9821
rect 112 8613 146 8629
rect -100 8545 -84 8579
rect 84 8545 100 8579
rect -100 8437 -84 8471
rect 84 8437 100 8471
rect -146 8387 -112 8403
rect -146 7195 -112 7211
rect 112 8387 146 8403
rect 112 7195 146 7211
rect -100 7127 -84 7161
rect 84 7127 100 7161
rect -100 7019 -84 7053
rect 84 7019 100 7053
rect -146 6969 -112 6985
rect -146 5777 -112 5793
rect 112 6969 146 6985
rect 112 5777 146 5793
rect -100 5709 -84 5743
rect 84 5709 100 5743
rect -100 5601 -84 5635
rect 84 5601 100 5635
rect -146 5551 -112 5567
rect -146 4359 -112 4375
rect 112 5551 146 5567
rect 112 4359 146 4375
rect -100 4291 -84 4325
rect 84 4291 100 4325
rect -100 4183 -84 4217
rect 84 4183 100 4217
rect -146 4133 -112 4149
rect -146 2941 -112 2957
rect 112 4133 146 4149
rect 112 2941 146 2957
rect -100 2873 -84 2907
rect 84 2873 100 2907
rect -100 2765 -84 2799
rect 84 2765 100 2799
rect -146 2715 -112 2731
rect -146 1523 -112 1539
rect 112 2715 146 2731
rect 112 1523 146 1539
rect -100 1455 -84 1489
rect 84 1455 100 1489
rect -100 1347 -84 1381
rect 84 1347 100 1381
rect -146 1297 -112 1313
rect -146 105 -112 121
rect 112 1297 146 1313
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -1313 -112 -1297
rect 112 -121 146 -105
rect 112 -1313 146 -1297
rect -100 -1381 -84 -1347
rect 84 -1381 100 -1347
rect -100 -1489 -84 -1455
rect 84 -1489 100 -1455
rect -146 -1539 -112 -1523
rect -146 -2731 -112 -2715
rect 112 -1539 146 -1523
rect 112 -2731 146 -2715
rect -100 -2799 -84 -2765
rect 84 -2799 100 -2765
rect -100 -2907 -84 -2873
rect 84 -2907 100 -2873
rect -146 -2957 -112 -2941
rect -146 -4149 -112 -4133
rect 112 -2957 146 -2941
rect 112 -4149 146 -4133
rect -100 -4217 -84 -4183
rect 84 -4217 100 -4183
rect -100 -4325 -84 -4291
rect 84 -4325 100 -4291
rect -146 -4375 -112 -4359
rect -146 -5567 -112 -5551
rect 112 -4375 146 -4359
rect 112 -5567 146 -5551
rect -100 -5635 -84 -5601
rect 84 -5635 100 -5601
rect -100 -5743 -84 -5709
rect 84 -5743 100 -5709
rect -146 -5793 -112 -5777
rect -146 -6985 -112 -6969
rect 112 -5793 146 -5777
rect 112 -6985 146 -6969
rect -100 -7053 -84 -7019
rect 84 -7053 100 -7019
rect -100 -7161 -84 -7127
rect 84 -7161 100 -7127
rect -146 -7211 -112 -7195
rect -146 -8403 -112 -8387
rect 112 -7211 146 -7195
rect 112 -8403 146 -8387
rect -100 -8471 -84 -8437
rect 84 -8471 100 -8437
rect -100 -8579 -84 -8545
rect 84 -8579 100 -8545
rect -146 -8629 -112 -8613
rect -146 -9821 -112 -9805
rect 112 -8629 146 -8613
rect 112 -9821 146 -9805
rect -100 -9889 -84 -9855
rect 84 -9889 100 -9855
rect -100 -9997 -84 -9963
rect 84 -9997 100 -9963
rect -146 -10047 -112 -10031
rect -146 -11239 -112 -11223
rect 112 -10047 146 -10031
rect 112 -11239 146 -11223
rect -100 -11307 -84 -11273
rect 84 -11307 100 -11273
rect -100 -11415 -84 -11381
rect 84 -11415 100 -11381
rect -146 -11465 -112 -11449
rect -146 -12657 -112 -12641
rect 112 -11465 146 -11449
rect 112 -12657 146 -12641
rect -100 -12725 -84 -12691
rect 84 -12725 100 -12691
rect -100 -12833 -84 -12799
rect 84 -12833 100 -12799
rect -146 -12883 -112 -12867
rect -146 -14075 -112 -14059
rect 112 -12883 146 -12867
rect 112 -14075 146 -14059
rect -100 -14143 -84 -14109
rect 84 -14143 100 -14109
rect -100 -14251 -84 -14217
rect 84 -14251 100 -14217
rect -146 -14301 -112 -14285
rect -146 -15493 -112 -15477
rect 112 -14301 146 -14285
rect 112 -15493 146 -15477
rect -100 -15561 -84 -15527
rect 84 -15561 100 -15527
rect -100 -15669 -84 -15635
rect 84 -15669 100 -15635
rect -146 -15719 -112 -15703
rect -146 -16911 -112 -16895
rect 112 -15719 146 -15703
rect 112 -16911 146 -16895
rect -100 -16979 -84 -16945
rect 84 -16979 100 -16945
rect -100 -17087 -84 -17053
rect 84 -17087 100 -17053
rect -146 -17137 -112 -17121
rect -146 -18329 -112 -18313
rect 112 -17137 146 -17121
rect 112 -18329 146 -18313
rect -100 -18397 -84 -18363
rect 84 -18397 100 -18363
rect -100 -18505 -84 -18471
rect 84 -18505 100 -18471
rect -146 -18555 -112 -18539
rect -146 -19747 -112 -19731
rect 112 -18555 146 -18539
rect 112 -19747 146 -19731
rect -100 -19815 -84 -19781
rect 84 -19815 100 -19781
rect -100 -19923 -84 -19889
rect 84 -19923 100 -19889
rect -146 -19973 -112 -19957
rect -146 -21165 -112 -21149
rect 112 -19973 146 -19957
rect 112 -21165 146 -21149
rect -100 -21233 -84 -21199
rect 84 -21233 100 -21199
rect -100 -21341 -84 -21307
rect 84 -21341 100 -21307
rect -146 -21391 -112 -21375
rect -146 -22583 -112 -22567
rect 112 -21391 146 -21375
rect 112 -22583 146 -22567
rect -100 -22651 -84 -22617
rect 84 -22651 100 -22617
rect -100 -22759 -84 -22725
rect 84 -22759 100 -22725
rect -146 -22809 -112 -22793
rect -146 -24001 -112 -23985
rect 112 -22809 146 -22793
rect 112 -24001 146 -23985
rect -100 -24069 -84 -24035
rect 84 -24069 100 -24035
rect -100 -24177 -84 -24143
rect 84 -24177 100 -24143
rect -146 -24227 -112 -24211
rect -146 -25419 -112 -25403
rect 112 -24227 146 -24211
rect 112 -25419 146 -25403
rect -100 -25487 -84 -25453
rect 84 -25487 100 -25453
rect -100 -25595 -84 -25561
rect 84 -25595 100 -25561
rect -146 -25645 -112 -25629
rect -146 -26837 -112 -26821
rect 112 -25645 146 -25629
rect 112 -26837 146 -26821
rect -100 -26905 -84 -26871
rect 84 -26905 100 -26871
rect -100 -27013 -84 -26979
rect 84 -27013 100 -26979
rect -146 -27063 -112 -27047
rect -146 -28255 -112 -28239
rect 112 -27063 146 -27047
rect 112 -28255 146 -28239
rect -100 -28323 -84 -28289
rect 84 -28323 100 -28289
rect -100 -28431 -84 -28397
rect 84 -28431 100 -28397
rect -146 -28481 -112 -28465
rect -146 -29673 -112 -29657
rect 112 -28481 146 -28465
rect 112 -29673 146 -29657
rect -100 -29741 -84 -29707
rect 84 -29741 100 -29707
rect -100 -29849 -84 -29815
rect 84 -29849 100 -29815
rect -146 -29899 -112 -29883
rect -146 -31091 -112 -31075
rect 112 -29899 146 -29883
rect 112 -31091 146 -31075
rect -100 -31159 -84 -31125
rect 84 -31159 100 -31125
rect -100 -31267 -84 -31233
rect 84 -31267 100 -31233
rect -146 -31317 -112 -31301
rect -146 -32509 -112 -32493
rect 112 -31317 146 -31301
rect 112 -32509 146 -32493
rect -100 -32577 -84 -32543
rect 84 -32577 100 -32543
rect -100 -32685 -84 -32651
rect 84 -32685 100 -32651
rect -146 -32735 -112 -32719
rect -146 -33927 -112 -33911
rect 112 -32735 146 -32719
rect 112 -33927 146 -33911
rect -100 -33995 -84 -33961
rect 84 -33995 100 -33961
rect -100 -34103 -84 -34069
rect 84 -34103 100 -34069
rect -146 -34153 -112 -34137
rect -146 -35345 -112 -35329
rect 112 -34153 146 -34137
rect 112 -35345 146 -35329
rect -100 -35413 -84 -35379
rect 84 -35413 100 -35379
rect -100 -35521 -84 -35487
rect 84 -35521 100 -35487
rect -146 -35571 -112 -35555
rect -146 -36763 -112 -36747
rect 112 -35571 146 -35555
rect 112 -36763 146 -36747
rect -100 -36831 -84 -36797
rect 84 -36831 100 -36797
rect -100 -36939 -84 -36905
rect 84 -36939 100 -36905
rect -146 -36989 -112 -36973
rect -146 -38181 -112 -38165
rect 112 -36989 146 -36973
rect 112 -38181 146 -38165
rect -100 -38249 -84 -38215
rect 84 -38249 100 -38215
rect -100 -38357 -84 -38323
rect 84 -38357 100 -38323
rect -146 -38407 -112 -38391
rect -146 -39599 -112 -39583
rect 112 -38407 146 -38391
rect 112 -39599 146 -39583
rect -100 -39667 -84 -39633
rect 84 -39667 100 -39633
rect -100 -39775 -84 -39741
rect 84 -39775 100 -39741
rect -146 -39825 -112 -39809
rect -146 -41017 -112 -41001
rect 112 -39825 146 -39809
rect 112 -41017 146 -41001
rect -100 -41085 -84 -41051
rect 84 -41085 100 -41051
rect -100 -41193 -84 -41159
rect 84 -41193 100 -41159
rect -146 -41243 -112 -41227
rect -146 -42435 -112 -42419
rect 112 -41243 146 -41227
rect 112 -42435 146 -42419
rect -100 -42503 -84 -42469
rect 84 -42503 100 -42469
rect -100 -42611 -84 -42577
rect 84 -42611 100 -42577
rect -146 -42661 -112 -42645
rect -146 -43853 -112 -43837
rect 112 -42661 146 -42645
rect 112 -43853 146 -43837
rect -100 -43921 -84 -43887
rect 84 -43921 100 -43887
rect -100 -44029 -84 -43995
rect 84 -44029 100 -43995
rect -146 -44079 -112 -44063
rect -146 -45271 -112 -45255
rect 112 -44079 146 -44063
rect 112 -45271 146 -45255
rect -100 -45339 -84 -45305
rect 84 -45339 100 -45305
rect -100 -45447 -84 -45413
rect 84 -45447 100 -45413
rect -146 -45497 -112 -45481
rect -146 -46689 -112 -46673
rect 112 -45497 146 -45481
rect 112 -46689 146 -46673
rect -100 -46757 -84 -46723
rect 84 -46757 100 -46723
rect -100 -46865 -84 -46831
rect 84 -46865 100 -46831
rect -146 -46915 -112 -46899
rect -146 -48107 -112 -48091
rect 112 -46915 146 -46899
rect 112 -48107 146 -48091
rect -100 -48175 -84 -48141
rect 84 -48175 100 -48141
rect -100 -48283 -84 -48249
rect 84 -48283 100 -48249
rect -146 -48333 -112 -48317
rect -146 -49525 -112 -49509
rect 112 -48333 146 -48317
rect 112 -49525 146 -49509
rect -100 -49593 -84 -49559
rect 84 -49593 100 -49559
rect -100 -49701 -84 -49667
rect 84 -49701 100 -49667
rect -146 -49751 -112 -49735
rect -146 -50943 -112 -50927
rect 112 -49751 146 -49735
rect 112 -50943 146 -50927
rect -100 -51011 -84 -50977
rect 84 -51011 100 -50977
rect -100 -51119 -84 -51085
rect 84 -51119 100 -51085
rect -146 -51169 -112 -51153
rect -146 -52361 -112 -52345
rect 112 -51169 146 -51153
rect 112 -52361 146 -52345
rect -100 -52429 -84 -52395
rect 84 -52429 100 -52395
rect -100 -52537 -84 -52503
rect 84 -52537 100 -52503
rect -146 -52587 -112 -52571
rect -146 -53779 -112 -53763
rect 112 -52587 146 -52571
rect 112 -53779 146 -53763
rect -100 -53847 -84 -53813
rect 84 -53847 100 -53813
rect -100 -53955 -84 -53921
rect 84 -53955 100 -53921
rect -146 -54005 -112 -53989
rect -146 -55197 -112 -55181
rect 112 -54005 146 -53989
rect 112 -55197 146 -55181
rect -100 -55265 -84 -55231
rect 84 -55265 100 -55231
rect -100 -55373 -84 -55339
rect 84 -55373 100 -55339
rect -146 -55423 -112 -55407
rect -146 -56615 -112 -56599
rect 112 -55423 146 -55407
rect 112 -56615 146 -56599
rect -100 -56683 -84 -56649
rect 84 -56683 100 -56649
rect -100 -56791 -84 -56757
rect 84 -56791 100 -56757
rect -146 -56841 -112 -56825
rect -146 -58033 -112 -58017
rect 112 -56841 146 -56825
rect 112 -58033 146 -58017
rect -100 -58101 -84 -58067
rect 84 -58101 100 -58067
rect -100 -58209 -84 -58175
rect 84 -58209 100 -58175
rect -146 -58259 -112 -58243
rect -146 -59451 -112 -59435
rect 112 -58259 146 -58243
rect 112 -59451 146 -59435
rect -100 -59519 -84 -59485
rect 84 -59519 100 -59485
rect -100 -59627 -84 -59593
rect 84 -59627 100 -59593
rect -146 -59677 -112 -59661
rect -146 -60869 -112 -60853
rect 112 -59677 146 -59661
rect 112 -60869 146 -60853
rect -100 -60937 -84 -60903
rect 84 -60937 100 -60903
rect -100 -61045 -84 -61011
rect 84 -61045 100 -61011
rect -146 -61095 -112 -61079
rect -146 -62287 -112 -62271
rect 112 -61095 146 -61079
rect 112 -62287 146 -62271
rect -100 -62355 -84 -62321
rect 84 -62355 100 -62321
rect -100 -62463 -84 -62429
rect 84 -62463 100 -62429
rect -146 -62513 -112 -62497
rect -146 -63705 -112 -63689
rect 112 -62513 146 -62497
rect 112 -63705 146 -63689
rect -100 -63773 -84 -63739
rect 84 -63773 100 -63739
rect -100 -63881 -84 -63847
rect 84 -63881 100 -63847
rect -146 -63931 -112 -63915
rect -146 -65123 -112 -65107
rect 112 -63931 146 -63915
rect 112 -65123 146 -65107
rect -100 -65191 -84 -65157
rect 84 -65191 100 -65157
rect -100 -65299 -84 -65265
rect 84 -65299 100 -65265
rect -146 -65349 -112 -65333
rect -146 -66541 -112 -66525
rect 112 -65349 146 -65333
rect 112 -66541 146 -66525
rect -100 -66609 -84 -66575
rect 84 -66609 100 -66575
rect -100 -66717 -84 -66683
rect 84 -66717 100 -66683
rect -146 -66767 -112 -66751
rect -146 -67959 -112 -67943
rect 112 -66767 146 -66751
rect 112 -67959 146 -67943
rect -100 -68027 -84 -67993
rect 84 -68027 100 -67993
rect -100 -68135 -84 -68101
rect 84 -68135 100 -68101
rect -146 -68185 -112 -68169
rect -146 -69377 -112 -69361
rect 112 -68185 146 -68169
rect 112 -69377 146 -69361
rect -100 -69445 -84 -69411
rect 84 -69445 100 -69411
rect -100 -69553 -84 -69519
rect 84 -69553 100 -69519
rect -146 -69603 -112 -69587
rect -146 -70795 -112 -70779
rect 112 -69603 146 -69587
rect 112 -70795 146 -70779
rect -100 -70863 -84 -70829
rect 84 -70863 100 -70829
rect -100 -70971 -84 -70937
rect 84 -70971 100 -70937
rect -146 -71021 -112 -71005
rect -146 -72213 -112 -72197
rect 112 -71021 146 -71005
rect 112 -72213 146 -72197
rect -100 -72281 -84 -72247
rect 84 -72281 100 -72247
rect -100 -72389 -84 -72355
rect 84 -72389 100 -72355
rect -146 -72439 -112 -72423
rect -146 -73631 -112 -73615
rect 112 -72439 146 -72423
rect 112 -73631 146 -73615
rect -100 -73699 -84 -73665
rect 84 -73699 100 -73665
rect -100 -73807 -84 -73773
rect 84 -73807 100 -73773
rect -146 -73857 -112 -73841
rect -146 -75049 -112 -75033
rect 112 -73857 146 -73841
rect 112 -75049 146 -75033
rect -100 -75117 -84 -75083
rect 84 -75117 100 -75083
rect -100 -75225 -84 -75191
rect 84 -75225 100 -75191
rect -146 -75275 -112 -75259
rect -146 -76467 -112 -76451
rect 112 -75275 146 -75259
rect 112 -76467 146 -76451
rect -100 -76535 -84 -76501
rect 84 -76535 100 -76501
rect -100 -76643 -84 -76609
rect 84 -76643 100 -76609
rect -146 -76693 -112 -76677
rect -146 -77885 -112 -77869
rect 112 -76693 146 -76677
rect 112 -77885 146 -77869
rect -100 -77953 -84 -77919
rect 84 -77953 100 -77919
rect -100 -78061 -84 -78027
rect 84 -78061 100 -78027
rect -146 -78111 -112 -78095
rect -146 -79303 -112 -79287
rect 112 -78111 146 -78095
rect 112 -79303 146 -79287
rect -100 -79371 -84 -79337
rect 84 -79371 100 -79337
rect -100 -79479 -84 -79445
rect 84 -79479 100 -79445
rect -146 -79529 -112 -79513
rect -146 -80721 -112 -80705
rect 112 -79529 146 -79513
rect 112 -80721 146 -80705
rect -100 -80789 -84 -80755
rect 84 -80789 100 -80755
rect -100 -80897 -84 -80863
rect 84 -80897 100 -80863
rect -146 -80947 -112 -80931
rect -146 -82139 -112 -82123
rect 112 -80947 146 -80931
rect 112 -82139 146 -82123
rect -100 -82207 -84 -82173
rect 84 -82207 100 -82173
rect -100 -82315 -84 -82281
rect 84 -82315 100 -82281
rect -146 -82365 -112 -82349
rect -146 -83557 -112 -83541
rect 112 -82365 146 -82349
rect 112 -83557 146 -83541
rect -100 -83625 -84 -83591
rect 84 -83625 100 -83591
rect -100 -83733 -84 -83699
rect 84 -83733 100 -83699
rect -146 -83783 -112 -83767
rect -146 -84975 -112 -84959
rect 112 -83783 146 -83767
rect 112 -84975 146 -84959
rect -100 -85043 -84 -85009
rect 84 -85043 100 -85009
rect -100 -85151 -84 -85117
rect 84 -85151 100 -85117
rect -146 -85201 -112 -85185
rect -146 -86393 -112 -86377
rect 112 -85201 146 -85185
rect 112 -86393 146 -86377
rect -100 -86461 -84 -86427
rect 84 -86461 100 -86427
rect -100 -86569 -84 -86535
rect 84 -86569 100 -86535
rect -146 -86619 -112 -86603
rect -146 -87811 -112 -87795
rect 112 -86619 146 -86603
rect 112 -87811 146 -87795
rect -100 -87879 -84 -87845
rect 84 -87879 100 -87845
rect -100 -87987 -84 -87953
rect 84 -87987 100 -87953
rect -146 -88037 -112 -88021
rect -146 -89229 -112 -89213
rect 112 -88037 146 -88021
rect 112 -89229 146 -89213
rect -100 -89297 -84 -89263
rect 84 -89297 100 -89263
rect -100 -89405 -84 -89371
rect 84 -89405 100 -89371
rect -146 -89455 -112 -89439
rect -146 -90647 -112 -90631
rect 112 -89455 146 -89439
rect 112 -90647 146 -90631
rect -100 -90715 -84 -90681
rect 84 -90715 100 -90681
rect -100 -90823 -84 -90789
rect 84 -90823 100 -90789
rect -146 -90873 -112 -90857
rect -146 -92065 -112 -92049
rect 112 -90873 146 -90857
rect 112 -92065 146 -92049
rect -100 -92133 -84 -92099
rect 84 -92133 100 -92099
rect -100 -92241 -84 -92207
rect 84 -92241 100 -92207
rect -146 -92291 -112 -92275
rect -146 -93483 -112 -93467
rect 112 -92291 146 -92275
rect 112 -93483 146 -93467
rect -100 -93551 -84 -93517
rect 84 -93551 100 -93517
rect -100 -93659 -84 -93625
rect 84 -93659 100 -93625
rect -146 -93709 -112 -93693
rect -146 -94901 -112 -94885
rect 112 -93709 146 -93693
rect 112 -94901 146 -94885
rect -100 -94969 -84 -94935
rect 84 -94969 100 -94935
rect -100 -95077 -84 -95043
rect 84 -95077 100 -95043
rect -146 -95127 -112 -95111
rect -146 -96319 -112 -96303
rect 112 -95127 146 -95111
rect 112 -96319 146 -96303
rect -100 -96387 -84 -96353
rect 84 -96387 100 -96353
rect -100 -96495 -84 -96461
rect 84 -96495 100 -96461
rect -146 -96545 -112 -96529
rect -146 -97737 -112 -97721
rect 112 -96545 146 -96529
rect 112 -97737 146 -97721
rect -100 -97805 -84 -97771
rect 84 -97805 100 -97771
rect -100 -97913 -84 -97879
rect 84 -97913 100 -97879
rect -146 -97963 -112 -97947
rect -146 -99155 -112 -99139
rect 112 -97963 146 -97947
rect 112 -99155 146 -99139
rect -100 -99223 -84 -99189
rect 84 -99223 100 -99189
rect -100 -99331 -84 -99297
rect 84 -99331 100 -99297
rect -146 -99381 -112 -99365
rect -146 -100573 -112 -100557
rect 112 -99381 146 -99365
rect 112 -100573 146 -100557
rect -100 -100641 -84 -100607
rect 84 -100641 100 -100607
rect -100 -100749 -84 -100715
rect 84 -100749 100 -100715
rect -146 -100799 -112 -100783
rect -146 -101991 -112 -101975
rect 112 -100799 146 -100783
rect 112 -101991 146 -101975
rect -100 -102059 -84 -102025
rect 84 -102059 100 -102025
rect -100 -102167 -84 -102133
rect 84 -102167 100 -102133
rect -146 -102217 -112 -102201
rect -146 -103409 -112 -103393
rect 112 -102217 146 -102201
rect 112 -103409 146 -103393
rect -100 -103477 -84 -103443
rect 84 -103477 100 -103443
rect -100 -103585 -84 -103551
rect 84 -103585 100 -103551
rect -146 -103635 -112 -103619
rect -146 -104827 -112 -104811
rect 112 -103635 146 -103619
rect 112 -104827 146 -104811
rect -100 -104895 -84 -104861
rect 84 -104895 100 -104861
rect -100 -105003 -84 -104969
rect 84 -105003 100 -104969
rect -146 -105053 -112 -105037
rect -146 -106245 -112 -106229
rect 112 -105053 146 -105037
rect 112 -106245 146 -106229
rect -100 -106313 -84 -106279
rect 84 -106313 100 -106279
rect -100 -106421 -84 -106387
rect 84 -106421 100 -106387
rect -146 -106471 -112 -106455
rect -146 -107663 -112 -107647
rect 112 -106471 146 -106455
rect 112 -107663 146 -107647
rect -100 -107731 -84 -107697
rect 84 -107731 100 -107697
rect -100 -107839 -84 -107805
rect 84 -107839 100 -107805
rect -146 -107889 -112 -107873
rect -146 -109081 -112 -109065
rect 112 -107889 146 -107873
rect 112 -109081 146 -109065
rect -100 -109149 -84 -109115
rect 84 -109149 100 -109115
rect -100 -109257 -84 -109223
rect 84 -109257 100 -109223
rect -146 -109307 -112 -109291
rect -146 -110499 -112 -110483
rect 112 -109307 146 -109291
rect 112 -110499 146 -110483
rect -100 -110567 -84 -110533
rect 84 -110567 100 -110533
rect -100 -110675 -84 -110641
rect 84 -110675 100 -110641
rect -146 -110725 -112 -110709
rect -146 -111917 -112 -111901
rect 112 -110725 146 -110709
rect 112 -111917 146 -111901
rect -100 -111985 -84 -111951
rect 84 -111985 100 -111951
rect -100 -112093 -84 -112059
rect 84 -112093 100 -112059
rect -146 -112143 -112 -112127
rect -146 -113335 -112 -113319
rect 112 -112143 146 -112127
rect 112 -113335 146 -113319
rect -100 -113403 -84 -113369
rect 84 -113403 100 -113369
rect -100 -113511 -84 -113477
rect 84 -113511 100 -113477
rect -146 -113561 -112 -113545
rect -146 -114753 -112 -114737
rect 112 -113561 146 -113545
rect 112 -114753 146 -114737
rect -100 -114821 -84 -114787
rect 84 -114821 100 -114787
rect -100 -114929 -84 -114895
rect 84 -114929 100 -114895
rect -146 -114979 -112 -114963
rect -146 -116171 -112 -116155
rect 112 -114979 146 -114963
rect 112 -116171 146 -116155
rect -100 -116239 -84 -116205
rect 84 -116239 100 -116205
rect -100 -116347 -84 -116313
rect 84 -116347 100 -116313
rect -146 -116397 -112 -116381
rect -146 -117589 -112 -117573
rect 112 -116397 146 -116381
rect 112 -117589 146 -117573
rect -100 -117657 -84 -117623
rect 84 -117657 100 -117623
rect -100 -117765 -84 -117731
rect 84 -117765 100 -117731
rect -146 -117815 -112 -117799
rect -146 -119007 -112 -118991
rect 112 -117815 146 -117799
rect 112 -119007 146 -118991
rect -100 -119075 -84 -119041
rect 84 -119075 100 -119041
rect -100 -119183 -84 -119149
rect 84 -119183 100 -119149
rect -146 -119233 -112 -119217
rect -146 -120425 -112 -120409
rect 112 -119233 146 -119217
rect 112 -120425 146 -120409
rect -100 -120493 -84 -120459
rect 84 -120493 100 -120459
rect -100 -120601 -84 -120567
rect 84 -120601 100 -120567
rect -146 -120651 -112 -120635
rect -146 -121843 -112 -121827
rect 112 -120651 146 -120635
rect 112 -121843 146 -121827
rect -100 -121911 -84 -121877
rect 84 -121911 100 -121877
rect -100 -122019 -84 -121985
rect 84 -122019 100 -121985
rect -146 -122069 -112 -122053
rect -146 -123261 -112 -123245
rect 112 -122069 146 -122053
rect 112 -123261 146 -123245
rect -100 -123329 -84 -123295
rect 84 -123329 100 -123295
rect -100 -123437 -84 -123403
rect 84 -123437 100 -123403
rect -146 -123487 -112 -123471
rect -146 -124679 -112 -124663
rect 112 -123487 146 -123471
rect 112 -124679 146 -124663
rect -100 -124747 -84 -124713
rect 84 -124747 100 -124713
rect -100 -124855 -84 -124821
rect 84 -124855 100 -124821
rect -146 -124905 -112 -124889
rect -146 -126097 -112 -126081
rect 112 -124905 146 -124889
rect 112 -126097 146 -126081
rect -100 -126165 -84 -126131
rect 84 -126165 100 -126131
rect -100 -126273 -84 -126239
rect 84 -126273 100 -126239
rect -146 -126323 -112 -126307
rect -146 -127515 -112 -127499
rect 112 -126323 146 -126307
rect 112 -127515 146 -127499
rect -100 -127583 -84 -127549
rect 84 -127583 100 -127549
rect -100 -127691 -84 -127657
rect 84 -127691 100 -127657
rect -146 -127741 -112 -127725
rect -146 -128933 -112 -128917
rect 112 -127741 146 -127725
rect 112 -128933 146 -128917
rect -100 -129001 -84 -128967
rect 84 -129001 100 -128967
rect -100 -129109 -84 -129075
rect 84 -129109 100 -129075
rect -146 -129159 -112 -129143
rect -146 -130351 -112 -130335
rect 112 -129159 146 -129143
rect 112 -130351 146 -130335
rect -100 -130419 -84 -130385
rect 84 -130419 100 -130385
rect -100 -130527 -84 -130493
rect 84 -130527 100 -130493
rect -146 -130577 -112 -130561
rect -146 -131769 -112 -131753
rect 112 -130577 146 -130561
rect 112 -131769 146 -131753
rect -100 -131837 -84 -131803
rect 84 -131837 100 -131803
rect -100 -131945 -84 -131911
rect 84 -131945 100 -131911
rect -146 -131995 -112 -131979
rect -146 -133187 -112 -133171
rect 112 -131995 146 -131979
rect 112 -133187 146 -133171
rect -100 -133255 -84 -133221
rect 84 -133255 100 -133221
rect -100 -133363 -84 -133329
rect 84 -133363 100 -133329
rect -146 -133413 -112 -133397
rect -146 -134605 -112 -134589
rect 112 -133413 146 -133397
rect 112 -134605 146 -134589
rect -100 -134673 -84 -134639
rect 84 -134673 100 -134639
rect -100 -134781 -84 -134747
rect 84 -134781 100 -134747
rect -146 -134831 -112 -134815
rect -146 -136023 -112 -136007
rect 112 -134831 146 -134815
rect 112 -136023 146 -136007
rect -100 -136091 -84 -136057
rect 84 -136091 100 -136057
rect -100 -136199 -84 -136165
rect 84 -136199 100 -136165
rect -146 -136249 -112 -136233
rect -146 -137441 -112 -137425
rect 112 -136249 146 -136233
rect 112 -137441 146 -137425
rect -100 -137509 -84 -137475
rect 84 -137509 100 -137475
rect -100 -137617 -84 -137583
rect 84 -137617 100 -137583
rect -146 -137667 -112 -137651
rect -146 -138859 -112 -138843
rect 112 -137667 146 -137651
rect 112 -138859 146 -138843
rect -100 -138927 -84 -138893
rect 84 -138927 100 -138893
rect -100 -139035 -84 -139001
rect 84 -139035 100 -139001
rect -146 -139085 -112 -139069
rect -146 -140277 -112 -140261
rect 112 -139085 146 -139069
rect 112 -140277 146 -140261
rect -100 -140345 -84 -140311
rect 84 -140345 100 -140311
rect -100 -140453 -84 -140419
rect 84 -140453 100 -140419
rect -146 -140503 -112 -140487
rect -146 -141695 -112 -141679
rect 112 -140503 146 -140487
rect 112 -141695 146 -141679
rect -100 -141763 -84 -141729
rect 84 -141763 100 -141729
rect -100 -141871 -84 -141837
rect 84 -141871 100 -141837
rect -146 -141921 -112 -141905
rect -146 -143113 -112 -143097
rect 112 -141921 146 -141905
rect 112 -143113 146 -143097
rect -100 -143181 -84 -143147
rect 84 -143181 100 -143147
rect -100 -143289 -84 -143255
rect 84 -143289 100 -143255
rect -146 -143339 -112 -143323
rect -146 -144531 -112 -144515
rect 112 -143339 146 -143323
rect 112 -144531 146 -144515
rect -100 -144599 -84 -144565
rect 84 -144599 100 -144565
rect -100 -144707 -84 -144673
rect 84 -144707 100 -144673
rect -146 -144757 -112 -144741
rect -146 -145949 -112 -145933
rect 112 -144757 146 -144741
rect 112 -145949 146 -145933
rect -100 -146017 -84 -145983
rect 84 -146017 100 -145983
rect -100 -146125 -84 -146091
rect 84 -146125 100 -146091
rect -146 -146175 -112 -146159
rect -146 -147367 -112 -147351
rect 112 -146175 146 -146159
rect 112 -147367 146 -147351
rect -100 -147435 -84 -147401
rect 84 -147435 100 -147401
rect -100 -147543 -84 -147509
rect 84 -147543 100 -147509
rect -146 -147593 -112 -147577
rect -146 -148785 -112 -148769
rect 112 -147593 146 -147577
rect 112 -148785 146 -148769
rect -100 -148853 -84 -148819
rect 84 -148853 100 -148819
rect -100 -148961 -84 -148927
rect 84 -148961 100 -148927
rect -146 -149011 -112 -148995
rect -146 -150203 -112 -150187
rect 112 -149011 146 -148995
rect 112 -150203 146 -150187
rect -100 -150271 -84 -150237
rect 84 -150271 100 -150237
rect -100 -150379 -84 -150345
rect 84 -150379 100 -150345
rect -146 -150429 -112 -150413
rect -146 -151621 -112 -151605
rect 112 -150429 146 -150413
rect 112 -151621 146 -151605
rect -100 -151689 -84 -151655
rect 84 -151689 100 -151655
rect -100 -151797 -84 -151763
rect 84 -151797 100 -151763
rect -146 -151847 -112 -151831
rect -146 -153039 -112 -153023
rect 112 -151847 146 -151831
rect 112 -153039 146 -153023
rect -100 -153107 -84 -153073
rect 84 -153107 100 -153073
rect -100 -153215 -84 -153181
rect 84 -153215 100 -153181
rect -146 -153265 -112 -153249
rect -146 -154457 -112 -154441
rect 112 -153265 146 -153249
rect 112 -154457 146 -154441
rect -100 -154525 -84 -154491
rect 84 -154525 100 -154491
rect -100 -154633 -84 -154599
rect 84 -154633 100 -154599
rect -146 -154683 -112 -154667
rect -146 -155875 -112 -155859
rect 112 -154683 146 -154667
rect 112 -155875 146 -155859
rect -100 -155943 -84 -155909
rect 84 -155943 100 -155909
rect -100 -156051 -84 -156017
rect 84 -156051 100 -156017
rect -146 -156101 -112 -156085
rect -146 -157293 -112 -157277
rect 112 -156101 146 -156085
rect 112 -157293 146 -157277
rect -100 -157361 -84 -157327
rect 84 -157361 100 -157327
rect -100 -157469 -84 -157435
rect 84 -157469 100 -157435
rect -146 -157519 -112 -157503
rect -146 -158711 -112 -158695
rect 112 -157519 146 -157503
rect 112 -158711 146 -158695
rect -100 -158779 -84 -158745
rect 84 -158779 100 -158745
rect -100 -158887 -84 -158853
rect 84 -158887 100 -158853
rect -146 -158937 -112 -158921
rect -146 -160129 -112 -160113
rect 112 -158937 146 -158921
rect 112 -160129 146 -160113
rect -100 -160197 -84 -160163
rect 84 -160197 100 -160163
rect -100 -160305 -84 -160271
rect 84 -160305 100 -160271
rect -146 -160355 -112 -160339
rect -146 -161547 -112 -161531
rect 112 -160355 146 -160339
rect 112 -161547 146 -161531
rect -100 -161615 -84 -161581
rect 84 -161615 100 -161581
rect -100 -161723 -84 -161689
rect 84 -161723 100 -161689
rect -146 -161773 -112 -161757
rect -146 -162965 -112 -162949
rect 112 -161773 146 -161757
rect 112 -162965 146 -162949
rect -100 -163033 -84 -162999
rect 84 -163033 100 -162999
rect -100 -163141 -84 -163107
rect 84 -163141 100 -163107
rect -146 -163191 -112 -163175
rect -146 -164383 -112 -164367
rect 112 -163191 146 -163175
rect 112 -164383 146 -164367
rect -100 -164451 -84 -164417
rect 84 -164451 100 -164417
rect -100 -164559 -84 -164525
rect 84 -164559 100 -164525
rect -146 -164609 -112 -164593
rect -146 -165801 -112 -165785
rect 112 -164609 146 -164593
rect 112 -165801 146 -165785
rect -100 -165869 -84 -165835
rect 84 -165869 100 -165835
rect -100 -165977 -84 -165943
rect 84 -165977 100 -165943
rect -146 -166027 -112 -166011
rect -146 -167219 -112 -167203
rect 112 -166027 146 -166011
rect 112 -167219 146 -167203
rect -100 -167287 -84 -167253
rect 84 -167287 100 -167253
rect -100 -167395 -84 -167361
rect 84 -167395 100 -167361
rect -146 -167445 -112 -167429
rect -146 -168637 -112 -168621
rect 112 -167445 146 -167429
rect 112 -168637 146 -168621
rect -100 -168705 -84 -168671
rect 84 -168705 100 -168671
rect -100 -168813 -84 -168779
rect 84 -168813 100 -168779
rect -146 -168863 -112 -168847
rect -146 -170055 -112 -170039
rect 112 -168863 146 -168847
rect 112 -170055 146 -170039
rect -100 -170123 -84 -170089
rect 84 -170123 100 -170089
rect -100 -170231 -84 -170197
rect 84 -170231 100 -170197
rect -146 -170281 -112 -170265
rect -146 -171473 -112 -171457
rect 112 -170281 146 -170265
rect 112 -171473 146 -171457
rect -100 -171541 -84 -171507
rect 84 -171541 100 -171507
rect -100 -171649 -84 -171615
rect 84 -171649 100 -171615
rect -146 -171699 -112 -171683
rect -146 -172891 -112 -172875
rect 112 -171699 146 -171683
rect 112 -172891 146 -172875
rect -100 -172959 -84 -172925
rect 84 -172959 100 -172925
rect -100 -173067 -84 -173033
rect 84 -173067 100 -173033
rect -146 -173117 -112 -173101
rect -146 -174309 -112 -174293
rect 112 -173117 146 -173101
rect 112 -174309 146 -174293
rect -100 -174377 -84 -174343
rect 84 -174377 100 -174343
rect -100 -174485 -84 -174451
rect 84 -174485 100 -174451
rect -146 -174535 -112 -174519
rect -146 -175727 -112 -175711
rect 112 -174535 146 -174519
rect 112 -175727 146 -175711
rect -100 -175795 -84 -175761
rect 84 -175795 100 -175761
rect -100 -175903 -84 -175869
rect 84 -175903 100 -175869
rect -146 -175953 -112 -175937
rect -146 -177145 -112 -177129
rect 112 -175953 146 -175937
rect 112 -177145 146 -177129
rect -100 -177213 -84 -177179
rect 84 -177213 100 -177179
rect -100 -177321 -84 -177287
rect 84 -177321 100 -177287
rect -146 -177371 -112 -177355
rect -146 -178563 -112 -178547
rect 112 -177371 146 -177355
rect 112 -178563 146 -178547
rect -100 -178631 -84 -178597
rect 84 -178631 100 -178597
rect -100 -178739 -84 -178705
rect 84 -178739 100 -178705
rect -146 -178789 -112 -178773
rect -146 -179981 -112 -179965
rect 112 -178789 146 -178773
rect 112 -179981 146 -179965
rect -100 -180049 -84 -180015
rect 84 -180049 100 -180015
rect -100 -180157 -84 -180123
rect 84 -180157 100 -180123
rect -146 -180207 -112 -180191
rect -146 -181399 -112 -181383
rect 112 -180207 146 -180191
rect 112 -181399 146 -181383
rect -100 -181467 -84 -181433
rect 84 -181467 100 -181433
rect -280 -181571 -246 -181509
rect 246 -181571 280 -181509
rect -280 -181605 -184 -181571
rect 184 -181605 280 -181571
<< viali >>
rect -84 181433 84 181467
rect -146 180207 -112 181383
rect 112 180207 146 181383
rect -84 180123 84 180157
rect -84 180015 84 180049
rect -146 178789 -112 179965
rect 112 178789 146 179965
rect -84 178705 84 178739
rect -84 178597 84 178631
rect -146 177371 -112 178547
rect 112 177371 146 178547
rect -84 177287 84 177321
rect -84 177179 84 177213
rect -146 175953 -112 177129
rect 112 175953 146 177129
rect -84 175869 84 175903
rect -84 175761 84 175795
rect -146 174535 -112 175711
rect 112 174535 146 175711
rect -84 174451 84 174485
rect -84 174343 84 174377
rect -146 173117 -112 174293
rect 112 173117 146 174293
rect -84 173033 84 173067
rect -84 172925 84 172959
rect -146 171699 -112 172875
rect 112 171699 146 172875
rect -84 171615 84 171649
rect -84 171507 84 171541
rect -146 170281 -112 171457
rect 112 170281 146 171457
rect -84 170197 84 170231
rect -84 170089 84 170123
rect -146 168863 -112 170039
rect 112 168863 146 170039
rect -84 168779 84 168813
rect -84 168671 84 168705
rect -146 167445 -112 168621
rect 112 167445 146 168621
rect -84 167361 84 167395
rect -84 167253 84 167287
rect -146 166027 -112 167203
rect 112 166027 146 167203
rect -84 165943 84 165977
rect -84 165835 84 165869
rect -146 164609 -112 165785
rect 112 164609 146 165785
rect -84 164525 84 164559
rect -84 164417 84 164451
rect -146 163191 -112 164367
rect 112 163191 146 164367
rect -84 163107 84 163141
rect -84 162999 84 163033
rect -146 161773 -112 162949
rect 112 161773 146 162949
rect -84 161689 84 161723
rect -84 161581 84 161615
rect -146 160355 -112 161531
rect 112 160355 146 161531
rect -84 160271 84 160305
rect -84 160163 84 160197
rect -146 158937 -112 160113
rect 112 158937 146 160113
rect -84 158853 84 158887
rect -84 158745 84 158779
rect -146 157519 -112 158695
rect 112 157519 146 158695
rect -84 157435 84 157469
rect -84 157327 84 157361
rect -146 156101 -112 157277
rect 112 156101 146 157277
rect -84 156017 84 156051
rect -84 155909 84 155943
rect -146 154683 -112 155859
rect 112 154683 146 155859
rect -84 154599 84 154633
rect -84 154491 84 154525
rect -146 153265 -112 154441
rect 112 153265 146 154441
rect -84 153181 84 153215
rect -84 153073 84 153107
rect -146 151847 -112 153023
rect 112 151847 146 153023
rect -84 151763 84 151797
rect -84 151655 84 151689
rect -146 150429 -112 151605
rect 112 150429 146 151605
rect -84 150345 84 150379
rect -84 150237 84 150271
rect -146 149011 -112 150187
rect 112 149011 146 150187
rect -84 148927 84 148961
rect -84 148819 84 148853
rect -146 147593 -112 148769
rect 112 147593 146 148769
rect -84 147509 84 147543
rect -84 147401 84 147435
rect -146 146175 -112 147351
rect 112 146175 146 147351
rect -84 146091 84 146125
rect -84 145983 84 146017
rect -146 144757 -112 145933
rect 112 144757 146 145933
rect -84 144673 84 144707
rect -84 144565 84 144599
rect -146 143339 -112 144515
rect 112 143339 146 144515
rect -84 143255 84 143289
rect -84 143147 84 143181
rect -146 141921 -112 143097
rect 112 141921 146 143097
rect -84 141837 84 141871
rect -84 141729 84 141763
rect -146 140503 -112 141679
rect 112 140503 146 141679
rect -84 140419 84 140453
rect -84 140311 84 140345
rect -146 139085 -112 140261
rect 112 139085 146 140261
rect -84 139001 84 139035
rect -84 138893 84 138927
rect -146 137667 -112 138843
rect 112 137667 146 138843
rect -84 137583 84 137617
rect -84 137475 84 137509
rect -146 136249 -112 137425
rect 112 136249 146 137425
rect -84 136165 84 136199
rect -84 136057 84 136091
rect -146 134831 -112 136007
rect 112 134831 146 136007
rect -84 134747 84 134781
rect -84 134639 84 134673
rect -146 133413 -112 134589
rect 112 133413 146 134589
rect -84 133329 84 133363
rect -84 133221 84 133255
rect -146 131995 -112 133171
rect 112 131995 146 133171
rect -84 131911 84 131945
rect -84 131803 84 131837
rect -146 130577 -112 131753
rect 112 130577 146 131753
rect -84 130493 84 130527
rect -84 130385 84 130419
rect -146 129159 -112 130335
rect 112 129159 146 130335
rect -84 129075 84 129109
rect -84 128967 84 129001
rect -146 127741 -112 128917
rect 112 127741 146 128917
rect -84 127657 84 127691
rect -84 127549 84 127583
rect -146 126323 -112 127499
rect 112 126323 146 127499
rect -84 126239 84 126273
rect -84 126131 84 126165
rect -146 124905 -112 126081
rect 112 124905 146 126081
rect -84 124821 84 124855
rect -84 124713 84 124747
rect -146 123487 -112 124663
rect 112 123487 146 124663
rect -84 123403 84 123437
rect -84 123295 84 123329
rect -146 122069 -112 123245
rect 112 122069 146 123245
rect -84 121985 84 122019
rect -84 121877 84 121911
rect -146 120651 -112 121827
rect 112 120651 146 121827
rect -84 120567 84 120601
rect -84 120459 84 120493
rect -146 119233 -112 120409
rect 112 119233 146 120409
rect -84 119149 84 119183
rect -84 119041 84 119075
rect -146 117815 -112 118991
rect 112 117815 146 118991
rect -84 117731 84 117765
rect -84 117623 84 117657
rect -146 116397 -112 117573
rect 112 116397 146 117573
rect -84 116313 84 116347
rect -84 116205 84 116239
rect -146 114979 -112 116155
rect 112 114979 146 116155
rect -84 114895 84 114929
rect -84 114787 84 114821
rect -146 113561 -112 114737
rect 112 113561 146 114737
rect -84 113477 84 113511
rect -84 113369 84 113403
rect -146 112143 -112 113319
rect 112 112143 146 113319
rect -84 112059 84 112093
rect -84 111951 84 111985
rect -146 110725 -112 111901
rect 112 110725 146 111901
rect -84 110641 84 110675
rect -84 110533 84 110567
rect -146 109307 -112 110483
rect 112 109307 146 110483
rect -84 109223 84 109257
rect -84 109115 84 109149
rect -146 107889 -112 109065
rect 112 107889 146 109065
rect -84 107805 84 107839
rect -84 107697 84 107731
rect -146 106471 -112 107647
rect 112 106471 146 107647
rect -84 106387 84 106421
rect -84 106279 84 106313
rect -146 105053 -112 106229
rect 112 105053 146 106229
rect -84 104969 84 105003
rect -84 104861 84 104895
rect -146 103635 -112 104811
rect 112 103635 146 104811
rect -84 103551 84 103585
rect -84 103443 84 103477
rect -146 102217 -112 103393
rect 112 102217 146 103393
rect -84 102133 84 102167
rect -84 102025 84 102059
rect -146 100799 -112 101975
rect 112 100799 146 101975
rect -84 100715 84 100749
rect -84 100607 84 100641
rect -146 99381 -112 100557
rect 112 99381 146 100557
rect -84 99297 84 99331
rect -84 99189 84 99223
rect -146 97963 -112 99139
rect 112 97963 146 99139
rect -84 97879 84 97913
rect -84 97771 84 97805
rect -146 96545 -112 97721
rect 112 96545 146 97721
rect -84 96461 84 96495
rect -84 96353 84 96387
rect -146 95127 -112 96303
rect 112 95127 146 96303
rect -84 95043 84 95077
rect -84 94935 84 94969
rect -146 93709 -112 94885
rect 112 93709 146 94885
rect -84 93625 84 93659
rect -84 93517 84 93551
rect -146 92291 -112 93467
rect 112 92291 146 93467
rect -84 92207 84 92241
rect -84 92099 84 92133
rect -146 90873 -112 92049
rect 112 90873 146 92049
rect -84 90789 84 90823
rect -84 90681 84 90715
rect -146 89455 -112 90631
rect 112 89455 146 90631
rect -84 89371 84 89405
rect -84 89263 84 89297
rect -146 88037 -112 89213
rect 112 88037 146 89213
rect -84 87953 84 87987
rect -84 87845 84 87879
rect -146 86619 -112 87795
rect 112 86619 146 87795
rect -84 86535 84 86569
rect -84 86427 84 86461
rect -146 85201 -112 86377
rect 112 85201 146 86377
rect -84 85117 84 85151
rect -84 85009 84 85043
rect -146 83783 -112 84959
rect 112 83783 146 84959
rect -84 83699 84 83733
rect -84 83591 84 83625
rect -146 82365 -112 83541
rect 112 82365 146 83541
rect -84 82281 84 82315
rect -84 82173 84 82207
rect -146 80947 -112 82123
rect 112 80947 146 82123
rect -84 80863 84 80897
rect -84 80755 84 80789
rect -146 79529 -112 80705
rect 112 79529 146 80705
rect -84 79445 84 79479
rect -84 79337 84 79371
rect -146 78111 -112 79287
rect 112 78111 146 79287
rect -84 78027 84 78061
rect -84 77919 84 77953
rect -146 76693 -112 77869
rect 112 76693 146 77869
rect -84 76609 84 76643
rect -84 76501 84 76535
rect -146 75275 -112 76451
rect 112 75275 146 76451
rect -84 75191 84 75225
rect -84 75083 84 75117
rect -146 73857 -112 75033
rect 112 73857 146 75033
rect -84 73773 84 73807
rect -84 73665 84 73699
rect -146 72439 -112 73615
rect 112 72439 146 73615
rect -84 72355 84 72389
rect -84 72247 84 72281
rect -146 71021 -112 72197
rect 112 71021 146 72197
rect -84 70937 84 70971
rect -84 70829 84 70863
rect -146 69603 -112 70779
rect 112 69603 146 70779
rect -84 69519 84 69553
rect -84 69411 84 69445
rect -146 68185 -112 69361
rect 112 68185 146 69361
rect -84 68101 84 68135
rect -84 67993 84 68027
rect -146 66767 -112 67943
rect 112 66767 146 67943
rect -84 66683 84 66717
rect -84 66575 84 66609
rect -146 65349 -112 66525
rect 112 65349 146 66525
rect -84 65265 84 65299
rect -84 65157 84 65191
rect -146 63931 -112 65107
rect 112 63931 146 65107
rect -84 63847 84 63881
rect -84 63739 84 63773
rect -146 62513 -112 63689
rect 112 62513 146 63689
rect -84 62429 84 62463
rect -84 62321 84 62355
rect -146 61095 -112 62271
rect 112 61095 146 62271
rect -84 61011 84 61045
rect -84 60903 84 60937
rect -146 59677 -112 60853
rect 112 59677 146 60853
rect -84 59593 84 59627
rect -84 59485 84 59519
rect -146 58259 -112 59435
rect 112 58259 146 59435
rect -84 58175 84 58209
rect -84 58067 84 58101
rect -146 56841 -112 58017
rect 112 56841 146 58017
rect -84 56757 84 56791
rect -84 56649 84 56683
rect -146 55423 -112 56599
rect 112 55423 146 56599
rect -84 55339 84 55373
rect -84 55231 84 55265
rect -146 54005 -112 55181
rect 112 54005 146 55181
rect -84 53921 84 53955
rect -84 53813 84 53847
rect -146 52587 -112 53763
rect 112 52587 146 53763
rect -84 52503 84 52537
rect -84 52395 84 52429
rect -146 51169 -112 52345
rect 112 51169 146 52345
rect -84 51085 84 51119
rect -84 50977 84 51011
rect -146 49751 -112 50927
rect 112 49751 146 50927
rect -84 49667 84 49701
rect -84 49559 84 49593
rect -146 48333 -112 49509
rect 112 48333 146 49509
rect -84 48249 84 48283
rect -84 48141 84 48175
rect -146 46915 -112 48091
rect 112 46915 146 48091
rect -84 46831 84 46865
rect -84 46723 84 46757
rect -146 45497 -112 46673
rect 112 45497 146 46673
rect -84 45413 84 45447
rect -84 45305 84 45339
rect -146 44079 -112 45255
rect 112 44079 146 45255
rect -84 43995 84 44029
rect -84 43887 84 43921
rect -146 42661 -112 43837
rect 112 42661 146 43837
rect -84 42577 84 42611
rect -84 42469 84 42503
rect -146 41243 -112 42419
rect 112 41243 146 42419
rect -84 41159 84 41193
rect -84 41051 84 41085
rect -146 39825 -112 41001
rect 112 39825 146 41001
rect -84 39741 84 39775
rect -84 39633 84 39667
rect -146 38407 -112 39583
rect 112 38407 146 39583
rect -84 38323 84 38357
rect -84 38215 84 38249
rect -146 36989 -112 38165
rect 112 36989 146 38165
rect -84 36905 84 36939
rect -84 36797 84 36831
rect -146 35571 -112 36747
rect 112 35571 146 36747
rect -84 35487 84 35521
rect -84 35379 84 35413
rect -146 34153 -112 35329
rect 112 34153 146 35329
rect -84 34069 84 34103
rect -84 33961 84 33995
rect -146 32735 -112 33911
rect 112 32735 146 33911
rect -84 32651 84 32685
rect -84 32543 84 32577
rect -146 31317 -112 32493
rect 112 31317 146 32493
rect -84 31233 84 31267
rect -84 31125 84 31159
rect -146 29899 -112 31075
rect 112 29899 146 31075
rect -84 29815 84 29849
rect -84 29707 84 29741
rect -146 28481 -112 29657
rect 112 28481 146 29657
rect -84 28397 84 28431
rect -84 28289 84 28323
rect -146 27063 -112 28239
rect 112 27063 146 28239
rect -84 26979 84 27013
rect -84 26871 84 26905
rect -146 25645 -112 26821
rect 112 25645 146 26821
rect -84 25561 84 25595
rect -84 25453 84 25487
rect -146 24227 -112 25403
rect 112 24227 146 25403
rect -84 24143 84 24177
rect -84 24035 84 24069
rect -146 22809 -112 23985
rect 112 22809 146 23985
rect -84 22725 84 22759
rect -84 22617 84 22651
rect -146 21391 -112 22567
rect 112 21391 146 22567
rect -84 21307 84 21341
rect -84 21199 84 21233
rect -146 19973 -112 21149
rect 112 19973 146 21149
rect -84 19889 84 19923
rect -84 19781 84 19815
rect -146 18555 -112 19731
rect 112 18555 146 19731
rect -84 18471 84 18505
rect -84 18363 84 18397
rect -146 17137 -112 18313
rect 112 17137 146 18313
rect -84 17053 84 17087
rect -84 16945 84 16979
rect -146 15719 -112 16895
rect 112 15719 146 16895
rect -84 15635 84 15669
rect -84 15527 84 15561
rect -146 14301 -112 15477
rect 112 14301 146 15477
rect -84 14217 84 14251
rect -84 14109 84 14143
rect -146 12883 -112 14059
rect 112 12883 146 14059
rect -84 12799 84 12833
rect -84 12691 84 12725
rect -146 11465 -112 12641
rect 112 11465 146 12641
rect -84 11381 84 11415
rect -84 11273 84 11307
rect -146 10047 -112 11223
rect 112 10047 146 11223
rect -84 9963 84 9997
rect -84 9855 84 9889
rect -146 8629 -112 9805
rect 112 8629 146 9805
rect -84 8545 84 8579
rect -84 8437 84 8471
rect -146 7211 -112 8387
rect 112 7211 146 8387
rect -84 7127 84 7161
rect -84 7019 84 7053
rect -146 5793 -112 6969
rect 112 5793 146 6969
rect -84 5709 84 5743
rect -84 5601 84 5635
rect -146 4375 -112 5551
rect 112 4375 146 5551
rect -84 4291 84 4325
rect -84 4183 84 4217
rect -146 2957 -112 4133
rect 112 2957 146 4133
rect -84 2873 84 2907
rect -84 2765 84 2799
rect -146 1539 -112 2715
rect 112 1539 146 2715
rect -84 1455 84 1489
rect -84 1347 84 1381
rect -146 121 -112 1297
rect 112 121 146 1297
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -1297 -112 -121
rect 112 -1297 146 -121
rect -84 -1381 84 -1347
rect -84 -1489 84 -1455
rect -146 -2715 -112 -1539
rect 112 -2715 146 -1539
rect -84 -2799 84 -2765
rect -84 -2907 84 -2873
rect -146 -4133 -112 -2957
rect 112 -4133 146 -2957
rect -84 -4217 84 -4183
rect -84 -4325 84 -4291
rect -146 -5551 -112 -4375
rect 112 -5551 146 -4375
rect -84 -5635 84 -5601
rect -84 -5743 84 -5709
rect -146 -6969 -112 -5793
rect 112 -6969 146 -5793
rect -84 -7053 84 -7019
rect -84 -7161 84 -7127
rect -146 -8387 -112 -7211
rect 112 -8387 146 -7211
rect -84 -8471 84 -8437
rect -84 -8579 84 -8545
rect -146 -9805 -112 -8629
rect 112 -9805 146 -8629
rect -84 -9889 84 -9855
rect -84 -9997 84 -9963
rect -146 -11223 -112 -10047
rect 112 -11223 146 -10047
rect -84 -11307 84 -11273
rect -84 -11415 84 -11381
rect -146 -12641 -112 -11465
rect 112 -12641 146 -11465
rect -84 -12725 84 -12691
rect -84 -12833 84 -12799
rect -146 -14059 -112 -12883
rect 112 -14059 146 -12883
rect -84 -14143 84 -14109
rect -84 -14251 84 -14217
rect -146 -15477 -112 -14301
rect 112 -15477 146 -14301
rect -84 -15561 84 -15527
rect -84 -15669 84 -15635
rect -146 -16895 -112 -15719
rect 112 -16895 146 -15719
rect -84 -16979 84 -16945
rect -84 -17087 84 -17053
rect -146 -18313 -112 -17137
rect 112 -18313 146 -17137
rect -84 -18397 84 -18363
rect -84 -18505 84 -18471
rect -146 -19731 -112 -18555
rect 112 -19731 146 -18555
rect -84 -19815 84 -19781
rect -84 -19923 84 -19889
rect -146 -21149 -112 -19973
rect 112 -21149 146 -19973
rect -84 -21233 84 -21199
rect -84 -21341 84 -21307
rect -146 -22567 -112 -21391
rect 112 -22567 146 -21391
rect -84 -22651 84 -22617
rect -84 -22759 84 -22725
rect -146 -23985 -112 -22809
rect 112 -23985 146 -22809
rect -84 -24069 84 -24035
rect -84 -24177 84 -24143
rect -146 -25403 -112 -24227
rect 112 -25403 146 -24227
rect -84 -25487 84 -25453
rect -84 -25595 84 -25561
rect -146 -26821 -112 -25645
rect 112 -26821 146 -25645
rect -84 -26905 84 -26871
rect -84 -27013 84 -26979
rect -146 -28239 -112 -27063
rect 112 -28239 146 -27063
rect -84 -28323 84 -28289
rect -84 -28431 84 -28397
rect -146 -29657 -112 -28481
rect 112 -29657 146 -28481
rect -84 -29741 84 -29707
rect -84 -29849 84 -29815
rect -146 -31075 -112 -29899
rect 112 -31075 146 -29899
rect -84 -31159 84 -31125
rect -84 -31267 84 -31233
rect -146 -32493 -112 -31317
rect 112 -32493 146 -31317
rect -84 -32577 84 -32543
rect -84 -32685 84 -32651
rect -146 -33911 -112 -32735
rect 112 -33911 146 -32735
rect -84 -33995 84 -33961
rect -84 -34103 84 -34069
rect -146 -35329 -112 -34153
rect 112 -35329 146 -34153
rect -84 -35413 84 -35379
rect -84 -35521 84 -35487
rect -146 -36747 -112 -35571
rect 112 -36747 146 -35571
rect -84 -36831 84 -36797
rect -84 -36939 84 -36905
rect -146 -38165 -112 -36989
rect 112 -38165 146 -36989
rect -84 -38249 84 -38215
rect -84 -38357 84 -38323
rect -146 -39583 -112 -38407
rect 112 -39583 146 -38407
rect -84 -39667 84 -39633
rect -84 -39775 84 -39741
rect -146 -41001 -112 -39825
rect 112 -41001 146 -39825
rect -84 -41085 84 -41051
rect -84 -41193 84 -41159
rect -146 -42419 -112 -41243
rect 112 -42419 146 -41243
rect -84 -42503 84 -42469
rect -84 -42611 84 -42577
rect -146 -43837 -112 -42661
rect 112 -43837 146 -42661
rect -84 -43921 84 -43887
rect -84 -44029 84 -43995
rect -146 -45255 -112 -44079
rect 112 -45255 146 -44079
rect -84 -45339 84 -45305
rect -84 -45447 84 -45413
rect -146 -46673 -112 -45497
rect 112 -46673 146 -45497
rect -84 -46757 84 -46723
rect -84 -46865 84 -46831
rect -146 -48091 -112 -46915
rect 112 -48091 146 -46915
rect -84 -48175 84 -48141
rect -84 -48283 84 -48249
rect -146 -49509 -112 -48333
rect 112 -49509 146 -48333
rect -84 -49593 84 -49559
rect -84 -49701 84 -49667
rect -146 -50927 -112 -49751
rect 112 -50927 146 -49751
rect -84 -51011 84 -50977
rect -84 -51119 84 -51085
rect -146 -52345 -112 -51169
rect 112 -52345 146 -51169
rect -84 -52429 84 -52395
rect -84 -52537 84 -52503
rect -146 -53763 -112 -52587
rect 112 -53763 146 -52587
rect -84 -53847 84 -53813
rect -84 -53955 84 -53921
rect -146 -55181 -112 -54005
rect 112 -55181 146 -54005
rect -84 -55265 84 -55231
rect -84 -55373 84 -55339
rect -146 -56599 -112 -55423
rect 112 -56599 146 -55423
rect -84 -56683 84 -56649
rect -84 -56791 84 -56757
rect -146 -58017 -112 -56841
rect 112 -58017 146 -56841
rect -84 -58101 84 -58067
rect -84 -58209 84 -58175
rect -146 -59435 -112 -58259
rect 112 -59435 146 -58259
rect -84 -59519 84 -59485
rect -84 -59627 84 -59593
rect -146 -60853 -112 -59677
rect 112 -60853 146 -59677
rect -84 -60937 84 -60903
rect -84 -61045 84 -61011
rect -146 -62271 -112 -61095
rect 112 -62271 146 -61095
rect -84 -62355 84 -62321
rect -84 -62463 84 -62429
rect -146 -63689 -112 -62513
rect 112 -63689 146 -62513
rect -84 -63773 84 -63739
rect -84 -63881 84 -63847
rect -146 -65107 -112 -63931
rect 112 -65107 146 -63931
rect -84 -65191 84 -65157
rect -84 -65299 84 -65265
rect -146 -66525 -112 -65349
rect 112 -66525 146 -65349
rect -84 -66609 84 -66575
rect -84 -66717 84 -66683
rect -146 -67943 -112 -66767
rect 112 -67943 146 -66767
rect -84 -68027 84 -67993
rect -84 -68135 84 -68101
rect -146 -69361 -112 -68185
rect 112 -69361 146 -68185
rect -84 -69445 84 -69411
rect -84 -69553 84 -69519
rect -146 -70779 -112 -69603
rect 112 -70779 146 -69603
rect -84 -70863 84 -70829
rect -84 -70971 84 -70937
rect -146 -72197 -112 -71021
rect 112 -72197 146 -71021
rect -84 -72281 84 -72247
rect -84 -72389 84 -72355
rect -146 -73615 -112 -72439
rect 112 -73615 146 -72439
rect -84 -73699 84 -73665
rect -84 -73807 84 -73773
rect -146 -75033 -112 -73857
rect 112 -75033 146 -73857
rect -84 -75117 84 -75083
rect -84 -75225 84 -75191
rect -146 -76451 -112 -75275
rect 112 -76451 146 -75275
rect -84 -76535 84 -76501
rect -84 -76643 84 -76609
rect -146 -77869 -112 -76693
rect 112 -77869 146 -76693
rect -84 -77953 84 -77919
rect -84 -78061 84 -78027
rect -146 -79287 -112 -78111
rect 112 -79287 146 -78111
rect -84 -79371 84 -79337
rect -84 -79479 84 -79445
rect -146 -80705 -112 -79529
rect 112 -80705 146 -79529
rect -84 -80789 84 -80755
rect -84 -80897 84 -80863
rect -146 -82123 -112 -80947
rect 112 -82123 146 -80947
rect -84 -82207 84 -82173
rect -84 -82315 84 -82281
rect -146 -83541 -112 -82365
rect 112 -83541 146 -82365
rect -84 -83625 84 -83591
rect -84 -83733 84 -83699
rect -146 -84959 -112 -83783
rect 112 -84959 146 -83783
rect -84 -85043 84 -85009
rect -84 -85151 84 -85117
rect -146 -86377 -112 -85201
rect 112 -86377 146 -85201
rect -84 -86461 84 -86427
rect -84 -86569 84 -86535
rect -146 -87795 -112 -86619
rect 112 -87795 146 -86619
rect -84 -87879 84 -87845
rect -84 -87987 84 -87953
rect -146 -89213 -112 -88037
rect 112 -89213 146 -88037
rect -84 -89297 84 -89263
rect -84 -89405 84 -89371
rect -146 -90631 -112 -89455
rect 112 -90631 146 -89455
rect -84 -90715 84 -90681
rect -84 -90823 84 -90789
rect -146 -92049 -112 -90873
rect 112 -92049 146 -90873
rect -84 -92133 84 -92099
rect -84 -92241 84 -92207
rect -146 -93467 -112 -92291
rect 112 -93467 146 -92291
rect -84 -93551 84 -93517
rect -84 -93659 84 -93625
rect -146 -94885 -112 -93709
rect 112 -94885 146 -93709
rect -84 -94969 84 -94935
rect -84 -95077 84 -95043
rect -146 -96303 -112 -95127
rect 112 -96303 146 -95127
rect -84 -96387 84 -96353
rect -84 -96495 84 -96461
rect -146 -97721 -112 -96545
rect 112 -97721 146 -96545
rect -84 -97805 84 -97771
rect -84 -97913 84 -97879
rect -146 -99139 -112 -97963
rect 112 -99139 146 -97963
rect -84 -99223 84 -99189
rect -84 -99331 84 -99297
rect -146 -100557 -112 -99381
rect 112 -100557 146 -99381
rect -84 -100641 84 -100607
rect -84 -100749 84 -100715
rect -146 -101975 -112 -100799
rect 112 -101975 146 -100799
rect -84 -102059 84 -102025
rect -84 -102167 84 -102133
rect -146 -103393 -112 -102217
rect 112 -103393 146 -102217
rect -84 -103477 84 -103443
rect -84 -103585 84 -103551
rect -146 -104811 -112 -103635
rect 112 -104811 146 -103635
rect -84 -104895 84 -104861
rect -84 -105003 84 -104969
rect -146 -106229 -112 -105053
rect 112 -106229 146 -105053
rect -84 -106313 84 -106279
rect -84 -106421 84 -106387
rect -146 -107647 -112 -106471
rect 112 -107647 146 -106471
rect -84 -107731 84 -107697
rect -84 -107839 84 -107805
rect -146 -109065 -112 -107889
rect 112 -109065 146 -107889
rect -84 -109149 84 -109115
rect -84 -109257 84 -109223
rect -146 -110483 -112 -109307
rect 112 -110483 146 -109307
rect -84 -110567 84 -110533
rect -84 -110675 84 -110641
rect -146 -111901 -112 -110725
rect 112 -111901 146 -110725
rect -84 -111985 84 -111951
rect -84 -112093 84 -112059
rect -146 -113319 -112 -112143
rect 112 -113319 146 -112143
rect -84 -113403 84 -113369
rect -84 -113511 84 -113477
rect -146 -114737 -112 -113561
rect 112 -114737 146 -113561
rect -84 -114821 84 -114787
rect -84 -114929 84 -114895
rect -146 -116155 -112 -114979
rect 112 -116155 146 -114979
rect -84 -116239 84 -116205
rect -84 -116347 84 -116313
rect -146 -117573 -112 -116397
rect 112 -117573 146 -116397
rect -84 -117657 84 -117623
rect -84 -117765 84 -117731
rect -146 -118991 -112 -117815
rect 112 -118991 146 -117815
rect -84 -119075 84 -119041
rect -84 -119183 84 -119149
rect -146 -120409 -112 -119233
rect 112 -120409 146 -119233
rect -84 -120493 84 -120459
rect -84 -120601 84 -120567
rect -146 -121827 -112 -120651
rect 112 -121827 146 -120651
rect -84 -121911 84 -121877
rect -84 -122019 84 -121985
rect -146 -123245 -112 -122069
rect 112 -123245 146 -122069
rect -84 -123329 84 -123295
rect -84 -123437 84 -123403
rect -146 -124663 -112 -123487
rect 112 -124663 146 -123487
rect -84 -124747 84 -124713
rect -84 -124855 84 -124821
rect -146 -126081 -112 -124905
rect 112 -126081 146 -124905
rect -84 -126165 84 -126131
rect -84 -126273 84 -126239
rect -146 -127499 -112 -126323
rect 112 -127499 146 -126323
rect -84 -127583 84 -127549
rect -84 -127691 84 -127657
rect -146 -128917 -112 -127741
rect 112 -128917 146 -127741
rect -84 -129001 84 -128967
rect -84 -129109 84 -129075
rect -146 -130335 -112 -129159
rect 112 -130335 146 -129159
rect -84 -130419 84 -130385
rect -84 -130527 84 -130493
rect -146 -131753 -112 -130577
rect 112 -131753 146 -130577
rect -84 -131837 84 -131803
rect -84 -131945 84 -131911
rect -146 -133171 -112 -131995
rect 112 -133171 146 -131995
rect -84 -133255 84 -133221
rect -84 -133363 84 -133329
rect -146 -134589 -112 -133413
rect 112 -134589 146 -133413
rect -84 -134673 84 -134639
rect -84 -134781 84 -134747
rect -146 -136007 -112 -134831
rect 112 -136007 146 -134831
rect -84 -136091 84 -136057
rect -84 -136199 84 -136165
rect -146 -137425 -112 -136249
rect 112 -137425 146 -136249
rect -84 -137509 84 -137475
rect -84 -137617 84 -137583
rect -146 -138843 -112 -137667
rect 112 -138843 146 -137667
rect -84 -138927 84 -138893
rect -84 -139035 84 -139001
rect -146 -140261 -112 -139085
rect 112 -140261 146 -139085
rect -84 -140345 84 -140311
rect -84 -140453 84 -140419
rect -146 -141679 -112 -140503
rect 112 -141679 146 -140503
rect -84 -141763 84 -141729
rect -84 -141871 84 -141837
rect -146 -143097 -112 -141921
rect 112 -143097 146 -141921
rect -84 -143181 84 -143147
rect -84 -143289 84 -143255
rect -146 -144515 -112 -143339
rect 112 -144515 146 -143339
rect -84 -144599 84 -144565
rect -84 -144707 84 -144673
rect -146 -145933 -112 -144757
rect 112 -145933 146 -144757
rect -84 -146017 84 -145983
rect -84 -146125 84 -146091
rect -146 -147351 -112 -146175
rect 112 -147351 146 -146175
rect -84 -147435 84 -147401
rect -84 -147543 84 -147509
rect -146 -148769 -112 -147593
rect 112 -148769 146 -147593
rect -84 -148853 84 -148819
rect -84 -148961 84 -148927
rect -146 -150187 -112 -149011
rect 112 -150187 146 -149011
rect -84 -150271 84 -150237
rect -84 -150379 84 -150345
rect -146 -151605 -112 -150429
rect 112 -151605 146 -150429
rect -84 -151689 84 -151655
rect -84 -151797 84 -151763
rect -146 -153023 -112 -151847
rect 112 -153023 146 -151847
rect -84 -153107 84 -153073
rect -84 -153215 84 -153181
rect -146 -154441 -112 -153265
rect 112 -154441 146 -153265
rect -84 -154525 84 -154491
rect -84 -154633 84 -154599
rect -146 -155859 -112 -154683
rect 112 -155859 146 -154683
rect -84 -155943 84 -155909
rect -84 -156051 84 -156017
rect -146 -157277 -112 -156101
rect 112 -157277 146 -156101
rect -84 -157361 84 -157327
rect -84 -157469 84 -157435
rect -146 -158695 -112 -157519
rect 112 -158695 146 -157519
rect -84 -158779 84 -158745
rect -84 -158887 84 -158853
rect -146 -160113 -112 -158937
rect 112 -160113 146 -158937
rect -84 -160197 84 -160163
rect -84 -160305 84 -160271
rect -146 -161531 -112 -160355
rect 112 -161531 146 -160355
rect -84 -161615 84 -161581
rect -84 -161723 84 -161689
rect -146 -162949 -112 -161773
rect 112 -162949 146 -161773
rect -84 -163033 84 -162999
rect -84 -163141 84 -163107
rect -146 -164367 -112 -163191
rect 112 -164367 146 -163191
rect -84 -164451 84 -164417
rect -84 -164559 84 -164525
rect -146 -165785 -112 -164609
rect 112 -165785 146 -164609
rect -84 -165869 84 -165835
rect -84 -165977 84 -165943
rect -146 -167203 -112 -166027
rect 112 -167203 146 -166027
rect -84 -167287 84 -167253
rect -84 -167395 84 -167361
rect -146 -168621 -112 -167445
rect 112 -168621 146 -167445
rect -84 -168705 84 -168671
rect -84 -168813 84 -168779
rect -146 -170039 -112 -168863
rect 112 -170039 146 -168863
rect -84 -170123 84 -170089
rect -84 -170231 84 -170197
rect -146 -171457 -112 -170281
rect 112 -171457 146 -170281
rect -84 -171541 84 -171507
rect -84 -171649 84 -171615
rect -146 -172875 -112 -171699
rect 112 -172875 146 -171699
rect -84 -172959 84 -172925
rect -84 -173067 84 -173033
rect -146 -174293 -112 -173117
rect 112 -174293 146 -173117
rect -84 -174377 84 -174343
rect -84 -174485 84 -174451
rect -146 -175711 -112 -174535
rect 112 -175711 146 -174535
rect -84 -175795 84 -175761
rect -84 -175903 84 -175869
rect -146 -177129 -112 -175953
rect 112 -177129 146 -175953
rect -84 -177213 84 -177179
rect -84 -177321 84 -177287
rect -146 -178547 -112 -177371
rect 112 -178547 146 -177371
rect -84 -178631 84 -178597
rect -84 -178739 84 -178705
rect -146 -179965 -112 -178789
rect 112 -179965 146 -178789
rect -84 -180049 84 -180015
rect -84 -180157 84 -180123
rect -146 -181383 -112 -180207
rect 112 -181383 146 -180207
rect -84 -181467 84 -181433
<< metal1 >>
rect -96 181467 96 181473
rect -96 181433 -84 181467
rect 84 181433 96 181467
rect -96 181427 96 181433
rect -152 181383 -106 181395
rect -152 180207 -146 181383
rect -112 180207 -106 181383
rect -152 180195 -106 180207
rect 106 181383 152 181395
rect 106 180207 112 181383
rect 146 180207 152 181383
rect 106 180195 152 180207
rect -96 180157 96 180163
rect -96 180123 -84 180157
rect 84 180123 96 180157
rect -96 180117 96 180123
rect -96 180049 96 180055
rect -96 180015 -84 180049
rect 84 180015 96 180049
rect -96 180009 96 180015
rect -152 179965 -106 179977
rect -152 178789 -146 179965
rect -112 178789 -106 179965
rect -152 178777 -106 178789
rect 106 179965 152 179977
rect 106 178789 112 179965
rect 146 178789 152 179965
rect 106 178777 152 178789
rect -96 178739 96 178745
rect -96 178705 -84 178739
rect 84 178705 96 178739
rect -96 178699 96 178705
rect -96 178631 96 178637
rect -96 178597 -84 178631
rect 84 178597 96 178631
rect -96 178591 96 178597
rect -152 178547 -106 178559
rect -152 177371 -146 178547
rect -112 177371 -106 178547
rect -152 177359 -106 177371
rect 106 178547 152 178559
rect 106 177371 112 178547
rect 146 177371 152 178547
rect 106 177359 152 177371
rect -96 177321 96 177327
rect -96 177287 -84 177321
rect 84 177287 96 177321
rect -96 177281 96 177287
rect -96 177213 96 177219
rect -96 177179 -84 177213
rect 84 177179 96 177213
rect -96 177173 96 177179
rect -152 177129 -106 177141
rect -152 175953 -146 177129
rect -112 175953 -106 177129
rect -152 175941 -106 175953
rect 106 177129 152 177141
rect 106 175953 112 177129
rect 146 175953 152 177129
rect 106 175941 152 175953
rect -96 175903 96 175909
rect -96 175869 -84 175903
rect 84 175869 96 175903
rect -96 175863 96 175869
rect -96 175795 96 175801
rect -96 175761 -84 175795
rect 84 175761 96 175795
rect -96 175755 96 175761
rect -152 175711 -106 175723
rect -152 174535 -146 175711
rect -112 174535 -106 175711
rect -152 174523 -106 174535
rect 106 175711 152 175723
rect 106 174535 112 175711
rect 146 174535 152 175711
rect 106 174523 152 174535
rect -96 174485 96 174491
rect -96 174451 -84 174485
rect 84 174451 96 174485
rect -96 174445 96 174451
rect -96 174377 96 174383
rect -96 174343 -84 174377
rect 84 174343 96 174377
rect -96 174337 96 174343
rect -152 174293 -106 174305
rect -152 173117 -146 174293
rect -112 173117 -106 174293
rect -152 173105 -106 173117
rect 106 174293 152 174305
rect 106 173117 112 174293
rect 146 173117 152 174293
rect 106 173105 152 173117
rect -96 173067 96 173073
rect -96 173033 -84 173067
rect 84 173033 96 173067
rect -96 173027 96 173033
rect -96 172959 96 172965
rect -96 172925 -84 172959
rect 84 172925 96 172959
rect -96 172919 96 172925
rect -152 172875 -106 172887
rect -152 171699 -146 172875
rect -112 171699 -106 172875
rect -152 171687 -106 171699
rect 106 172875 152 172887
rect 106 171699 112 172875
rect 146 171699 152 172875
rect 106 171687 152 171699
rect -96 171649 96 171655
rect -96 171615 -84 171649
rect 84 171615 96 171649
rect -96 171609 96 171615
rect -96 171541 96 171547
rect -96 171507 -84 171541
rect 84 171507 96 171541
rect -96 171501 96 171507
rect -152 171457 -106 171469
rect -152 170281 -146 171457
rect -112 170281 -106 171457
rect -152 170269 -106 170281
rect 106 171457 152 171469
rect 106 170281 112 171457
rect 146 170281 152 171457
rect 106 170269 152 170281
rect -96 170231 96 170237
rect -96 170197 -84 170231
rect 84 170197 96 170231
rect -96 170191 96 170197
rect -96 170123 96 170129
rect -96 170089 -84 170123
rect 84 170089 96 170123
rect -96 170083 96 170089
rect -152 170039 -106 170051
rect -152 168863 -146 170039
rect -112 168863 -106 170039
rect -152 168851 -106 168863
rect 106 170039 152 170051
rect 106 168863 112 170039
rect 146 168863 152 170039
rect 106 168851 152 168863
rect -96 168813 96 168819
rect -96 168779 -84 168813
rect 84 168779 96 168813
rect -96 168773 96 168779
rect -96 168705 96 168711
rect -96 168671 -84 168705
rect 84 168671 96 168705
rect -96 168665 96 168671
rect -152 168621 -106 168633
rect -152 167445 -146 168621
rect -112 167445 -106 168621
rect -152 167433 -106 167445
rect 106 168621 152 168633
rect 106 167445 112 168621
rect 146 167445 152 168621
rect 106 167433 152 167445
rect -96 167395 96 167401
rect -96 167361 -84 167395
rect 84 167361 96 167395
rect -96 167355 96 167361
rect -96 167287 96 167293
rect -96 167253 -84 167287
rect 84 167253 96 167287
rect -96 167247 96 167253
rect -152 167203 -106 167215
rect -152 166027 -146 167203
rect -112 166027 -106 167203
rect -152 166015 -106 166027
rect 106 167203 152 167215
rect 106 166027 112 167203
rect 146 166027 152 167203
rect 106 166015 152 166027
rect -96 165977 96 165983
rect -96 165943 -84 165977
rect 84 165943 96 165977
rect -96 165937 96 165943
rect -96 165869 96 165875
rect -96 165835 -84 165869
rect 84 165835 96 165869
rect -96 165829 96 165835
rect -152 165785 -106 165797
rect -152 164609 -146 165785
rect -112 164609 -106 165785
rect -152 164597 -106 164609
rect 106 165785 152 165797
rect 106 164609 112 165785
rect 146 164609 152 165785
rect 106 164597 152 164609
rect -96 164559 96 164565
rect -96 164525 -84 164559
rect 84 164525 96 164559
rect -96 164519 96 164525
rect -96 164451 96 164457
rect -96 164417 -84 164451
rect 84 164417 96 164451
rect -96 164411 96 164417
rect -152 164367 -106 164379
rect -152 163191 -146 164367
rect -112 163191 -106 164367
rect -152 163179 -106 163191
rect 106 164367 152 164379
rect 106 163191 112 164367
rect 146 163191 152 164367
rect 106 163179 152 163191
rect -96 163141 96 163147
rect -96 163107 -84 163141
rect 84 163107 96 163141
rect -96 163101 96 163107
rect -96 163033 96 163039
rect -96 162999 -84 163033
rect 84 162999 96 163033
rect -96 162993 96 162999
rect -152 162949 -106 162961
rect -152 161773 -146 162949
rect -112 161773 -106 162949
rect -152 161761 -106 161773
rect 106 162949 152 162961
rect 106 161773 112 162949
rect 146 161773 152 162949
rect 106 161761 152 161773
rect -96 161723 96 161729
rect -96 161689 -84 161723
rect 84 161689 96 161723
rect -96 161683 96 161689
rect -96 161615 96 161621
rect -96 161581 -84 161615
rect 84 161581 96 161615
rect -96 161575 96 161581
rect -152 161531 -106 161543
rect -152 160355 -146 161531
rect -112 160355 -106 161531
rect -152 160343 -106 160355
rect 106 161531 152 161543
rect 106 160355 112 161531
rect 146 160355 152 161531
rect 106 160343 152 160355
rect -96 160305 96 160311
rect -96 160271 -84 160305
rect 84 160271 96 160305
rect -96 160265 96 160271
rect -96 160197 96 160203
rect -96 160163 -84 160197
rect 84 160163 96 160197
rect -96 160157 96 160163
rect -152 160113 -106 160125
rect -152 158937 -146 160113
rect -112 158937 -106 160113
rect -152 158925 -106 158937
rect 106 160113 152 160125
rect 106 158937 112 160113
rect 146 158937 152 160113
rect 106 158925 152 158937
rect -96 158887 96 158893
rect -96 158853 -84 158887
rect 84 158853 96 158887
rect -96 158847 96 158853
rect -96 158779 96 158785
rect -96 158745 -84 158779
rect 84 158745 96 158779
rect -96 158739 96 158745
rect -152 158695 -106 158707
rect -152 157519 -146 158695
rect -112 157519 -106 158695
rect -152 157507 -106 157519
rect 106 158695 152 158707
rect 106 157519 112 158695
rect 146 157519 152 158695
rect 106 157507 152 157519
rect -96 157469 96 157475
rect -96 157435 -84 157469
rect 84 157435 96 157469
rect -96 157429 96 157435
rect -96 157361 96 157367
rect -96 157327 -84 157361
rect 84 157327 96 157361
rect -96 157321 96 157327
rect -152 157277 -106 157289
rect -152 156101 -146 157277
rect -112 156101 -106 157277
rect -152 156089 -106 156101
rect 106 157277 152 157289
rect 106 156101 112 157277
rect 146 156101 152 157277
rect 106 156089 152 156101
rect -96 156051 96 156057
rect -96 156017 -84 156051
rect 84 156017 96 156051
rect -96 156011 96 156017
rect -96 155943 96 155949
rect -96 155909 -84 155943
rect 84 155909 96 155943
rect -96 155903 96 155909
rect -152 155859 -106 155871
rect -152 154683 -146 155859
rect -112 154683 -106 155859
rect -152 154671 -106 154683
rect 106 155859 152 155871
rect 106 154683 112 155859
rect 146 154683 152 155859
rect 106 154671 152 154683
rect -96 154633 96 154639
rect -96 154599 -84 154633
rect 84 154599 96 154633
rect -96 154593 96 154599
rect -96 154525 96 154531
rect -96 154491 -84 154525
rect 84 154491 96 154525
rect -96 154485 96 154491
rect -152 154441 -106 154453
rect -152 153265 -146 154441
rect -112 153265 -106 154441
rect -152 153253 -106 153265
rect 106 154441 152 154453
rect 106 153265 112 154441
rect 146 153265 152 154441
rect 106 153253 152 153265
rect -96 153215 96 153221
rect -96 153181 -84 153215
rect 84 153181 96 153215
rect -96 153175 96 153181
rect -96 153107 96 153113
rect -96 153073 -84 153107
rect 84 153073 96 153107
rect -96 153067 96 153073
rect -152 153023 -106 153035
rect -152 151847 -146 153023
rect -112 151847 -106 153023
rect -152 151835 -106 151847
rect 106 153023 152 153035
rect 106 151847 112 153023
rect 146 151847 152 153023
rect 106 151835 152 151847
rect -96 151797 96 151803
rect -96 151763 -84 151797
rect 84 151763 96 151797
rect -96 151757 96 151763
rect -96 151689 96 151695
rect -96 151655 -84 151689
rect 84 151655 96 151689
rect -96 151649 96 151655
rect -152 151605 -106 151617
rect -152 150429 -146 151605
rect -112 150429 -106 151605
rect -152 150417 -106 150429
rect 106 151605 152 151617
rect 106 150429 112 151605
rect 146 150429 152 151605
rect 106 150417 152 150429
rect -96 150379 96 150385
rect -96 150345 -84 150379
rect 84 150345 96 150379
rect -96 150339 96 150345
rect -96 150271 96 150277
rect -96 150237 -84 150271
rect 84 150237 96 150271
rect -96 150231 96 150237
rect -152 150187 -106 150199
rect -152 149011 -146 150187
rect -112 149011 -106 150187
rect -152 148999 -106 149011
rect 106 150187 152 150199
rect 106 149011 112 150187
rect 146 149011 152 150187
rect 106 148999 152 149011
rect -96 148961 96 148967
rect -96 148927 -84 148961
rect 84 148927 96 148961
rect -96 148921 96 148927
rect -96 148853 96 148859
rect -96 148819 -84 148853
rect 84 148819 96 148853
rect -96 148813 96 148819
rect -152 148769 -106 148781
rect -152 147593 -146 148769
rect -112 147593 -106 148769
rect -152 147581 -106 147593
rect 106 148769 152 148781
rect 106 147593 112 148769
rect 146 147593 152 148769
rect 106 147581 152 147593
rect -96 147543 96 147549
rect -96 147509 -84 147543
rect 84 147509 96 147543
rect -96 147503 96 147509
rect -96 147435 96 147441
rect -96 147401 -84 147435
rect 84 147401 96 147435
rect -96 147395 96 147401
rect -152 147351 -106 147363
rect -152 146175 -146 147351
rect -112 146175 -106 147351
rect -152 146163 -106 146175
rect 106 147351 152 147363
rect 106 146175 112 147351
rect 146 146175 152 147351
rect 106 146163 152 146175
rect -96 146125 96 146131
rect -96 146091 -84 146125
rect 84 146091 96 146125
rect -96 146085 96 146091
rect -96 146017 96 146023
rect -96 145983 -84 146017
rect 84 145983 96 146017
rect -96 145977 96 145983
rect -152 145933 -106 145945
rect -152 144757 -146 145933
rect -112 144757 -106 145933
rect -152 144745 -106 144757
rect 106 145933 152 145945
rect 106 144757 112 145933
rect 146 144757 152 145933
rect 106 144745 152 144757
rect -96 144707 96 144713
rect -96 144673 -84 144707
rect 84 144673 96 144707
rect -96 144667 96 144673
rect -96 144599 96 144605
rect -96 144565 -84 144599
rect 84 144565 96 144599
rect -96 144559 96 144565
rect -152 144515 -106 144527
rect -152 143339 -146 144515
rect -112 143339 -106 144515
rect -152 143327 -106 143339
rect 106 144515 152 144527
rect 106 143339 112 144515
rect 146 143339 152 144515
rect 106 143327 152 143339
rect -96 143289 96 143295
rect -96 143255 -84 143289
rect 84 143255 96 143289
rect -96 143249 96 143255
rect -96 143181 96 143187
rect -96 143147 -84 143181
rect 84 143147 96 143181
rect -96 143141 96 143147
rect -152 143097 -106 143109
rect -152 141921 -146 143097
rect -112 141921 -106 143097
rect -152 141909 -106 141921
rect 106 143097 152 143109
rect 106 141921 112 143097
rect 146 141921 152 143097
rect 106 141909 152 141921
rect -96 141871 96 141877
rect -96 141837 -84 141871
rect 84 141837 96 141871
rect -96 141831 96 141837
rect -96 141763 96 141769
rect -96 141729 -84 141763
rect 84 141729 96 141763
rect -96 141723 96 141729
rect -152 141679 -106 141691
rect -152 140503 -146 141679
rect -112 140503 -106 141679
rect -152 140491 -106 140503
rect 106 141679 152 141691
rect 106 140503 112 141679
rect 146 140503 152 141679
rect 106 140491 152 140503
rect -96 140453 96 140459
rect -96 140419 -84 140453
rect 84 140419 96 140453
rect -96 140413 96 140419
rect -96 140345 96 140351
rect -96 140311 -84 140345
rect 84 140311 96 140345
rect -96 140305 96 140311
rect -152 140261 -106 140273
rect -152 139085 -146 140261
rect -112 139085 -106 140261
rect -152 139073 -106 139085
rect 106 140261 152 140273
rect 106 139085 112 140261
rect 146 139085 152 140261
rect 106 139073 152 139085
rect -96 139035 96 139041
rect -96 139001 -84 139035
rect 84 139001 96 139035
rect -96 138995 96 139001
rect -96 138927 96 138933
rect -96 138893 -84 138927
rect 84 138893 96 138927
rect -96 138887 96 138893
rect -152 138843 -106 138855
rect -152 137667 -146 138843
rect -112 137667 -106 138843
rect -152 137655 -106 137667
rect 106 138843 152 138855
rect 106 137667 112 138843
rect 146 137667 152 138843
rect 106 137655 152 137667
rect -96 137617 96 137623
rect -96 137583 -84 137617
rect 84 137583 96 137617
rect -96 137577 96 137583
rect -96 137509 96 137515
rect -96 137475 -84 137509
rect 84 137475 96 137509
rect -96 137469 96 137475
rect -152 137425 -106 137437
rect -152 136249 -146 137425
rect -112 136249 -106 137425
rect -152 136237 -106 136249
rect 106 137425 152 137437
rect 106 136249 112 137425
rect 146 136249 152 137425
rect 106 136237 152 136249
rect -96 136199 96 136205
rect -96 136165 -84 136199
rect 84 136165 96 136199
rect -96 136159 96 136165
rect -96 136091 96 136097
rect -96 136057 -84 136091
rect 84 136057 96 136091
rect -96 136051 96 136057
rect -152 136007 -106 136019
rect -152 134831 -146 136007
rect -112 134831 -106 136007
rect -152 134819 -106 134831
rect 106 136007 152 136019
rect 106 134831 112 136007
rect 146 134831 152 136007
rect 106 134819 152 134831
rect -96 134781 96 134787
rect -96 134747 -84 134781
rect 84 134747 96 134781
rect -96 134741 96 134747
rect -96 134673 96 134679
rect -96 134639 -84 134673
rect 84 134639 96 134673
rect -96 134633 96 134639
rect -152 134589 -106 134601
rect -152 133413 -146 134589
rect -112 133413 -106 134589
rect -152 133401 -106 133413
rect 106 134589 152 134601
rect 106 133413 112 134589
rect 146 133413 152 134589
rect 106 133401 152 133413
rect -96 133363 96 133369
rect -96 133329 -84 133363
rect 84 133329 96 133363
rect -96 133323 96 133329
rect -96 133255 96 133261
rect -96 133221 -84 133255
rect 84 133221 96 133255
rect -96 133215 96 133221
rect -152 133171 -106 133183
rect -152 131995 -146 133171
rect -112 131995 -106 133171
rect -152 131983 -106 131995
rect 106 133171 152 133183
rect 106 131995 112 133171
rect 146 131995 152 133171
rect 106 131983 152 131995
rect -96 131945 96 131951
rect -96 131911 -84 131945
rect 84 131911 96 131945
rect -96 131905 96 131911
rect -96 131837 96 131843
rect -96 131803 -84 131837
rect 84 131803 96 131837
rect -96 131797 96 131803
rect -152 131753 -106 131765
rect -152 130577 -146 131753
rect -112 130577 -106 131753
rect -152 130565 -106 130577
rect 106 131753 152 131765
rect 106 130577 112 131753
rect 146 130577 152 131753
rect 106 130565 152 130577
rect -96 130527 96 130533
rect -96 130493 -84 130527
rect 84 130493 96 130527
rect -96 130487 96 130493
rect -96 130419 96 130425
rect -96 130385 -84 130419
rect 84 130385 96 130419
rect -96 130379 96 130385
rect -152 130335 -106 130347
rect -152 129159 -146 130335
rect -112 129159 -106 130335
rect -152 129147 -106 129159
rect 106 130335 152 130347
rect 106 129159 112 130335
rect 146 129159 152 130335
rect 106 129147 152 129159
rect -96 129109 96 129115
rect -96 129075 -84 129109
rect 84 129075 96 129109
rect -96 129069 96 129075
rect -96 129001 96 129007
rect -96 128967 -84 129001
rect 84 128967 96 129001
rect -96 128961 96 128967
rect -152 128917 -106 128929
rect -152 127741 -146 128917
rect -112 127741 -106 128917
rect -152 127729 -106 127741
rect 106 128917 152 128929
rect 106 127741 112 128917
rect 146 127741 152 128917
rect 106 127729 152 127741
rect -96 127691 96 127697
rect -96 127657 -84 127691
rect 84 127657 96 127691
rect -96 127651 96 127657
rect -96 127583 96 127589
rect -96 127549 -84 127583
rect 84 127549 96 127583
rect -96 127543 96 127549
rect -152 127499 -106 127511
rect -152 126323 -146 127499
rect -112 126323 -106 127499
rect -152 126311 -106 126323
rect 106 127499 152 127511
rect 106 126323 112 127499
rect 146 126323 152 127499
rect 106 126311 152 126323
rect -96 126273 96 126279
rect -96 126239 -84 126273
rect 84 126239 96 126273
rect -96 126233 96 126239
rect -96 126165 96 126171
rect -96 126131 -84 126165
rect 84 126131 96 126165
rect -96 126125 96 126131
rect -152 126081 -106 126093
rect -152 124905 -146 126081
rect -112 124905 -106 126081
rect -152 124893 -106 124905
rect 106 126081 152 126093
rect 106 124905 112 126081
rect 146 124905 152 126081
rect 106 124893 152 124905
rect -96 124855 96 124861
rect -96 124821 -84 124855
rect 84 124821 96 124855
rect -96 124815 96 124821
rect -96 124747 96 124753
rect -96 124713 -84 124747
rect 84 124713 96 124747
rect -96 124707 96 124713
rect -152 124663 -106 124675
rect -152 123487 -146 124663
rect -112 123487 -106 124663
rect -152 123475 -106 123487
rect 106 124663 152 124675
rect 106 123487 112 124663
rect 146 123487 152 124663
rect 106 123475 152 123487
rect -96 123437 96 123443
rect -96 123403 -84 123437
rect 84 123403 96 123437
rect -96 123397 96 123403
rect -96 123329 96 123335
rect -96 123295 -84 123329
rect 84 123295 96 123329
rect -96 123289 96 123295
rect -152 123245 -106 123257
rect -152 122069 -146 123245
rect -112 122069 -106 123245
rect -152 122057 -106 122069
rect 106 123245 152 123257
rect 106 122069 112 123245
rect 146 122069 152 123245
rect 106 122057 152 122069
rect -96 122019 96 122025
rect -96 121985 -84 122019
rect 84 121985 96 122019
rect -96 121979 96 121985
rect -96 121911 96 121917
rect -96 121877 -84 121911
rect 84 121877 96 121911
rect -96 121871 96 121877
rect -152 121827 -106 121839
rect -152 120651 -146 121827
rect -112 120651 -106 121827
rect -152 120639 -106 120651
rect 106 121827 152 121839
rect 106 120651 112 121827
rect 146 120651 152 121827
rect 106 120639 152 120651
rect -96 120601 96 120607
rect -96 120567 -84 120601
rect 84 120567 96 120601
rect -96 120561 96 120567
rect -96 120493 96 120499
rect -96 120459 -84 120493
rect 84 120459 96 120493
rect -96 120453 96 120459
rect -152 120409 -106 120421
rect -152 119233 -146 120409
rect -112 119233 -106 120409
rect -152 119221 -106 119233
rect 106 120409 152 120421
rect 106 119233 112 120409
rect 146 119233 152 120409
rect 106 119221 152 119233
rect -96 119183 96 119189
rect -96 119149 -84 119183
rect 84 119149 96 119183
rect -96 119143 96 119149
rect -96 119075 96 119081
rect -96 119041 -84 119075
rect 84 119041 96 119075
rect -96 119035 96 119041
rect -152 118991 -106 119003
rect -152 117815 -146 118991
rect -112 117815 -106 118991
rect -152 117803 -106 117815
rect 106 118991 152 119003
rect 106 117815 112 118991
rect 146 117815 152 118991
rect 106 117803 152 117815
rect -96 117765 96 117771
rect -96 117731 -84 117765
rect 84 117731 96 117765
rect -96 117725 96 117731
rect -96 117657 96 117663
rect -96 117623 -84 117657
rect 84 117623 96 117657
rect -96 117617 96 117623
rect -152 117573 -106 117585
rect -152 116397 -146 117573
rect -112 116397 -106 117573
rect -152 116385 -106 116397
rect 106 117573 152 117585
rect 106 116397 112 117573
rect 146 116397 152 117573
rect 106 116385 152 116397
rect -96 116347 96 116353
rect -96 116313 -84 116347
rect 84 116313 96 116347
rect -96 116307 96 116313
rect -96 116239 96 116245
rect -96 116205 -84 116239
rect 84 116205 96 116239
rect -96 116199 96 116205
rect -152 116155 -106 116167
rect -152 114979 -146 116155
rect -112 114979 -106 116155
rect -152 114967 -106 114979
rect 106 116155 152 116167
rect 106 114979 112 116155
rect 146 114979 152 116155
rect 106 114967 152 114979
rect -96 114929 96 114935
rect -96 114895 -84 114929
rect 84 114895 96 114929
rect -96 114889 96 114895
rect -96 114821 96 114827
rect -96 114787 -84 114821
rect 84 114787 96 114821
rect -96 114781 96 114787
rect -152 114737 -106 114749
rect -152 113561 -146 114737
rect -112 113561 -106 114737
rect -152 113549 -106 113561
rect 106 114737 152 114749
rect 106 113561 112 114737
rect 146 113561 152 114737
rect 106 113549 152 113561
rect -96 113511 96 113517
rect -96 113477 -84 113511
rect 84 113477 96 113511
rect -96 113471 96 113477
rect -96 113403 96 113409
rect -96 113369 -84 113403
rect 84 113369 96 113403
rect -96 113363 96 113369
rect -152 113319 -106 113331
rect -152 112143 -146 113319
rect -112 112143 -106 113319
rect -152 112131 -106 112143
rect 106 113319 152 113331
rect 106 112143 112 113319
rect 146 112143 152 113319
rect 106 112131 152 112143
rect -96 112093 96 112099
rect -96 112059 -84 112093
rect 84 112059 96 112093
rect -96 112053 96 112059
rect -96 111985 96 111991
rect -96 111951 -84 111985
rect 84 111951 96 111985
rect -96 111945 96 111951
rect -152 111901 -106 111913
rect -152 110725 -146 111901
rect -112 110725 -106 111901
rect -152 110713 -106 110725
rect 106 111901 152 111913
rect 106 110725 112 111901
rect 146 110725 152 111901
rect 106 110713 152 110725
rect -96 110675 96 110681
rect -96 110641 -84 110675
rect 84 110641 96 110675
rect -96 110635 96 110641
rect -96 110567 96 110573
rect -96 110533 -84 110567
rect 84 110533 96 110567
rect -96 110527 96 110533
rect -152 110483 -106 110495
rect -152 109307 -146 110483
rect -112 109307 -106 110483
rect -152 109295 -106 109307
rect 106 110483 152 110495
rect 106 109307 112 110483
rect 146 109307 152 110483
rect 106 109295 152 109307
rect -96 109257 96 109263
rect -96 109223 -84 109257
rect 84 109223 96 109257
rect -96 109217 96 109223
rect -96 109149 96 109155
rect -96 109115 -84 109149
rect 84 109115 96 109149
rect -96 109109 96 109115
rect -152 109065 -106 109077
rect -152 107889 -146 109065
rect -112 107889 -106 109065
rect -152 107877 -106 107889
rect 106 109065 152 109077
rect 106 107889 112 109065
rect 146 107889 152 109065
rect 106 107877 152 107889
rect -96 107839 96 107845
rect -96 107805 -84 107839
rect 84 107805 96 107839
rect -96 107799 96 107805
rect -96 107731 96 107737
rect -96 107697 -84 107731
rect 84 107697 96 107731
rect -96 107691 96 107697
rect -152 107647 -106 107659
rect -152 106471 -146 107647
rect -112 106471 -106 107647
rect -152 106459 -106 106471
rect 106 107647 152 107659
rect 106 106471 112 107647
rect 146 106471 152 107647
rect 106 106459 152 106471
rect -96 106421 96 106427
rect -96 106387 -84 106421
rect 84 106387 96 106421
rect -96 106381 96 106387
rect -96 106313 96 106319
rect -96 106279 -84 106313
rect 84 106279 96 106313
rect -96 106273 96 106279
rect -152 106229 -106 106241
rect -152 105053 -146 106229
rect -112 105053 -106 106229
rect -152 105041 -106 105053
rect 106 106229 152 106241
rect 106 105053 112 106229
rect 146 105053 152 106229
rect 106 105041 152 105053
rect -96 105003 96 105009
rect -96 104969 -84 105003
rect 84 104969 96 105003
rect -96 104963 96 104969
rect -96 104895 96 104901
rect -96 104861 -84 104895
rect 84 104861 96 104895
rect -96 104855 96 104861
rect -152 104811 -106 104823
rect -152 103635 -146 104811
rect -112 103635 -106 104811
rect -152 103623 -106 103635
rect 106 104811 152 104823
rect 106 103635 112 104811
rect 146 103635 152 104811
rect 106 103623 152 103635
rect -96 103585 96 103591
rect -96 103551 -84 103585
rect 84 103551 96 103585
rect -96 103545 96 103551
rect -96 103477 96 103483
rect -96 103443 -84 103477
rect 84 103443 96 103477
rect -96 103437 96 103443
rect -152 103393 -106 103405
rect -152 102217 -146 103393
rect -112 102217 -106 103393
rect -152 102205 -106 102217
rect 106 103393 152 103405
rect 106 102217 112 103393
rect 146 102217 152 103393
rect 106 102205 152 102217
rect -96 102167 96 102173
rect -96 102133 -84 102167
rect 84 102133 96 102167
rect -96 102127 96 102133
rect -96 102059 96 102065
rect -96 102025 -84 102059
rect 84 102025 96 102059
rect -96 102019 96 102025
rect -152 101975 -106 101987
rect -152 100799 -146 101975
rect -112 100799 -106 101975
rect -152 100787 -106 100799
rect 106 101975 152 101987
rect 106 100799 112 101975
rect 146 100799 152 101975
rect 106 100787 152 100799
rect -96 100749 96 100755
rect -96 100715 -84 100749
rect 84 100715 96 100749
rect -96 100709 96 100715
rect -96 100641 96 100647
rect -96 100607 -84 100641
rect 84 100607 96 100641
rect -96 100601 96 100607
rect -152 100557 -106 100569
rect -152 99381 -146 100557
rect -112 99381 -106 100557
rect -152 99369 -106 99381
rect 106 100557 152 100569
rect 106 99381 112 100557
rect 146 99381 152 100557
rect 106 99369 152 99381
rect -96 99331 96 99337
rect -96 99297 -84 99331
rect 84 99297 96 99331
rect -96 99291 96 99297
rect -96 99223 96 99229
rect -96 99189 -84 99223
rect 84 99189 96 99223
rect -96 99183 96 99189
rect -152 99139 -106 99151
rect -152 97963 -146 99139
rect -112 97963 -106 99139
rect -152 97951 -106 97963
rect 106 99139 152 99151
rect 106 97963 112 99139
rect 146 97963 152 99139
rect 106 97951 152 97963
rect -96 97913 96 97919
rect -96 97879 -84 97913
rect 84 97879 96 97913
rect -96 97873 96 97879
rect -96 97805 96 97811
rect -96 97771 -84 97805
rect 84 97771 96 97805
rect -96 97765 96 97771
rect -152 97721 -106 97733
rect -152 96545 -146 97721
rect -112 96545 -106 97721
rect -152 96533 -106 96545
rect 106 97721 152 97733
rect 106 96545 112 97721
rect 146 96545 152 97721
rect 106 96533 152 96545
rect -96 96495 96 96501
rect -96 96461 -84 96495
rect 84 96461 96 96495
rect -96 96455 96 96461
rect -96 96387 96 96393
rect -96 96353 -84 96387
rect 84 96353 96 96387
rect -96 96347 96 96353
rect -152 96303 -106 96315
rect -152 95127 -146 96303
rect -112 95127 -106 96303
rect -152 95115 -106 95127
rect 106 96303 152 96315
rect 106 95127 112 96303
rect 146 95127 152 96303
rect 106 95115 152 95127
rect -96 95077 96 95083
rect -96 95043 -84 95077
rect 84 95043 96 95077
rect -96 95037 96 95043
rect -96 94969 96 94975
rect -96 94935 -84 94969
rect 84 94935 96 94969
rect -96 94929 96 94935
rect -152 94885 -106 94897
rect -152 93709 -146 94885
rect -112 93709 -106 94885
rect -152 93697 -106 93709
rect 106 94885 152 94897
rect 106 93709 112 94885
rect 146 93709 152 94885
rect 106 93697 152 93709
rect -96 93659 96 93665
rect -96 93625 -84 93659
rect 84 93625 96 93659
rect -96 93619 96 93625
rect -96 93551 96 93557
rect -96 93517 -84 93551
rect 84 93517 96 93551
rect -96 93511 96 93517
rect -152 93467 -106 93479
rect -152 92291 -146 93467
rect -112 92291 -106 93467
rect -152 92279 -106 92291
rect 106 93467 152 93479
rect 106 92291 112 93467
rect 146 92291 152 93467
rect 106 92279 152 92291
rect -96 92241 96 92247
rect -96 92207 -84 92241
rect 84 92207 96 92241
rect -96 92201 96 92207
rect -96 92133 96 92139
rect -96 92099 -84 92133
rect 84 92099 96 92133
rect -96 92093 96 92099
rect -152 92049 -106 92061
rect -152 90873 -146 92049
rect -112 90873 -106 92049
rect -152 90861 -106 90873
rect 106 92049 152 92061
rect 106 90873 112 92049
rect 146 90873 152 92049
rect 106 90861 152 90873
rect -96 90823 96 90829
rect -96 90789 -84 90823
rect 84 90789 96 90823
rect -96 90783 96 90789
rect -96 90715 96 90721
rect -96 90681 -84 90715
rect 84 90681 96 90715
rect -96 90675 96 90681
rect -152 90631 -106 90643
rect -152 89455 -146 90631
rect -112 89455 -106 90631
rect -152 89443 -106 89455
rect 106 90631 152 90643
rect 106 89455 112 90631
rect 146 89455 152 90631
rect 106 89443 152 89455
rect -96 89405 96 89411
rect -96 89371 -84 89405
rect 84 89371 96 89405
rect -96 89365 96 89371
rect -96 89297 96 89303
rect -96 89263 -84 89297
rect 84 89263 96 89297
rect -96 89257 96 89263
rect -152 89213 -106 89225
rect -152 88037 -146 89213
rect -112 88037 -106 89213
rect -152 88025 -106 88037
rect 106 89213 152 89225
rect 106 88037 112 89213
rect 146 88037 152 89213
rect 106 88025 152 88037
rect -96 87987 96 87993
rect -96 87953 -84 87987
rect 84 87953 96 87987
rect -96 87947 96 87953
rect -96 87879 96 87885
rect -96 87845 -84 87879
rect 84 87845 96 87879
rect -96 87839 96 87845
rect -152 87795 -106 87807
rect -152 86619 -146 87795
rect -112 86619 -106 87795
rect -152 86607 -106 86619
rect 106 87795 152 87807
rect 106 86619 112 87795
rect 146 86619 152 87795
rect 106 86607 152 86619
rect -96 86569 96 86575
rect -96 86535 -84 86569
rect 84 86535 96 86569
rect -96 86529 96 86535
rect -96 86461 96 86467
rect -96 86427 -84 86461
rect 84 86427 96 86461
rect -96 86421 96 86427
rect -152 86377 -106 86389
rect -152 85201 -146 86377
rect -112 85201 -106 86377
rect -152 85189 -106 85201
rect 106 86377 152 86389
rect 106 85201 112 86377
rect 146 85201 152 86377
rect 106 85189 152 85201
rect -96 85151 96 85157
rect -96 85117 -84 85151
rect 84 85117 96 85151
rect -96 85111 96 85117
rect -96 85043 96 85049
rect -96 85009 -84 85043
rect 84 85009 96 85043
rect -96 85003 96 85009
rect -152 84959 -106 84971
rect -152 83783 -146 84959
rect -112 83783 -106 84959
rect -152 83771 -106 83783
rect 106 84959 152 84971
rect 106 83783 112 84959
rect 146 83783 152 84959
rect 106 83771 152 83783
rect -96 83733 96 83739
rect -96 83699 -84 83733
rect 84 83699 96 83733
rect -96 83693 96 83699
rect -96 83625 96 83631
rect -96 83591 -84 83625
rect 84 83591 96 83625
rect -96 83585 96 83591
rect -152 83541 -106 83553
rect -152 82365 -146 83541
rect -112 82365 -106 83541
rect -152 82353 -106 82365
rect 106 83541 152 83553
rect 106 82365 112 83541
rect 146 82365 152 83541
rect 106 82353 152 82365
rect -96 82315 96 82321
rect -96 82281 -84 82315
rect 84 82281 96 82315
rect -96 82275 96 82281
rect -96 82207 96 82213
rect -96 82173 -84 82207
rect 84 82173 96 82207
rect -96 82167 96 82173
rect -152 82123 -106 82135
rect -152 80947 -146 82123
rect -112 80947 -106 82123
rect -152 80935 -106 80947
rect 106 82123 152 82135
rect 106 80947 112 82123
rect 146 80947 152 82123
rect 106 80935 152 80947
rect -96 80897 96 80903
rect -96 80863 -84 80897
rect 84 80863 96 80897
rect -96 80857 96 80863
rect -96 80789 96 80795
rect -96 80755 -84 80789
rect 84 80755 96 80789
rect -96 80749 96 80755
rect -152 80705 -106 80717
rect -152 79529 -146 80705
rect -112 79529 -106 80705
rect -152 79517 -106 79529
rect 106 80705 152 80717
rect 106 79529 112 80705
rect 146 79529 152 80705
rect 106 79517 152 79529
rect -96 79479 96 79485
rect -96 79445 -84 79479
rect 84 79445 96 79479
rect -96 79439 96 79445
rect -96 79371 96 79377
rect -96 79337 -84 79371
rect 84 79337 96 79371
rect -96 79331 96 79337
rect -152 79287 -106 79299
rect -152 78111 -146 79287
rect -112 78111 -106 79287
rect -152 78099 -106 78111
rect 106 79287 152 79299
rect 106 78111 112 79287
rect 146 78111 152 79287
rect 106 78099 152 78111
rect -96 78061 96 78067
rect -96 78027 -84 78061
rect 84 78027 96 78061
rect -96 78021 96 78027
rect -96 77953 96 77959
rect -96 77919 -84 77953
rect 84 77919 96 77953
rect -96 77913 96 77919
rect -152 77869 -106 77881
rect -152 76693 -146 77869
rect -112 76693 -106 77869
rect -152 76681 -106 76693
rect 106 77869 152 77881
rect 106 76693 112 77869
rect 146 76693 152 77869
rect 106 76681 152 76693
rect -96 76643 96 76649
rect -96 76609 -84 76643
rect 84 76609 96 76643
rect -96 76603 96 76609
rect -96 76535 96 76541
rect -96 76501 -84 76535
rect 84 76501 96 76535
rect -96 76495 96 76501
rect -152 76451 -106 76463
rect -152 75275 -146 76451
rect -112 75275 -106 76451
rect -152 75263 -106 75275
rect 106 76451 152 76463
rect 106 75275 112 76451
rect 146 75275 152 76451
rect 106 75263 152 75275
rect -96 75225 96 75231
rect -96 75191 -84 75225
rect 84 75191 96 75225
rect -96 75185 96 75191
rect -96 75117 96 75123
rect -96 75083 -84 75117
rect 84 75083 96 75117
rect -96 75077 96 75083
rect -152 75033 -106 75045
rect -152 73857 -146 75033
rect -112 73857 -106 75033
rect -152 73845 -106 73857
rect 106 75033 152 75045
rect 106 73857 112 75033
rect 146 73857 152 75033
rect 106 73845 152 73857
rect -96 73807 96 73813
rect -96 73773 -84 73807
rect 84 73773 96 73807
rect -96 73767 96 73773
rect -96 73699 96 73705
rect -96 73665 -84 73699
rect 84 73665 96 73699
rect -96 73659 96 73665
rect -152 73615 -106 73627
rect -152 72439 -146 73615
rect -112 72439 -106 73615
rect -152 72427 -106 72439
rect 106 73615 152 73627
rect 106 72439 112 73615
rect 146 72439 152 73615
rect 106 72427 152 72439
rect -96 72389 96 72395
rect -96 72355 -84 72389
rect 84 72355 96 72389
rect -96 72349 96 72355
rect -96 72281 96 72287
rect -96 72247 -84 72281
rect 84 72247 96 72281
rect -96 72241 96 72247
rect -152 72197 -106 72209
rect -152 71021 -146 72197
rect -112 71021 -106 72197
rect -152 71009 -106 71021
rect 106 72197 152 72209
rect 106 71021 112 72197
rect 146 71021 152 72197
rect 106 71009 152 71021
rect -96 70971 96 70977
rect -96 70937 -84 70971
rect 84 70937 96 70971
rect -96 70931 96 70937
rect -96 70863 96 70869
rect -96 70829 -84 70863
rect 84 70829 96 70863
rect -96 70823 96 70829
rect -152 70779 -106 70791
rect -152 69603 -146 70779
rect -112 69603 -106 70779
rect -152 69591 -106 69603
rect 106 70779 152 70791
rect 106 69603 112 70779
rect 146 69603 152 70779
rect 106 69591 152 69603
rect -96 69553 96 69559
rect -96 69519 -84 69553
rect 84 69519 96 69553
rect -96 69513 96 69519
rect -96 69445 96 69451
rect -96 69411 -84 69445
rect 84 69411 96 69445
rect -96 69405 96 69411
rect -152 69361 -106 69373
rect -152 68185 -146 69361
rect -112 68185 -106 69361
rect -152 68173 -106 68185
rect 106 69361 152 69373
rect 106 68185 112 69361
rect 146 68185 152 69361
rect 106 68173 152 68185
rect -96 68135 96 68141
rect -96 68101 -84 68135
rect 84 68101 96 68135
rect -96 68095 96 68101
rect -96 68027 96 68033
rect -96 67993 -84 68027
rect 84 67993 96 68027
rect -96 67987 96 67993
rect -152 67943 -106 67955
rect -152 66767 -146 67943
rect -112 66767 -106 67943
rect -152 66755 -106 66767
rect 106 67943 152 67955
rect 106 66767 112 67943
rect 146 66767 152 67943
rect 106 66755 152 66767
rect -96 66717 96 66723
rect -96 66683 -84 66717
rect 84 66683 96 66717
rect -96 66677 96 66683
rect -96 66609 96 66615
rect -96 66575 -84 66609
rect 84 66575 96 66609
rect -96 66569 96 66575
rect -152 66525 -106 66537
rect -152 65349 -146 66525
rect -112 65349 -106 66525
rect -152 65337 -106 65349
rect 106 66525 152 66537
rect 106 65349 112 66525
rect 146 65349 152 66525
rect 106 65337 152 65349
rect -96 65299 96 65305
rect -96 65265 -84 65299
rect 84 65265 96 65299
rect -96 65259 96 65265
rect -96 65191 96 65197
rect -96 65157 -84 65191
rect 84 65157 96 65191
rect -96 65151 96 65157
rect -152 65107 -106 65119
rect -152 63931 -146 65107
rect -112 63931 -106 65107
rect -152 63919 -106 63931
rect 106 65107 152 65119
rect 106 63931 112 65107
rect 146 63931 152 65107
rect 106 63919 152 63931
rect -96 63881 96 63887
rect -96 63847 -84 63881
rect 84 63847 96 63881
rect -96 63841 96 63847
rect -96 63773 96 63779
rect -96 63739 -84 63773
rect 84 63739 96 63773
rect -96 63733 96 63739
rect -152 63689 -106 63701
rect -152 62513 -146 63689
rect -112 62513 -106 63689
rect -152 62501 -106 62513
rect 106 63689 152 63701
rect 106 62513 112 63689
rect 146 62513 152 63689
rect 106 62501 152 62513
rect -96 62463 96 62469
rect -96 62429 -84 62463
rect 84 62429 96 62463
rect -96 62423 96 62429
rect -96 62355 96 62361
rect -96 62321 -84 62355
rect 84 62321 96 62355
rect -96 62315 96 62321
rect -152 62271 -106 62283
rect -152 61095 -146 62271
rect -112 61095 -106 62271
rect -152 61083 -106 61095
rect 106 62271 152 62283
rect 106 61095 112 62271
rect 146 61095 152 62271
rect 106 61083 152 61095
rect -96 61045 96 61051
rect -96 61011 -84 61045
rect 84 61011 96 61045
rect -96 61005 96 61011
rect -96 60937 96 60943
rect -96 60903 -84 60937
rect 84 60903 96 60937
rect -96 60897 96 60903
rect -152 60853 -106 60865
rect -152 59677 -146 60853
rect -112 59677 -106 60853
rect -152 59665 -106 59677
rect 106 60853 152 60865
rect 106 59677 112 60853
rect 146 59677 152 60853
rect 106 59665 152 59677
rect -96 59627 96 59633
rect -96 59593 -84 59627
rect 84 59593 96 59627
rect -96 59587 96 59593
rect -96 59519 96 59525
rect -96 59485 -84 59519
rect 84 59485 96 59519
rect -96 59479 96 59485
rect -152 59435 -106 59447
rect -152 58259 -146 59435
rect -112 58259 -106 59435
rect -152 58247 -106 58259
rect 106 59435 152 59447
rect 106 58259 112 59435
rect 146 58259 152 59435
rect 106 58247 152 58259
rect -96 58209 96 58215
rect -96 58175 -84 58209
rect 84 58175 96 58209
rect -96 58169 96 58175
rect -96 58101 96 58107
rect -96 58067 -84 58101
rect 84 58067 96 58101
rect -96 58061 96 58067
rect -152 58017 -106 58029
rect -152 56841 -146 58017
rect -112 56841 -106 58017
rect -152 56829 -106 56841
rect 106 58017 152 58029
rect 106 56841 112 58017
rect 146 56841 152 58017
rect 106 56829 152 56841
rect -96 56791 96 56797
rect -96 56757 -84 56791
rect 84 56757 96 56791
rect -96 56751 96 56757
rect -96 56683 96 56689
rect -96 56649 -84 56683
rect 84 56649 96 56683
rect -96 56643 96 56649
rect -152 56599 -106 56611
rect -152 55423 -146 56599
rect -112 55423 -106 56599
rect -152 55411 -106 55423
rect 106 56599 152 56611
rect 106 55423 112 56599
rect 146 55423 152 56599
rect 106 55411 152 55423
rect -96 55373 96 55379
rect -96 55339 -84 55373
rect 84 55339 96 55373
rect -96 55333 96 55339
rect -96 55265 96 55271
rect -96 55231 -84 55265
rect 84 55231 96 55265
rect -96 55225 96 55231
rect -152 55181 -106 55193
rect -152 54005 -146 55181
rect -112 54005 -106 55181
rect -152 53993 -106 54005
rect 106 55181 152 55193
rect 106 54005 112 55181
rect 146 54005 152 55181
rect 106 53993 152 54005
rect -96 53955 96 53961
rect -96 53921 -84 53955
rect 84 53921 96 53955
rect -96 53915 96 53921
rect -96 53847 96 53853
rect -96 53813 -84 53847
rect 84 53813 96 53847
rect -96 53807 96 53813
rect -152 53763 -106 53775
rect -152 52587 -146 53763
rect -112 52587 -106 53763
rect -152 52575 -106 52587
rect 106 53763 152 53775
rect 106 52587 112 53763
rect 146 52587 152 53763
rect 106 52575 152 52587
rect -96 52537 96 52543
rect -96 52503 -84 52537
rect 84 52503 96 52537
rect -96 52497 96 52503
rect -96 52429 96 52435
rect -96 52395 -84 52429
rect 84 52395 96 52429
rect -96 52389 96 52395
rect -152 52345 -106 52357
rect -152 51169 -146 52345
rect -112 51169 -106 52345
rect -152 51157 -106 51169
rect 106 52345 152 52357
rect 106 51169 112 52345
rect 146 51169 152 52345
rect 106 51157 152 51169
rect -96 51119 96 51125
rect -96 51085 -84 51119
rect 84 51085 96 51119
rect -96 51079 96 51085
rect -96 51011 96 51017
rect -96 50977 -84 51011
rect 84 50977 96 51011
rect -96 50971 96 50977
rect -152 50927 -106 50939
rect -152 49751 -146 50927
rect -112 49751 -106 50927
rect -152 49739 -106 49751
rect 106 50927 152 50939
rect 106 49751 112 50927
rect 146 49751 152 50927
rect 106 49739 152 49751
rect -96 49701 96 49707
rect -96 49667 -84 49701
rect 84 49667 96 49701
rect -96 49661 96 49667
rect -96 49593 96 49599
rect -96 49559 -84 49593
rect 84 49559 96 49593
rect -96 49553 96 49559
rect -152 49509 -106 49521
rect -152 48333 -146 49509
rect -112 48333 -106 49509
rect -152 48321 -106 48333
rect 106 49509 152 49521
rect 106 48333 112 49509
rect 146 48333 152 49509
rect 106 48321 152 48333
rect -96 48283 96 48289
rect -96 48249 -84 48283
rect 84 48249 96 48283
rect -96 48243 96 48249
rect -96 48175 96 48181
rect -96 48141 -84 48175
rect 84 48141 96 48175
rect -96 48135 96 48141
rect -152 48091 -106 48103
rect -152 46915 -146 48091
rect -112 46915 -106 48091
rect -152 46903 -106 46915
rect 106 48091 152 48103
rect 106 46915 112 48091
rect 146 46915 152 48091
rect 106 46903 152 46915
rect -96 46865 96 46871
rect -96 46831 -84 46865
rect 84 46831 96 46865
rect -96 46825 96 46831
rect -96 46757 96 46763
rect -96 46723 -84 46757
rect 84 46723 96 46757
rect -96 46717 96 46723
rect -152 46673 -106 46685
rect -152 45497 -146 46673
rect -112 45497 -106 46673
rect -152 45485 -106 45497
rect 106 46673 152 46685
rect 106 45497 112 46673
rect 146 45497 152 46673
rect 106 45485 152 45497
rect -96 45447 96 45453
rect -96 45413 -84 45447
rect 84 45413 96 45447
rect -96 45407 96 45413
rect -96 45339 96 45345
rect -96 45305 -84 45339
rect 84 45305 96 45339
rect -96 45299 96 45305
rect -152 45255 -106 45267
rect -152 44079 -146 45255
rect -112 44079 -106 45255
rect -152 44067 -106 44079
rect 106 45255 152 45267
rect 106 44079 112 45255
rect 146 44079 152 45255
rect 106 44067 152 44079
rect -96 44029 96 44035
rect -96 43995 -84 44029
rect 84 43995 96 44029
rect -96 43989 96 43995
rect -96 43921 96 43927
rect -96 43887 -84 43921
rect 84 43887 96 43921
rect -96 43881 96 43887
rect -152 43837 -106 43849
rect -152 42661 -146 43837
rect -112 42661 -106 43837
rect -152 42649 -106 42661
rect 106 43837 152 43849
rect 106 42661 112 43837
rect 146 42661 152 43837
rect 106 42649 152 42661
rect -96 42611 96 42617
rect -96 42577 -84 42611
rect 84 42577 96 42611
rect -96 42571 96 42577
rect -96 42503 96 42509
rect -96 42469 -84 42503
rect 84 42469 96 42503
rect -96 42463 96 42469
rect -152 42419 -106 42431
rect -152 41243 -146 42419
rect -112 41243 -106 42419
rect -152 41231 -106 41243
rect 106 42419 152 42431
rect 106 41243 112 42419
rect 146 41243 152 42419
rect 106 41231 152 41243
rect -96 41193 96 41199
rect -96 41159 -84 41193
rect 84 41159 96 41193
rect -96 41153 96 41159
rect -96 41085 96 41091
rect -96 41051 -84 41085
rect 84 41051 96 41085
rect -96 41045 96 41051
rect -152 41001 -106 41013
rect -152 39825 -146 41001
rect -112 39825 -106 41001
rect -152 39813 -106 39825
rect 106 41001 152 41013
rect 106 39825 112 41001
rect 146 39825 152 41001
rect 106 39813 152 39825
rect -96 39775 96 39781
rect -96 39741 -84 39775
rect 84 39741 96 39775
rect -96 39735 96 39741
rect -96 39667 96 39673
rect -96 39633 -84 39667
rect 84 39633 96 39667
rect -96 39627 96 39633
rect -152 39583 -106 39595
rect -152 38407 -146 39583
rect -112 38407 -106 39583
rect -152 38395 -106 38407
rect 106 39583 152 39595
rect 106 38407 112 39583
rect 146 38407 152 39583
rect 106 38395 152 38407
rect -96 38357 96 38363
rect -96 38323 -84 38357
rect 84 38323 96 38357
rect -96 38317 96 38323
rect -96 38249 96 38255
rect -96 38215 -84 38249
rect 84 38215 96 38249
rect -96 38209 96 38215
rect -152 38165 -106 38177
rect -152 36989 -146 38165
rect -112 36989 -106 38165
rect -152 36977 -106 36989
rect 106 38165 152 38177
rect 106 36989 112 38165
rect 146 36989 152 38165
rect 106 36977 152 36989
rect -96 36939 96 36945
rect -96 36905 -84 36939
rect 84 36905 96 36939
rect -96 36899 96 36905
rect -96 36831 96 36837
rect -96 36797 -84 36831
rect 84 36797 96 36831
rect -96 36791 96 36797
rect -152 36747 -106 36759
rect -152 35571 -146 36747
rect -112 35571 -106 36747
rect -152 35559 -106 35571
rect 106 36747 152 36759
rect 106 35571 112 36747
rect 146 35571 152 36747
rect 106 35559 152 35571
rect -96 35521 96 35527
rect -96 35487 -84 35521
rect 84 35487 96 35521
rect -96 35481 96 35487
rect -96 35413 96 35419
rect -96 35379 -84 35413
rect 84 35379 96 35413
rect -96 35373 96 35379
rect -152 35329 -106 35341
rect -152 34153 -146 35329
rect -112 34153 -106 35329
rect -152 34141 -106 34153
rect 106 35329 152 35341
rect 106 34153 112 35329
rect 146 34153 152 35329
rect 106 34141 152 34153
rect -96 34103 96 34109
rect -96 34069 -84 34103
rect 84 34069 96 34103
rect -96 34063 96 34069
rect -96 33995 96 34001
rect -96 33961 -84 33995
rect 84 33961 96 33995
rect -96 33955 96 33961
rect -152 33911 -106 33923
rect -152 32735 -146 33911
rect -112 32735 -106 33911
rect -152 32723 -106 32735
rect 106 33911 152 33923
rect 106 32735 112 33911
rect 146 32735 152 33911
rect 106 32723 152 32735
rect -96 32685 96 32691
rect -96 32651 -84 32685
rect 84 32651 96 32685
rect -96 32645 96 32651
rect -96 32577 96 32583
rect -96 32543 -84 32577
rect 84 32543 96 32577
rect -96 32537 96 32543
rect -152 32493 -106 32505
rect -152 31317 -146 32493
rect -112 31317 -106 32493
rect -152 31305 -106 31317
rect 106 32493 152 32505
rect 106 31317 112 32493
rect 146 31317 152 32493
rect 106 31305 152 31317
rect -96 31267 96 31273
rect -96 31233 -84 31267
rect 84 31233 96 31267
rect -96 31227 96 31233
rect -96 31159 96 31165
rect -96 31125 -84 31159
rect 84 31125 96 31159
rect -96 31119 96 31125
rect -152 31075 -106 31087
rect -152 29899 -146 31075
rect -112 29899 -106 31075
rect -152 29887 -106 29899
rect 106 31075 152 31087
rect 106 29899 112 31075
rect 146 29899 152 31075
rect 106 29887 152 29899
rect -96 29849 96 29855
rect -96 29815 -84 29849
rect 84 29815 96 29849
rect -96 29809 96 29815
rect -96 29741 96 29747
rect -96 29707 -84 29741
rect 84 29707 96 29741
rect -96 29701 96 29707
rect -152 29657 -106 29669
rect -152 28481 -146 29657
rect -112 28481 -106 29657
rect -152 28469 -106 28481
rect 106 29657 152 29669
rect 106 28481 112 29657
rect 146 28481 152 29657
rect 106 28469 152 28481
rect -96 28431 96 28437
rect -96 28397 -84 28431
rect 84 28397 96 28431
rect -96 28391 96 28397
rect -96 28323 96 28329
rect -96 28289 -84 28323
rect 84 28289 96 28323
rect -96 28283 96 28289
rect -152 28239 -106 28251
rect -152 27063 -146 28239
rect -112 27063 -106 28239
rect -152 27051 -106 27063
rect 106 28239 152 28251
rect 106 27063 112 28239
rect 146 27063 152 28239
rect 106 27051 152 27063
rect -96 27013 96 27019
rect -96 26979 -84 27013
rect 84 26979 96 27013
rect -96 26973 96 26979
rect -96 26905 96 26911
rect -96 26871 -84 26905
rect 84 26871 96 26905
rect -96 26865 96 26871
rect -152 26821 -106 26833
rect -152 25645 -146 26821
rect -112 25645 -106 26821
rect -152 25633 -106 25645
rect 106 26821 152 26833
rect 106 25645 112 26821
rect 146 25645 152 26821
rect 106 25633 152 25645
rect -96 25595 96 25601
rect -96 25561 -84 25595
rect 84 25561 96 25595
rect -96 25555 96 25561
rect -96 25487 96 25493
rect -96 25453 -84 25487
rect 84 25453 96 25487
rect -96 25447 96 25453
rect -152 25403 -106 25415
rect -152 24227 -146 25403
rect -112 24227 -106 25403
rect -152 24215 -106 24227
rect 106 25403 152 25415
rect 106 24227 112 25403
rect 146 24227 152 25403
rect 106 24215 152 24227
rect -96 24177 96 24183
rect -96 24143 -84 24177
rect 84 24143 96 24177
rect -96 24137 96 24143
rect -96 24069 96 24075
rect -96 24035 -84 24069
rect 84 24035 96 24069
rect -96 24029 96 24035
rect -152 23985 -106 23997
rect -152 22809 -146 23985
rect -112 22809 -106 23985
rect -152 22797 -106 22809
rect 106 23985 152 23997
rect 106 22809 112 23985
rect 146 22809 152 23985
rect 106 22797 152 22809
rect -96 22759 96 22765
rect -96 22725 -84 22759
rect 84 22725 96 22759
rect -96 22719 96 22725
rect -96 22651 96 22657
rect -96 22617 -84 22651
rect 84 22617 96 22651
rect -96 22611 96 22617
rect -152 22567 -106 22579
rect -152 21391 -146 22567
rect -112 21391 -106 22567
rect -152 21379 -106 21391
rect 106 22567 152 22579
rect 106 21391 112 22567
rect 146 21391 152 22567
rect 106 21379 152 21391
rect -96 21341 96 21347
rect -96 21307 -84 21341
rect 84 21307 96 21341
rect -96 21301 96 21307
rect -96 21233 96 21239
rect -96 21199 -84 21233
rect 84 21199 96 21233
rect -96 21193 96 21199
rect -152 21149 -106 21161
rect -152 19973 -146 21149
rect -112 19973 -106 21149
rect -152 19961 -106 19973
rect 106 21149 152 21161
rect 106 19973 112 21149
rect 146 19973 152 21149
rect 106 19961 152 19973
rect -96 19923 96 19929
rect -96 19889 -84 19923
rect 84 19889 96 19923
rect -96 19883 96 19889
rect -96 19815 96 19821
rect -96 19781 -84 19815
rect 84 19781 96 19815
rect -96 19775 96 19781
rect -152 19731 -106 19743
rect -152 18555 -146 19731
rect -112 18555 -106 19731
rect -152 18543 -106 18555
rect 106 19731 152 19743
rect 106 18555 112 19731
rect 146 18555 152 19731
rect 106 18543 152 18555
rect -96 18505 96 18511
rect -96 18471 -84 18505
rect 84 18471 96 18505
rect -96 18465 96 18471
rect -96 18397 96 18403
rect -96 18363 -84 18397
rect 84 18363 96 18397
rect -96 18357 96 18363
rect -152 18313 -106 18325
rect -152 17137 -146 18313
rect -112 17137 -106 18313
rect -152 17125 -106 17137
rect 106 18313 152 18325
rect 106 17137 112 18313
rect 146 17137 152 18313
rect 106 17125 152 17137
rect -96 17087 96 17093
rect -96 17053 -84 17087
rect 84 17053 96 17087
rect -96 17047 96 17053
rect -96 16979 96 16985
rect -96 16945 -84 16979
rect 84 16945 96 16979
rect -96 16939 96 16945
rect -152 16895 -106 16907
rect -152 15719 -146 16895
rect -112 15719 -106 16895
rect -152 15707 -106 15719
rect 106 16895 152 16907
rect 106 15719 112 16895
rect 146 15719 152 16895
rect 106 15707 152 15719
rect -96 15669 96 15675
rect -96 15635 -84 15669
rect 84 15635 96 15669
rect -96 15629 96 15635
rect -96 15561 96 15567
rect -96 15527 -84 15561
rect 84 15527 96 15561
rect -96 15521 96 15527
rect -152 15477 -106 15489
rect -152 14301 -146 15477
rect -112 14301 -106 15477
rect -152 14289 -106 14301
rect 106 15477 152 15489
rect 106 14301 112 15477
rect 146 14301 152 15477
rect 106 14289 152 14301
rect -96 14251 96 14257
rect -96 14217 -84 14251
rect 84 14217 96 14251
rect -96 14211 96 14217
rect -96 14143 96 14149
rect -96 14109 -84 14143
rect 84 14109 96 14143
rect -96 14103 96 14109
rect -152 14059 -106 14071
rect -152 12883 -146 14059
rect -112 12883 -106 14059
rect -152 12871 -106 12883
rect 106 14059 152 14071
rect 106 12883 112 14059
rect 146 12883 152 14059
rect 106 12871 152 12883
rect -96 12833 96 12839
rect -96 12799 -84 12833
rect 84 12799 96 12833
rect -96 12793 96 12799
rect -96 12725 96 12731
rect -96 12691 -84 12725
rect 84 12691 96 12725
rect -96 12685 96 12691
rect -152 12641 -106 12653
rect -152 11465 -146 12641
rect -112 11465 -106 12641
rect -152 11453 -106 11465
rect 106 12641 152 12653
rect 106 11465 112 12641
rect 146 11465 152 12641
rect 106 11453 152 11465
rect -96 11415 96 11421
rect -96 11381 -84 11415
rect 84 11381 96 11415
rect -96 11375 96 11381
rect -96 11307 96 11313
rect -96 11273 -84 11307
rect 84 11273 96 11307
rect -96 11267 96 11273
rect -152 11223 -106 11235
rect -152 10047 -146 11223
rect -112 10047 -106 11223
rect -152 10035 -106 10047
rect 106 11223 152 11235
rect 106 10047 112 11223
rect 146 10047 152 11223
rect 106 10035 152 10047
rect -96 9997 96 10003
rect -96 9963 -84 9997
rect 84 9963 96 9997
rect -96 9957 96 9963
rect -96 9889 96 9895
rect -96 9855 -84 9889
rect 84 9855 96 9889
rect -96 9849 96 9855
rect -152 9805 -106 9817
rect -152 8629 -146 9805
rect -112 8629 -106 9805
rect -152 8617 -106 8629
rect 106 9805 152 9817
rect 106 8629 112 9805
rect 146 8629 152 9805
rect 106 8617 152 8629
rect -96 8579 96 8585
rect -96 8545 -84 8579
rect 84 8545 96 8579
rect -96 8539 96 8545
rect -96 8471 96 8477
rect -96 8437 -84 8471
rect 84 8437 96 8471
rect -96 8431 96 8437
rect -152 8387 -106 8399
rect -152 7211 -146 8387
rect -112 7211 -106 8387
rect -152 7199 -106 7211
rect 106 8387 152 8399
rect 106 7211 112 8387
rect 146 7211 152 8387
rect 106 7199 152 7211
rect -96 7161 96 7167
rect -96 7127 -84 7161
rect 84 7127 96 7161
rect -96 7121 96 7127
rect -96 7053 96 7059
rect -96 7019 -84 7053
rect 84 7019 96 7053
rect -96 7013 96 7019
rect -152 6969 -106 6981
rect -152 5793 -146 6969
rect -112 5793 -106 6969
rect -152 5781 -106 5793
rect 106 6969 152 6981
rect 106 5793 112 6969
rect 146 5793 152 6969
rect 106 5781 152 5793
rect -96 5743 96 5749
rect -96 5709 -84 5743
rect 84 5709 96 5743
rect -96 5703 96 5709
rect -96 5635 96 5641
rect -96 5601 -84 5635
rect 84 5601 96 5635
rect -96 5595 96 5601
rect -152 5551 -106 5563
rect -152 4375 -146 5551
rect -112 4375 -106 5551
rect -152 4363 -106 4375
rect 106 5551 152 5563
rect 106 4375 112 5551
rect 146 4375 152 5551
rect 106 4363 152 4375
rect -96 4325 96 4331
rect -96 4291 -84 4325
rect 84 4291 96 4325
rect -96 4285 96 4291
rect -96 4217 96 4223
rect -96 4183 -84 4217
rect 84 4183 96 4217
rect -96 4177 96 4183
rect -152 4133 -106 4145
rect -152 2957 -146 4133
rect -112 2957 -106 4133
rect -152 2945 -106 2957
rect 106 4133 152 4145
rect 106 2957 112 4133
rect 146 2957 152 4133
rect 106 2945 152 2957
rect -96 2907 96 2913
rect -96 2873 -84 2907
rect 84 2873 96 2907
rect -96 2867 96 2873
rect -96 2799 96 2805
rect -96 2765 -84 2799
rect 84 2765 96 2799
rect -96 2759 96 2765
rect -152 2715 -106 2727
rect -152 1539 -146 2715
rect -112 1539 -106 2715
rect -152 1527 -106 1539
rect 106 2715 152 2727
rect 106 1539 112 2715
rect 146 1539 152 2715
rect 106 1527 152 1539
rect -96 1489 96 1495
rect -96 1455 -84 1489
rect 84 1455 96 1489
rect -96 1449 96 1455
rect -96 1381 96 1387
rect -96 1347 -84 1381
rect 84 1347 96 1381
rect -96 1341 96 1347
rect -152 1297 -106 1309
rect -152 121 -146 1297
rect -112 121 -106 1297
rect -152 109 -106 121
rect 106 1297 152 1309
rect 106 121 112 1297
rect 146 121 152 1297
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -1297 -146 -121
rect -112 -1297 -106 -121
rect -152 -1309 -106 -1297
rect 106 -121 152 -109
rect 106 -1297 112 -121
rect 146 -1297 152 -121
rect 106 -1309 152 -1297
rect -96 -1347 96 -1341
rect -96 -1381 -84 -1347
rect 84 -1381 96 -1347
rect -96 -1387 96 -1381
rect -96 -1455 96 -1449
rect -96 -1489 -84 -1455
rect 84 -1489 96 -1455
rect -96 -1495 96 -1489
rect -152 -1539 -106 -1527
rect -152 -2715 -146 -1539
rect -112 -2715 -106 -1539
rect -152 -2727 -106 -2715
rect 106 -1539 152 -1527
rect 106 -2715 112 -1539
rect 146 -2715 152 -1539
rect 106 -2727 152 -2715
rect -96 -2765 96 -2759
rect -96 -2799 -84 -2765
rect 84 -2799 96 -2765
rect -96 -2805 96 -2799
rect -96 -2873 96 -2867
rect -96 -2907 -84 -2873
rect 84 -2907 96 -2873
rect -96 -2913 96 -2907
rect -152 -2957 -106 -2945
rect -152 -4133 -146 -2957
rect -112 -4133 -106 -2957
rect -152 -4145 -106 -4133
rect 106 -2957 152 -2945
rect 106 -4133 112 -2957
rect 146 -4133 152 -2957
rect 106 -4145 152 -4133
rect -96 -4183 96 -4177
rect -96 -4217 -84 -4183
rect 84 -4217 96 -4183
rect -96 -4223 96 -4217
rect -96 -4291 96 -4285
rect -96 -4325 -84 -4291
rect 84 -4325 96 -4291
rect -96 -4331 96 -4325
rect -152 -4375 -106 -4363
rect -152 -5551 -146 -4375
rect -112 -5551 -106 -4375
rect -152 -5563 -106 -5551
rect 106 -4375 152 -4363
rect 106 -5551 112 -4375
rect 146 -5551 152 -4375
rect 106 -5563 152 -5551
rect -96 -5601 96 -5595
rect -96 -5635 -84 -5601
rect 84 -5635 96 -5601
rect -96 -5641 96 -5635
rect -96 -5709 96 -5703
rect -96 -5743 -84 -5709
rect 84 -5743 96 -5709
rect -96 -5749 96 -5743
rect -152 -5793 -106 -5781
rect -152 -6969 -146 -5793
rect -112 -6969 -106 -5793
rect -152 -6981 -106 -6969
rect 106 -5793 152 -5781
rect 106 -6969 112 -5793
rect 146 -6969 152 -5793
rect 106 -6981 152 -6969
rect -96 -7019 96 -7013
rect -96 -7053 -84 -7019
rect 84 -7053 96 -7019
rect -96 -7059 96 -7053
rect -96 -7127 96 -7121
rect -96 -7161 -84 -7127
rect 84 -7161 96 -7127
rect -96 -7167 96 -7161
rect -152 -7211 -106 -7199
rect -152 -8387 -146 -7211
rect -112 -8387 -106 -7211
rect -152 -8399 -106 -8387
rect 106 -7211 152 -7199
rect 106 -8387 112 -7211
rect 146 -8387 152 -7211
rect 106 -8399 152 -8387
rect -96 -8437 96 -8431
rect -96 -8471 -84 -8437
rect 84 -8471 96 -8437
rect -96 -8477 96 -8471
rect -96 -8545 96 -8539
rect -96 -8579 -84 -8545
rect 84 -8579 96 -8545
rect -96 -8585 96 -8579
rect -152 -8629 -106 -8617
rect -152 -9805 -146 -8629
rect -112 -9805 -106 -8629
rect -152 -9817 -106 -9805
rect 106 -8629 152 -8617
rect 106 -9805 112 -8629
rect 146 -9805 152 -8629
rect 106 -9817 152 -9805
rect -96 -9855 96 -9849
rect -96 -9889 -84 -9855
rect 84 -9889 96 -9855
rect -96 -9895 96 -9889
rect -96 -9963 96 -9957
rect -96 -9997 -84 -9963
rect 84 -9997 96 -9963
rect -96 -10003 96 -9997
rect -152 -10047 -106 -10035
rect -152 -11223 -146 -10047
rect -112 -11223 -106 -10047
rect -152 -11235 -106 -11223
rect 106 -10047 152 -10035
rect 106 -11223 112 -10047
rect 146 -11223 152 -10047
rect 106 -11235 152 -11223
rect -96 -11273 96 -11267
rect -96 -11307 -84 -11273
rect 84 -11307 96 -11273
rect -96 -11313 96 -11307
rect -96 -11381 96 -11375
rect -96 -11415 -84 -11381
rect 84 -11415 96 -11381
rect -96 -11421 96 -11415
rect -152 -11465 -106 -11453
rect -152 -12641 -146 -11465
rect -112 -12641 -106 -11465
rect -152 -12653 -106 -12641
rect 106 -11465 152 -11453
rect 106 -12641 112 -11465
rect 146 -12641 152 -11465
rect 106 -12653 152 -12641
rect -96 -12691 96 -12685
rect -96 -12725 -84 -12691
rect 84 -12725 96 -12691
rect -96 -12731 96 -12725
rect -96 -12799 96 -12793
rect -96 -12833 -84 -12799
rect 84 -12833 96 -12799
rect -96 -12839 96 -12833
rect -152 -12883 -106 -12871
rect -152 -14059 -146 -12883
rect -112 -14059 -106 -12883
rect -152 -14071 -106 -14059
rect 106 -12883 152 -12871
rect 106 -14059 112 -12883
rect 146 -14059 152 -12883
rect 106 -14071 152 -14059
rect -96 -14109 96 -14103
rect -96 -14143 -84 -14109
rect 84 -14143 96 -14109
rect -96 -14149 96 -14143
rect -96 -14217 96 -14211
rect -96 -14251 -84 -14217
rect 84 -14251 96 -14217
rect -96 -14257 96 -14251
rect -152 -14301 -106 -14289
rect -152 -15477 -146 -14301
rect -112 -15477 -106 -14301
rect -152 -15489 -106 -15477
rect 106 -14301 152 -14289
rect 106 -15477 112 -14301
rect 146 -15477 152 -14301
rect 106 -15489 152 -15477
rect -96 -15527 96 -15521
rect -96 -15561 -84 -15527
rect 84 -15561 96 -15527
rect -96 -15567 96 -15561
rect -96 -15635 96 -15629
rect -96 -15669 -84 -15635
rect 84 -15669 96 -15635
rect -96 -15675 96 -15669
rect -152 -15719 -106 -15707
rect -152 -16895 -146 -15719
rect -112 -16895 -106 -15719
rect -152 -16907 -106 -16895
rect 106 -15719 152 -15707
rect 106 -16895 112 -15719
rect 146 -16895 152 -15719
rect 106 -16907 152 -16895
rect -96 -16945 96 -16939
rect -96 -16979 -84 -16945
rect 84 -16979 96 -16945
rect -96 -16985 96 -16979
rect -96 -17053 96 -17047
rect -96 -17087 -84 -17053
rect 84 -17087 96 -17053
rect -96 -17093 96 -17087
rect -152 -17137 -106 -17125
rect -152 -18313 -146 -17137
rect -112 -18313 -106 -17137
rect -152 -18325 -106 -18313
rect 106 -17137 152 -17125
rect 106 -18313 112 -17137
rect 146 -18313 152 -17137
rect 106 -18325 152 -18313
rect -96 -18363 96 -18357
rect -96 -18397 -84 -18363
rect 84 -18397 96 -18363
rect -96 -18403 96 -18397
rect -96 -18471 96 -18465
rect -96 -18505 -84 -18471
rect 84 -18505 96 -18471
rect -96 -18511 96 -18505
rect -152 -18555 -106 -18543
rect -152 -19731 -146 -18555
rect -112 -19731 -106 -18555
rect -152 -19743 -106 -19731
rect 106 -18555 152 -18543
rect 106 -19731 112 -18555
rect 146 -19731 152 -18555
rect 106 -19743 152 -19731
rect -96 -19781 96 -19775
rect -96 -19815 -84 -19781
rect 84 -19815 96 -19781
rect -96 -19821 96 -19815
rect -96 -19889 96 -19883
rect -96 -19923 -84 -19889
rect 84 -19923 96 -19889
rect -96 -19929 96 -19923
rect -152 -19973 -106 -19961
rect -152 -21149 -146 -19973
rect -112 -21149 -106 -19973
rect -152 -21161 -106 -21149
rect 106 -19973 152 -19961
rect 106 -21149 112 -19973
rect 146 -21149 152 -19973
rect 106 -21161 152 -21149
rect -96 -21199 96 -21193
rect -96 -21233 -84 -21199
rect 84 -21233 96 -21199
rect -96 -21239 96 -21233
rect -96 -21307 96 -21301
rect -96 -21341 -84 -21307
rect 84 -21341 96 -21307
rect -96 -21347 96 -21341
rect -152 -21391 -106 -21379
rect -152 -22567 -146 -21391
rect -112 -22567 -106 -21391
rect -152 -22579 -106 -22567
rect 106 -21391 152 -21379
rect 106 -22567 112 -21391
rect 146 -22567 152 -21391
rect 106 -22579 152 -22567
rect -96 -22617 96 -22611
rect -96 -22651 -84 -22617
rect 84 -22651 96 -22617
rect -96 -22657 96 -22651
rect -96 -22725 96 -22719
rect -96 -22759 -84 -22725
rect 84 -22759 96 -22725
rect -96 -22765 96 -22759
rect -152 -22809 -106 -22797
rect -152 -23985 -146 -22809
rect -112 -23985 -106 -22809
rect -152 -23997 -106 -23985
rect 106 -22809 152 -22797
rect 106 -23985 112 -22809
rect 146 -23985 152 -22809
rect 106 -23997 152 -23985
rect -96 -24035 96 -24029
rect -96 -24069 -84 -24035
rect 84 -24069 96 -24035
rect -96 -24075 96 -24069
rect -96 -24143 96 -24137
rect -96 -24177 -84 -24143
rect 84 -24177 96 -24143
rect -96 -24183 96 -24177
rect -152 -24227 -106 -24215
rect -152 -25403 -146 -24227
rect -112 -25403 -106 -24227
rect -152 -25415 -106 -25403
rect 106 -24227 152 -24215
rect 106 -25403 112 -24227
rect 146 -25403 152 -24227
rect 106 -25415 152 -25403
rect -96 -25453 96 -25447
rect -96 -25487 -84 -25453
rect 84 -25487 96 -25453
rect -96 -25493 96 -25487
rect -96 -25561 96 -25555
rect -96 -25595 -84 -25561
rect 84 -25595 96 -25561
rect -96 -25601 96 -25595
rect -152 -25645 -106 -25633
rect -152 -26821 -146 -25645
rect -112 -26821 -106 -25645
rect -152 -26833 -106 -26821
rect 106 -25645 152 -25633
rect 106 -26821 112 -25645
rect 146 -26821 152 -25645
rect 106 -26833 152 -26821
rect -96 -26871 96 -26865
rect -96 -26905 -84 -26871
rect 84 -26905 96 -26871
rect -96 -26911 96 -26905
rect -96 -26979 96 -26973
rect -96 -27013 -84 -26979
rect 84 -27013 96 -26979
rect -96 -27019 96 -27013
rect -152 -27063 -106 -27051
rect -152 -28239 -146 -27063
rect -112 -28239 -106 -27063
rect -152 -28251 -106 -28239
rect 106 -27063 152 -27051
rect 106 -28239 112 -27063
rect 146 -28239 152 -27063
rect 106 -28251 152 -28239
rect -96 -28289 96 -28283
rect -96 -28323 -84 -28289
rect 84 -28323 96 -28289
rect -96 -28329 96 -28323
rect -96 -28397 96 -28391
rect -96 -28431 -84 -28397
rect 84 -28431 96 -28397
rect -96 -28437 96 -28431
rect -152 -28481 -106 -28469
rect -152 -29657 -146 -28481
rect -112 -29657 -106 -28481
rect -152 -29669 -106 -29657
rect 106 -28481 152 -28469
rect 106 -29657 112 -28481
rect 146 -29657 152 -28481
rect 106 -29669 152 -29657
rect -96 -29707 96 -29701
rect -96 -29741 -84 -29707
rect 84 -29741 96 -29707
rect -96 -29747 96 -29741
rect -96 -29815 96 -29809
rect -96 -29849 -84 -29815
rect 84 -29849 96 -29815
rect -96 -29855 96 -29849
rect -152 -29899 -106 -29887
rect -152 -31075 -146 -29899
rect -112 -31075 -106 -29899
rect -152 -31087 -106 -31075
rect 106 -29899 152 -29887
rect 106 -31075 112 -29899
rect 146 -31075 152 -29899
rect 106 -31087 152 -31075
rect -96 -31125 96 -31119
rect -96 -31159 -84 -31125
rect 84 -31159 96 -31125
rect -96 -31165 96 -31159
rect -96 -31233 96 -31227
rect -96 -31267 -84 -31233
rect 84 -31267 96 -31233
rect -96 -31273 96 -31267
rect -152 -31317 -106 -31305
rect -152 -32493 -146 -31317
rect -112 -32493 -106 -31317
rect -152 -32505 -106 -32493
rect 106 -31317 152 -31305
rect 106 -32493 112 -31317
rect 146 -32493 152 -31317
rect 106 -32505 152 -32493
rect -96 -32543 96 -32537
rect -96 -32577 -84 -32543
rect 84 -32577 96 -32543
rect -96 -32583 96 -32577
rect -96 -32651 96 -32645
rect -96 -32685 -84 -32651
rect 84 -32685 96 -32651
rect -96 -32691 96 -32685
rect -152 -32735 -106 -32723
rect -152 -33911 -146 -32735
rect -112 -33911 -106 -32735
rect -152 -33923 -106 -33911
rect 106 -32735 152 -32723
rect 106 -33911 112 -32735
rect 146 -33911 152 -32735
rect 106 -33923 152 -33911
rect -96 -33961 96 -33955
rect -96 -33995 -84 -33961
rect 84 -33995 96 -33961
rect -96 -34001 96 -33995
rect -96 -34069 96 -34063
rect -96 -34103 -84 -34069
rect 84 -34103 96 -34069
rect -96 -34109 96 -34103
rect -152 -34153 -106 -34141
rect -152 -35329 -146 -34153
rect -112 -35329 -106 -34153
rect -152 -35341 -106 -35329
rect 106 -34153 152 -34141
rect 106 -35329 112 -34153
rect 146 -35329 152 -34153
rect 106 -35341 152 -35329
rect -96 -35379 96 -35373
rect -96 -35413 -84 -35379
rect 84 -35413 96 -35379
rect -96 -35419 96 -35413
rect -96 -35487 96 -35481
rect -96 -35521 -84 -35487
rect 84 -35521 96 -35487
rect -96 -35527 96 -35521
rect -152 -35571 -106 -35559
rect -152 -36747 -146 -35571
rect -112 -36747 -106 -35571
rect -152 -36759 -106 -36747
rect 106 -35571 152 -35559
rect 106 -36747 112 -35571
rect 146 -36747 152 -35571
rect 106 -36759 152 -36747
rect -96 -36797 96 -36791
rect -96 -36831 -84 -36797
rect 84 -36831 96 -36797
rect -96 -36837 96 -36831
rect -96 -36905 96 -36899
rect -96 -36939 -84 -36905
rect 84 -36939 96 -36905
rect -96 -36945 96 -36939
rect -152 -36989 -106 -36977
rect -152 -38165 -146 -36989
rect -112 -38165 -106 -36989
rect -152 -38177 -106 -38165
rect 106 -36989 152 -36977
rect 106 -38165 112 -36989
rect 146 -38165 152 -36989
rect 106 -38177 152 -38165
rect -96 -38215 96 -38209
rect -96 -38249 -84 -38215
rect 84 -38249 96 -38215
rect -96 -38255 96 -38249
rect -96 -38323 96 -38317
rect -96 -38357 -84 -38323
rect 84 -38357 96 -38323
rect -96 -38363 96 -38357
rect -152 -38407 -106 -38395
rect -152 -39583 -146 -38407
rect -112 -39583 -106 -38407
rect -152 -39595 -106 -39583
rect 106 -38407 152 -38395
rect 106 -39583 112 -38407
rect 146 -39583 152 -38407
rect 106 -39595 152 -39583
rect -96 -39633 96 -39627
rect -96 -39667 -84 -39633
rect 84 -39667 96 -39633
rect -96 -39673 96 -39667
rect -96 -39741 96 -39735
rect -96 -39775 -84 -39741
rect 84 -39775 96 -39741
rect -96 -39781 96 -39775
rect -152 -39825 -106 -39813
rect -152 -41001 -146 -39825
rect -112 -41001 -106 -39825
rect -152 -41013 -106 -41001
rect 106 -39825 152 -39813
rect 106 -41001 112 -39825
rect 146 -41001 152 -39825
rect 106 -41013 152 -41001
rect -96 -41051 96 -41045
rect -96 -41085 -84 -41051
rect 84 -41085 96 -41051
rect -96 -41091 96 -41085
rect -96 -41159 96 -41153
rect -96 -41193 -84 -41159
rect 84 -41193 96 -41159
rect -96 -41199 96 -41193
rect -152 -41243 -106 -41231
rect -152 -42419 -146 -41243
rect -112 -42419 -106 -41243
rect -152 -42431 -106 -42419
rect 106 -41243 152 -41231
rect 106 -42419 112 -41243
rect 146 -42419 152 -41243
rect 106 -42431 152 -42419
rect -96 -42469 96 -42463
rect -96 -42503 -84 -42469
rect 84 -42503 96 -42469
rect -96 -42509 96 -42503
rect -96 -42577 96 -42571
rect -96 -42611 -84 -42577
rect 84 -42611 96 -42577
rect -96 -42617 96 -42611
rect -152 -42661 -106 -42649
rect -152 -43837 -146 -42661
rect -112 -43837 -106 -42661
rect -152 -43849 -106 -43837
rect 106 -42661 152 -42649
rect 106 -43837 112 -42661
rect 146 -43837 152 -42661
rect 106 -43849 152 -43837
rect -96 -43887 96 -43881
rect -96 -43921 -84 -43887
rect 84 -43921 96 -43887
rect -96 -43927 96 -43921
rect -96 -43995 96 -43989
rect -96 -44029 -84 -43995
rect 84 -44029 96 -43995
rect -96 -44035 96 -44029
rect -152 -44079 -106 -44067
rect -152 -45255 -146 -44079
rect -112 -45255 -106 -44079
rect -152 -45267 -106 -45255
rect 106 -44079 152 -44067
rect 106 -45255 112 -44079
rect 146 -45255 152 -44079
rect 106 -45267 152 -45255
rect -96 -45305 96 -45299
rect -96 -45339 -84 -45305
rect 84 -45339 96 -45305
rect -96 -45345 96 -45339
rect -96 -45413 96 -45407
rect -96 -45447 -84 -45413
rect 84 -45447 96 -45413
rect -96 -45453 96 -45447
rect -152 -45497 -106 -45485
rect -152 -46673 -146 -45497
rect -112 -46673 -106 -45497
rect -152 -46685 -106 -46673
rect 106 -45497 152 -45485
rect 106 -46673 112 -45497
rect 146 -46673 152 -45497
rect 106 -46685 152 -46673
rect -96 -46723 96 -46717
rect -96 -46757 -84 -46723
rect 84 -46757 96 -46723
rect -96 -46763 96 -46757
rect -96 -46831 96 -46825
rect -96 -46865 -84 -46831
rect 84 -46865 96 -46831
rect -96 -46871 96 -46865
rect -152 -46915 -106 -46903
rect -152 -48091 -146 -46915
rect -112 -48091 -106 -46915
rect -152 -48103 -106 -48091
rect 106 -46915 152 -46903
rect 106 -48091 112 -46915
rect 146 -48091 152 -46915
rect 106 -48103 152 -48091
rect -96 -48141 96 -48135
rect -96 -48175 -84 -48141
rect 84 -48175 96 -48141
rect -96 -48181 96 -48175
rect -96 -48249 96 -48243
rect -96 -48283 -84 -48249
rect 84 -48283 96 -48249
rect -96 -48289 96 -48283
rect -152 -48333 -106 -48321
rect -152 -49509 -146 -48333
rect -112 -49509 -106 -48333
rect -152 -49521 -106 -49509
rect 106 -48333 152 -48321
rect 106 -49509 112 -48333
rect 146 -49509 152 -48333
rect 106 -49521 152 -49509
rect -96 -49559 96 -49553
rect -96 -49593 -84 -49559
rect 84 -49593 96 -49559
rect -96 -49599 96 -49593
rect -96 -49667 96 -49661
rect -96 -49701 -84 -49667
rect 84 -49701 96 -49667
rect -96 -49707 96 -49701
rect -152 -49751 -106 -49739
rect -152 -50927 -146 -49751
rect -112 -50927 -106 -49751
rect -152 -50939 -106 -50927
rect 106 -49751 152 -49739
rect 106 -50927 112 -49751
rect 146 -50927 152 -49751
rect 106 -50939 152 -50927
rect -96 -50977 96 -50971
rect -96 -51011 -84 -50977
rect 84 -51011 96 -50977
rect -96 -51017 96 -51011
rect -96 -51085 96 -51079
rect -96 -51119 -84 -51085
rect 84 -51119 96 -51085
rect -96 -51125 96 -51119
rect -152 -51169 -106 -51157
rect -152 -52345 -146 -51169
rect -112 -52345 -106 -51169
rect -152 -52357 -106 -52345
rect 106 -51169 152 -51157
rect 106 -52345 112 -51169
rect 146 -52345 152 -51169
rect 106 -52357 152 -52345
rect -96 -52395 96 -52389
rect -96 -52429 -84 -52395
rect 84 -52429 96 -52395
rect -96 -52435 96 -52429
rect -96 -52503 96 -52497
rect -96 -52537 -84 -52503
rect 84 -52537 96 -52503
rect -96 -52543 96 -52537
rect -152 -52587 -106 -52575
rect -152 -53763 -146 -52587
rect -112 -53763 -106 -52587
rect -152 -53775 -106 -53763
rect 106 -52587 152 -52575
rect 106 -53763 112 -52587
rect 146 -53763 152 -52587
rect 106 -53775 152 -53763
rect -96 -53813 96 -53807
rect -96 -53847 -84 -53813
rect 84 -53847 96 -53813
rect -96 -53853 96 -53847
rect -96 -53921 96 -53915
rect -96 -53955 -84 -53921
rect 84 -53955 96 -53921
rect -96 -53961 96 -53955
rect -152 -54005 -106 -53993
rect -152 -55181 -146 -54005
rect -112 -55181 -106 -54005
rect -152 -55193 -106 -55181
rect 106 -54005 152 -53993
rect 106 -55181 112 -54005
rect 146 -55181 152 -54005
rect 106 -55193 152 -55181
rect -96 -55231 96 -55225
rect -96 -55265 -84 -55231
rect 84 -55265 96 -55231
rect -96 -55271 96 -55265
rect -96 -55339 96 -55333
rect -96 -55373 -84 -55339
rect 84 -55373 96 -55339
rect -96 -55379 96 -55373
rect -152 -55423 -106 -55411
rect -152 -56599 -146 -55423
rect -112 -56599 -106 -55423
rect -152 -56611 -106 -56599
rect 106 -55423 152 -55411
rect 106 -56599 112 -55423
rect 146 -56599 152 -55423
rect 106 -56611 152 -56599
rect -96 -56649 96 -56643
rect -96 -56683 -84 -56649
rect 84 -56683 96 -56649
rect -96 -56689 96 -56683
rect -96 -56757 96 -56751
rect -96 -56791 -84 -56757
rect 84 -56791 96 -56757
rect -96 -56797 96 -56791
rect -152 -56841 -106 -56829
rect -152 -58017 -146 -56841
rect -112 -58017 -106 -56841
rect -152 -58029 -106 -58017
rect 106 -56841 152 -56829
rect 106 -58017 112 -56841
rect 146 -58017 152 -56841
rect 106 -58029 152 -58017
rect -96 -58067 96 -58061
rect -96 -58101 -84 -58067
rect 84 -58101 96 -58067
rect -96 -58107 96 -58101
rect -96 -58175 96 -58169
rect -96 -58209 -84 -58175
rect 84 -58209 96 -58175
rect -96 -58215 96 -58209
rect -152 -58259 -106 -58247
rect -152 -59435 -146 -58259
rect -112 -59435 -106 -58259
rect -152 -59447 -106 -59435
rect 106 -58259 152 -58247
rect 106 -59435 112 -58259
rect 146 -59435 152 -58259
rect 106 -59447 152 -59435
rect -96 -59485 96 -59479
rect -96 -59519 -84 -59485
rect 84 -59519 96 -59485
rect -96 -59525 96 -59519
rect -96 -59593 96 -59587
rect -96 -59627 -84 -59593
rect 84 -59627 96 -59593
rect -96 -59633 96 -59627
rect -152 -59677 -106 -59665
rect -152 -60853 -146 -59677
rect -112 -60853 -106 -59677
rect -152 -60865 -106 -60853
rect 106 -59677 152 -59665
rect 106 -60853 112 -59677
rect 146 -60853 152 -59677
rect 106 -60865 152 -60853
rect -96 -60903 96 -60897
rect -96 -60937 -84 -60903
rect 84 -60937 96 -60903
rect -96 -60943 96 -60937
rect -96 -61011 96 -61005
rect -96 -61045 -84 -61011
rect 84 -61045 96 -61011
rect -96 -61051 96 -61045
rect -152 -61095 -106 -61083
rect -152 -62271 -146 -61095
rect -112 -62271 -106 -61095
rect -152 -62283 -106 -62271
rect 106 -61095 152 -61083
rect 106 -62271 112 -61095
rect 146 -62271 152 -61095
rect 106 -62283 152 -62271
rect -96 -62321 96 -62315
rect -96 -62355 -84 -62321
rect 84 -62355 96 -62321
rect -96 -62361 96 -62355
rect -96 -62429 96 -62423
rect -96 -62463 -84 -62429
rect 84 -62463 96 -62429
rect -96 -62469 96 -62463
rect -152 -62513 -106 -62501
rect -152 -63689 -146 -62513
rect -112 -63689 -106 -62513
rect -152 -63701 -106 -63689
rect 106 -62513 152 -62501
rect 106 -63689 112 -62513
rect 146 -63689 152 -62513
rect 106 -63701 152 -63689
rect -96 -63739 96 -63733
rect -96 -63773 -84 -63739
rect 84 -63773 96 -63739
rect -96 -63779 96 -63773
rect -96 -63847 96 -63841
rect -96 -63881 -84 -63847
rect 84 -63881 96 -63847
rect -96 -63887 96 -63881
rect -152 -63931 -106 -63919
rect -152 -65107 -146 -63931
rect -112 -65107 -106 -63931
rect -152 -65119 -106 -65107
rect 106 -63931 152 -63919
rect 106 -65107 112 -63931
rect 146 -65107 152 -63931
rect 106 -65119 152 -65107
rect -96 -65157 96 -65151
rect -96 -65191 -84 -65157
rect 84 -65191 96 -65157
rect -96 -65197 96 -65191
rect -96 -65265 96 -65259
rect -96 -65299 -84 -65265
rect 84 -65299 96 -65265
rect -96 -65305 96 -65299
rect -152 -65349 -106 -65337
rect -152 -66525 -146 -65349
rect -112 -66525 -106 -65349
rect -152 -66537 -106 -66525
rect 106 -65349 152 -65337
rect 106 -66525 112 -65349
rect 146 -66525 152 -65349
rect 106 -66537 152 -66525
rect -96 -66575 96 -66569
rect -96 -66609 -84 -66575
rect 84 -66609 96 -66575
rect -96 -66615 96 -66609
rect -96 -66683 96 -66677
rect -96 -66717 -84 -66683
rect 84 -66717 96 -66683
rect -96 -66723 96 -66717
rect -152 -66767 -106 -66755
rect -152 -67943 -146 -66767
rect -112 -67943 -106 -66767
rect -152 -67955 -106 -67943
rect 106 -66767 152 -66755
rect 106 -67943 112 -66767
rect 146 -67943 152 -66767
rect 106 -67955 152 -67943
rect -96 -67993 96 -67987
rect -96 -68027 -84 -67993
rect 84 -68027 96 -67993
rect -96 -68033 96 -68027
rect -96 -68101 96 -68095
rect -96 -68135 -84 -68101
rect 84 -68135 96 -68101
rect -96 -68141 96 -68135
rect -152 -68185 -106 -68173
rect -152 -69361 -146 -68185
rect -112 -69361 -106 -68185
rect -152 -69373 -106 -69361
rect 106 -68185 152 -68173
rect 106 -69361 112 -68185
rect 146 -69361 152 -68185
rect 106 -69373 152 -69361
rect -96 -69411 96 -69405
rect -96 -69445 -84 -69411
rect 84 -69445 96 -69411
rect -96 -69451 96 -69445
rect -96 -69519 96 -69513
rect -96 -69553 -84 -69519
rect 84 -69553 96 -69519
rect -96 -69559 96 -69553
rect -152 -69603 -106 -69591
rect -152 -70779 -146 -69603
rect -112 -70779 -106 -69603
rect -152 -70791 -106 -70779
rect 106 -69603 152 -69591
rect 106 -70779 112 -69603
rect 146 -70779 152 -69603
rect 106 -70791 152 -70779
rect -96 -70829 96 -70823
rect -96 -70863 -84 -70829
rect 84 -70863 96 -70829
rect -96 -70869 96 -70863
rect -96 -70937 96 -70931
rect -96 -70971 -84 -70937
rect 84 -70971 96 -70937
rect -96 -70977 96 -70971
rect -152 -71021 -106 -71009
rect -152 -72197 -146 -71021
rect -112 -72197 -106 -71021
rect -152 -72209 -106 -72197
rect 106 -71021 152 -71009
rect 106 -72197 112 -71021
rect 146 -72197 152 -71021
rect 106 -72209 152 -72197
rect -96 -72247 96 -72241
rect -96 -72281 -84 -72247
rect 84 -72281 96 -72247
rect -96 -72287 96 -72281
rect -96 -72355 96 -72349
rect -96 -72389 -84 -72355
rect 84 -72389 96 -72355
rect -96 -72395 96 -72389
rect -152 -72439 -106 -72427
rect -152 -73615 -146 -72439
rect -112 -73615 -106 -72439
rect -152 -73627 -106 -73615
rect 106 -72439 152 -72427
rect 106 -73615 112 -72439
rect 146 -73615 152 -72439
rect 106 -73627 152 -73615
rect -96 -73665 96 -73659
rect -96 -73699 -84 -73665
rect 84 -73699 96 -73665
rect -96 -73705 96 -73699
rect -96 -73773 96 -73767
rect -96 -73807 -84 -73773
rect 84 -73807 96 -73773
rect -96 -73813 96 -73807
rect -152 -73857 -106 -73845
rect -152 -75033 -146 -73857
rect -112 -75033 -106 -73857
rect -152 -75045 -106 -75033
rect 106 -73857 152 -73845
rect 106 -75033 112 -73857
rect 146 -75033 152 -73857
rect 106 -75045 152 -75033
rect -96 -75083 96 -75077
rect -96 -75117 -84 -75083
rect 84 -75117 96 -75083
rect -96 -75123 96 -75117
rect -96 -75191 96 -75185
rect -96 -75225 -84 -75191
rect 84 -75225 96 -75191
rect -96 -75231 96 -75225
rect -152 -75275 -106 -75263
rect -152 -76451 -146 -75275
rect -112 -76451 -106 -75275
rect -152 -76463 -106 -76451
rect 106 -75275 152 -75263
rect 106 -76451 112 -75275
rect 146 -76451 152 -75275
rect 106 -76463 152 -76451
rect -96 -76501 96 -76495
rect -96 -76535 -84 -76501
rect 84 -76535 96 -76501
rect -96 -76541 96 -76535
rect -96 -76609 96 -76603
rect -96 -76643 -84 -76609
rect 84 -76643 96 -76609
rect -96 -76649 96 -76643
rect -152 -76693 -106 -76681
rect -152 -77869 -146 -76693
rect -112 -77869 -106 -76693
rect -152 -77881 -106 -77869
rect 106 -76693 152 -76681
rect 106 -77869 112 -76693
rect 146 -77869 152 -76693
rect 106 -77881 152 -77869
rect -96 -77919 96 -77913
rect -96 -77953 -84 -77919
rect 84 -77953 96 -77919
rect -96 -77959 96 -77953
rect -96 -78027 96 -78021
rect -96 -78061 -84 -78027
rect 84 -78061 96 -78027
rect -96 -78067 96 -78061
rect -152 -78111 -106 -78099
rect -152 -79287 -146 -78111
rect -112 -79287 -106 -78111
rect -152 -79299 -106 -79287
rect 106 -78111 152 -78099
rect 106 -79287 112 -78111
rect 146 -79287 152 -78111
rect 106 -79299 152 -79287
rect -96 -79337 96 -79331
rect -96 -79371 -84 -79337
rect 84 -79371 96 -79337
rect -96 -79377 96 -79371
rect -96 -79445 96 -79439
rect -96 -79479 -84 -79445
rect 84 -79479 96 -79445
rect -96 -79485 96 -79479
rect -152 -79529 -106 -79517
rect -152 -80705 -146 -79529
rect -112 -80705 -106 -79529
rect -152 -80717 -106 -80705
rect 106 -79529 152 -79517
rect 106 -80705 112 -79529
rect 146 -80705 152 -79529
rect 106 -80717 152 -80705
rect -96 -80755 96 -80749
rect -96 -80789 -84 -80755
rect 84 -80789 96 -80755
rect -96 -80795 96 -80789
rect -96 -80863 96 -80857
rect -96 -80897 -84 -80863
rect 84 -80897 96 -80863
rect -96 -80903 96 -80897
rect -152 -80947 -106 -80935
rect -152 -82123 -146 -80947
rect -112 -82123 -106 -80947
rect -152 -82135 -106 -82123
rect 106 -80947 152 -80935
rect 106 -82123 112 -80947
rect 146 -82123 152 -80947
rect 106 -82135 152 -82123
rect -96 -82173 96 -82167
rect -96 -82207 -84 -82173
rect 84 -82207 96 -82173
rect -96 -82213 96 -82207
rect -96 -82281 96 -82275
rect -96 -82315 -84 -82281
rect 84 -82315 96 -82281
rect -96 -82321 96 -82315
rect -152 -82365 -106 -82353
rect -152 -83541 -146 -82365
rect -112 -83541 -106 -82365
rect -152 -83553 -106 -83541
rect 106 -82365 152 -82353
rect 106 -83541 112 -82365
rect 146 -83541 152 -82365
rect 106 -83553 152 -83541
rect -96 -83591 96 -83585
rect -96 -83625 -84 -83591
rect 84 -83625 96 -83591
rect -96 -83631 96 -83625
rect -96 -83699 96 -83693
rect -96 -83733 -84 -83699
rect 84 -83733 96 -83699
rect -96 -83739 96 -83733
rect -152 -83783 -106 -83771
rect -152 -84959 -146 -83783
rect -112 -84959 -106 -83783
rect -152 -84971 -106 -84959
rect 106 -83783 152 -83771
rect 106 -84959 112 -83783
rect 146 -84959 152 -83783
rect 106 -84971 152 -84959
rect -96 -85009 96 -85003
rect -96 -85043 -84 -85009
rect 84 -85043 96 -85009
rect -96 -85049 96 -85043
rect -96 -85117 96 -85111
rect -96 -85151 -84 -85117
rect 84 -85151 96 -85117
rect -96 -85157 96 -85151
rect -152 -85201 -106 -85189
rect -152 -86377 -146 -85201
rect -112 -86377 -106 -85201
rect -152 -86389 -106 -86377
rect 106 -85201 152 -85189
rect 106 -86377 112 -85201
rect 146 -86377 152 -85201
rect 106 -86389 152 -86377
rect -96 -86427 96 -86421
rect -96 -86461 -84 -86427
rect 84 -86461 96 -86427
rect -96 -86467 96 -86461
rect -96 -86535 96 -86529
rect -96 -86569 -84 -86535
rect 84 -86569 96 -86535
rect -96 -86575 96 -86569
rect -152 -86619 -106 -86607
rect -152 -87795 -146 -86619
rect -112 -87795 -106 -86619
rect -152 -87807 -106 -87795
rect 106 -86619 152 -86607
rect 106 -87795 112 -86619
rect 146 -87795 152 -86619
rect 106 -87807 152 -87795
rect -96 -87845 96 -87839
rect -96 -87879 -84 -87845
rect 84 -87879 96 -87845
rect -96 -87885 96 -87879
rect -96 -87953 96 -87947
rect -96 -87987 -84 -87953
rect 84 -87987 96 -87953
rect -96 -87993 96 -87987
rect -152 -88037 -106 -88025
rect -152 -89213 -146 -88037
rect -112 -89213 -106 -88037
rect -152 -89225 -106 -89213
rect 106 -88037 152 -88025
rect 106 -89213 112 -88037
rect 146 -89213 152 -88037
rect 106 -89225 152 -89213
rect -96 -89263 96 -89257
rect -96 -89297 -84 -89263
rect 84 -89297 96 -89263
rect -96 -89303 96 -89297
rect -96 -89371 96 -89365
rect -96 -89405 -84 -89371
rect 84 -89405 96 -89371
rect -96 -89411 96 -89405
rect -152 -89455 -106 -89443
rect -152 -90631 -146 -89455
rect -112 -90631 -106 -89455
rect -152 -90643 -106 -90631
rect 106 -89455 152 -89443
rect 106 -90631 112 -89455
rect 146 -90631 152 -89455
rect 106 -90643 152 -90631
rect -96 -90681 96 -90675
rect -96 -90715 -84 -90681
rect 84 -90715 96 -90681
rect -96 -90721 96 -90715
rect -96 -90789 96 -90783
rect -96 -90823 -84 -90789
rect 84 -90823 96 -90789
rect -96 -90829 96 -90823
rect -152 -90873 -106 -90861
rect -152 -92049 -146 -90873
rect -112 -92049 -106 -90873
rect -152 -92061 -106 -92049
rect 106 -90873 152 -90861
rect 106 -92049 112 -90873
rect 146 -92049 152 -90873
rect 106 -92061 152 -92049
rect -96 -92099 96 -92093
rect -96 -92133 -84 -92099
rect 84 -92133 96 -92099
rect -96 -92139 96 -92133
rect -96 -92207 96 -92201
rect -96 -92241 -84 -92207
rect 84 -92241 96 -92207
rect -96 -92247 96 -92241
rect -152 -92291 -106 -92279
rect -152 -93467 -146 -92291
rect -112 -93467 -106 -92291
rect -152 -93479 -106 -93467
rect 106 -92291 152 -92279
rect 106 -93467 112 -92291
rect 146 -93467 152 -92291
rect 106 -93479 152 -93467
rect -96 -93517 96 -93511
rect -96 -93551 -84 -93517
rect 84 -93551 96 -93517
rect -96 -93557 96 -93551
rect -96 -93625 96 -93619
rect -96 -93659 -84 -93625
rect 84 -93659 96 -93625
rect -96 -93665 96 -93659
rect -152 -93709 -106 -93697
rect -152 -94885 -146 -93709
rect -112 -94885 -106 -93709
rect -152 -94897 -106 -94885
rect 106 -93709 152 -93697
rect 106 -94885 112 -93709
rect 146 -94885 152 -93709
rect 106 -94897 152 -94885
rect -96 -94935 96 -94929
rect -96 -94969 -84 -94935
rect 84 -94969 96 -94935
rect -96 -94975 96 -94969
rect -96 -95043 96 -95037
rect -96 -95077 -84 -95043
rect 84 -95077 96 -95043
rect -96 -95083 96 -95077
rect -152 -95127 -106 -95115
rect -152 -96303 -146 -95127
rect -112 -96303 -106 -95127
rect -152 -96315 -106 -96303
rect 106 -95127 152 -95115
rect 106 -96303 112 -95127
rect 146 -96303 152 -95127
rect 106 -96315 152 -96303
rect -96 -96353 96 -96347
rect -96 -96387 -84 -96353
rect 84 -96387 96 -96353
rect -96 -96393 96 -96387
rect -96 -96461 96 -96455
rect -96 -96495 -84 -96461
rect 84 -96495 96 -96461
rect -96 -96501 96 -96495
rect -152 -96545 -106 -96533
rect -152 -97721 -146 -96545
rect -112 -97721 -106 -96545
rect -152 -97733 -106 -97721
rect 106 -96545 152 -96533
rect 106 -97721 112 -96545
rect 146 -97721 152 -96545
rect 106 -97733 152 -97721
rect -96 -97771 96 -97765
rect -96 -97805 -84 -97771
rect 84 -97805 96 -97771
rect -96 -97811 96 -97805
rect -96 -97879 96 -97873
rect -96 -97913 -84 -97879
rect 84 -97913 96 -97879
rect -96 -97919 96 -97913
rect -152 -97963 -106 -97951
rect -152 -99139 -146 -97963
rect -112 -99139 -106 -97963
rect -152 -99151 -106 -99139
rect 106 -97963 152 -97951
rect 106 -99139 112 -97963
rect 146 -99139 152 -97963
rect 106 -99151 152 -99139
rect -96 -99189 96 -99183
rect -96 -99223 -84 -99189
rect 84 -99223 96 -99189
rect -96 -99229 96 -99223
rect -96 -99297 96 -99291
rect -96 -99331 -84 -99297
rect 84 -99331 96 -99297
rect -96 -99337 96 -99331
rect -152 -99381 -106 -99369
rect -152 -100557 -146 -99381
rect -112 -100557 -106 -99381
rect -152 -100569 -106 -100557
rect 106 -99381 152 -99369
rect 106 -100557 112 -99381
rect 146 -100557 152 -99381
rect 106 -100569 152 -100557
rect -96 -100607 96 -100601
rect -96 -100641 -84 -100607
rect 84 -100641 96 -100607
rect -96 -100647 96 -100641
rect -96 -100715 96 -100709
rect -96 -100749 -84 -100715
rect 84 -100749 96 -100715
rect -96 -100755 96 -100749
rect -152 -100799 -106 -100787
rect -152 -101975 -146 -100799
rect -112 -101975 -106 -100799
rect -152 -101987 -106 -101975
rect 106 -100799 152 -100787
rect 106 -101975 112 -100799
rect 146 -101975 152 -100799
rect 106 -101987 152 -101975
rect -96 -102025 96 -102019
rect -96 -102059 -84 -102025
rect 84 -102059 96 -102025
rect -96 -102065 96 -102059
rect -96 -102133 96 -102127
rect -96 -102167 -84 -102133
rect 84 -102167 96 -102133
rect -96 -102173 96 -102167
rect -152 -102217 -106 -102205
rect -152 -103393 -146 -102217
rect -112 -103393 -106 -102217
rect -152 -103405 -106 -103393
rect 106 -102217 152 -102205
rect 106 -103393 112 -102217
rect 146 -103393 152 -102217
rect 106 -103405 152 -103393
rect -96 -103443 96 -103437
rect -96 -103477 -84 -103443
rect 84 -103477 96 -103443
rect -96 -103483 96 -103477
rect -96 -103551 96 -103545
rect -96 -103585 -84 -103551
rect 84 -103585 96 -103551
rect -96 -103591 96 -103585
rect -152 -103635 -106 -103623
rect -152 -104811 -146 -103635
rect -112 -104811 -106 -103635
rect -152 -104823 -106 -104811
rect 106 -103635 152 -103623
rect 106 -104811 112 -103635
rect 146 -104811 152 -103635
rect 106 -104823 152 -104811
rect -96 -104861 96 -104855
rect -96 -104895 -84 -104861
rect 84 -104895 96 -104861
rect -96 -104901 96 -104895
rect -96 -104969 96 -104963
rect -96 -105003 -84 -104969
rect 84 -105003 96 -104969
rect -96 -105009 96 -105003
rect -152 -105053 -106 -105041
rect -152 -106229 -146 -105053
rect -112 -106229 -106 -105053
rect -152 -106241 -106 -106229
rect 106 -105053 152 -105041
rect 106 -106229 112 -105053
rect 146 -106229 152 -105053
rect 106 -106241 152 -106229
rect -96 -106279 96 -106273
rect -96 -106313 -84 -106279
rect 84 -106313 96 -106279
rect -96 -106319 96 -106313
rect -96 -106387 96 -106381
rect -96 -106421 -84 -106387
rect 84 -106421 96 -106387
rect -96 -106427 96 -106421
rect -152 -106471 -106 -106459
rect -152 -107647 -146 -106471
rect -112 -107647 -106 -106471
rect -152 -107659 -106 -107647
rect 106 -106471 152 -106459
rect 106 -107647 112 -106471
rect 146 -107647 152 -106471
rect 106 -107659 152 -107647
rect -96 -107697 96 -107691
rect -96 -107731 -84 -107697
rect 84 -107731 96 -107697
rect -96 -107737 96 -107731
rect -96 -107805 96 -107799
rect -96 -107839 -84 -107805
rect 84 -107839 96 -107805
rect -96 -107845 96 -107839
rect -152 -107889 -106 -107877
rect -152 -109065 -146 -107889
rect -112 -109065 -106 -107889
rect -152 -109077 -106 -109065
rect 106 -107889 152 -107877
rect 106 -109065 112 -107889
rect 146 -109065 152 -107889
rect 106 -109077 152 -109065
rect -96 -109115 96 -109109
rect -96 -109149 -84 -109115
rect 84 -109149 96 -109115
rect -96 -109155 96 -109149
rect -96 -109223 96 -109217
rect -96 -109257 -84 -109223
rect 84 -109257 96 -109223
rect -96 -109263 96 -109257
rect -152 -109307 -106 -109295
rect -152 -110483 -146 -109307
rect -112 -110483 -106 -109307
rect -152 -110495 -106 -110483
rect 106 -109307 152 -109295
rect 106 -110483 112 -109307
rect 146 -110483 152 -109307
rect 106 -110495 152 -110483
rect -96 -110533 96 -110527
rect -96 -110567 -84 -110533
rect 84 -110567 96 -110533
rect -96 -110573 96 -110567
rect -96 -110641 96 -110635
rect -96 -110675 -84 -110641
rect 84 -110675 96 -110641
rect -96 -110681 96 -110675
rect -152 -110725 -106 -110713
rect -152 -111901 -146 -110725
rect -112 -111901 -106 -110725
rect -152 -111913 -106 -111901
rect 106 -110725 152 -110713
rect 106 -111901 112 -110725
rect 146 -111901 152 -110725
rect 106 -111913 152 -111901
rect -96 -111951 96 -111945
rect -96 -111985 -84 -111951
rect 84 -111985 96 -111951
rect -96 -111991 96 -111985
rect -96 -112059 96 -112053
rect -96 -112093 -84 -112059
rect 84 -112093 96 -112059
rect -96 -112099 96 -112093
rect -152 -112143 -106 -112131
rect -152 -113319 -146 -112143
rect -112 -113319 -106 -112143
rect -152 -113331 -106 -113319
rect 106 -112143 152 -112131
rect 106 -113319 112 -112143
rect 146 -113319 152 -112143
rect 106 -113331 152 -113319
rect -96 -113369 96 -113363
rect -96 -113403 -84 -113369
rect 84 -113403 96 -113369
rect -96 -113409 96 -113403
rect -96 -113477 96 -113471
rect -96 -113511 -84 -113477
rect 84 -113511 96 -113477
rect -96 -113517 96 -113511
rect -152 -113561 -106 -113549
rect -152 -114737 -146 -113561
rect -112 -114737 -106 -113561
rect -152 -114749 -106 -114737
rect 106 -113561 152 -113549
rect 106 -114737 112 -113561
rect 146 -114737 152 -113561
rect 106 -114749 152 -114737
rect -96 -114787 96 -114781
rect -96 -114821 -84 -114787
rect 84 -114821 96 -114787
rect -96 -114827 96 -114821
rect -96 -114895 96 -114889
rect -96 -114929 -84 -114895
rect 84 -114929 96 -114895
rect -96 -114935 96 -114929
rect -152 -114979 -106 -114967
rect -152 -116155 -146 -114979
rect -112 -116155 -106 -114979
rect -152 -116167 -106 -116155
rect 106 -114979 152 -114967
rect 106 -116155 112 -114979
rect 146 -116155 152 -114979
rect 106 -116167 152 -116155
rect -96 -116205 96 -116199
rect -96 -116239 -84 -116205
rect 84 -116239 96 -116205
rect -96 -116245 96 -116239
rect -96 -116313 96 -116307
rect -96 -116347 -84 -116313
rect 84 -116347 96 -116313
rect -96 -116353 96 -116347
rect -152 -116397 -106 -116385
rect -152 -117573 -146 -116397
rect -112 -117573 -106 -116397
rect -152 -117585 -106 -117573
rect 106 -116397 152 -116385
rect 106 -117573 112 -116397
rect 146 -117573 152 -116397
rect 106 -117585 152 -117573
rect -96 -117623 96 -117617
rect -96 -117657 -84 -117623
rect 84 -117657 96 -117623
rect -96 -117663 96 -117657
rect -96 -117731 96 -117725
rect -96 -117765 -84 -117731
rect 84 -117765 96 -117731
rect -96 -117771 96 -117765
rect -152 -117815 -106 -117803
rect -152 -118991 -146 -117815
rect -112 -118991 -106 -117815
rect -152 -119003 -106 -118991
rect 106 -117815 152 -117803
rect 106 -118991 112 -117815
rect 146 -118991 152 -117815
rect 106 -119003 152 -118991
rect -96 -119041 96 -119035
rect -96 -119075 -84 -119041
rect 84 -119075 96 -119041
rect -96 -119081 96 -119075
rect -96 -119149 96 -119143
rect -96 -119183 -84 -119149
rect 84 -119183 96 -119149
rect -96 -119189 96 -119183
rect -152 -119233 -106 -119221
rect -152 -120409 -146 -119233
rect -112 -120409 -106 -119233
rect -152 -120421 -106 -120409
rect 106 -119233 152 -119221
rect 106 -120409 112 -119233
rect 146 -120409 152 -119233
rect 106 -120421 152 -120409
rect -96 -120459 96 -120453
rect -96 -120493 -84 -120459
rect 84 -120493 96 -120459
rect -96 -120499 96 -120493
rect -96 -120567 96 -120561
rect -96 -120601 -84 -120567
rect 84 -120601 96 -120567
rect -96 -120607 96 -120601
rect -152 -120651 -106 -120639
rect -152 -121827 -146 -120651
rect -112 -121827 -106 -120651
rect -152 -121839 -106 -121827
rect 106 -120651 152 -120639
rect 106 -121827 112 -120651
rect 146 -121827 152 -120651
rect 106 -121839 152 -121827
rect -96 -121877 96 -121871
rect -96 -121911 -84 -121877
rect 84 -121911 96 -121877
rect -96 -121917 96 -121911
rect -96 -121985 96 -121979
rect -96 -122019 -84 -121985
rect 84 -122019 96 -121985
rect -96 -122025 96 -122019
rect -152 -122069 -106 -122057
rect -152 -123245 -146 -122069
rect -112 -123245 -106 -122069
rect -152 -123257 -106 -123245
rect 106 -122069 152 -122057
rect 106 -123245 112 -122069
rect 146 -123245 152 -122069
rect 106 -123257 152 -123245
rect -96 -123295 96 -123289
rect -96 -123329 -84 -123295
rect 84 -123329 96 -123295
rect -96 -123335 96 -123329
rect -96 -123403 96 -123397
rect -96 -123437 -84 -123403
rect 84 -123437 96 -123403
rect -96 -123443 96 -123437
rect -152 -123487 -106 -123475
rect -152 -124663 -146 -123487
rect -112 -124663 -106 -123487
rect -152 -124675 -106 -124663
rect 106 -123487 152 -123475
rect 106 -124663 112 -123487
rect 146 -124663 152 -123487
rect 106 -124675 152 -124663
rect -96 -124713 96 -124707
rect -96 -124747 -84 -124713
rect 84 -124747 96 -124713
rect -96 -124753 96 -124747
rect -96 -124821 96 -124815
rect -96 -124855 -84 -124821
rect 84 -124855 96 -124821
rect -96 -124861 96 -124855
rect -152 -124905 -106 -124893
rect -152 -126081 -146 -124905
rect -112 -126081 -106 -124905
rect -152 -126093 -106 -126081
rect 106 -124905 152 -124893
rect 106 -126081 112 -124905
rect 146 -126081 152 -124905
rect 106 -126093 152 -126081
rect -96 -126131 96 -126125
rect -96 -126165 -84 -126131
rect 84 -126165 96 -126131
rect -96 -126171 96 -126165
rect -96 -126239 96 -126233
rect -96 -126273 -84 -126239
rect 84 -126273 96 -126239
rect -96 -126279 96 -126273
rect -152 -126323 -106 -126311
rect -152 -127499 -146 -126323
rect -112 -127499 -106 -126323
rect -152 -127511 -106 -127499
rect 106 -126323 152 -126311
rect 106 -127499 112 -126323
rect 146 -127499 152 -126323
rect 106 -127511 152 -127499
rect -96 -127549 96 -127543
rect -96 -127583 -84 -127549
rect 84 -127583 96 -127549
rect -96 -127589 96 -127583
rect -96 -127657 96 -127651
rect -96 -127691 -84 -127657
rect 84 -127691 96 -127657
rect -96 -127697 96 -127691
rect -152 -127741 -106 -127729
rect -152 -128917 -146 -127741
rect -112 -128917 -106 -127741
rect -152 -128929 -106 -128917
rect 106 -127741 152 -127729
rect 106 -128917 112 -127741
rect 146 -128917 152 -127741
rect 106 -128929 152 -128917
rect -96 -128967 96 -128961
rect -96 -129001 -84 -128967
rect 84 -129001 96 -128967
rect -96 -129007 96 -129001
rect -96 -129075 96 -129069
rect -96 -129109 -84 -129075
rect 84 -129109 96 -129075
rect -96 -129115 96 -129109
rect -152 -129159 -106 -129147
rect -152 -130335 -146 -129159
rect -112 -130335 -106 -129159
rect -152 -130347 -106 -130335
rect 106 -129159 152 -129147
rect 106 -130335 112 -129159
rect 146 -130335 152 -129159
rect 106 -130347 152 -130335
rect -96 -130385 96 -130379
rect -96 -130419 -84 -130385
rect 84 -130419 96 -130385
rect -96 -130425 96 -130419
rect -96 -130493 96 -130487
rect -96 -130527 -84 -130493
rect 84 -130527 96 -130493
rect -96 -130533 96 -130527
rect -152 -130577 -106 -130565
rect -152 -131753 -146 -130577
rect -112 -131753 -106 -130577
rect -152 -131765 -106 -131753
rect 106 -130577 152 -130565
rect 106 -131753 112 -130577
rect 146 -131753 152 -130577
rect 106 -131765 152 -131753
rect -96 -131803 96 -131797
rect -96 -131837 -84 -131803
rect 84 -131837 96 -131803
rect -96 -131843 96 -131837
rect -96 -131911 96 -131905
rect -96 -131945 -84 -131911
rect 84 -131945 96 -131911
rect -96 -131951 96 -131945
rect -152 -131995 -106 -131983
rect -152 -133171 -146 -131995
rect -112 -133171 -106 -131995
rect -152 -133183 -106 -133171
rect 106 -131995 152 -131983
rect 106 -133171 112 -131995
rect 146 -133171 152 -131995
rect 106 -133183 152 -133171
rect -96 -133221 96 -133215
rect -96 -133255 -84 -133221
rect 84 -133255 96 -133221
rect -96 -133261 96 -133255
rect -96 -133329 96 -133323
rect -96 -133363 -84 -133329
rect 84 -133363 96 -133329
rect -96 -133369 96 -133363
rect -152 -133413 -106 -133401
rect -152 -134589 -146 -133413
rect -112 -134589 -106 -133413
rect -152 -134601 -106 -134589
rect 106 -133413 152 -133401
rect 106 -134589 112 -133413
rect 146 -134589 152 -133413
rect 106 -134601 152 -134589
rect -96 -134639 96 -134633
rect -96 -134673 -84 -134639
rect 84 -134673 96 -134639
rect -96 -134679 96 -134673
rect -96 -134747 96 -134741
rect -96 -134781 -84 -134747
rect 84 -134781 96 -134747
rect -96 -134787 96 -134781
rect -152 -134831 -106 -134819
rect -152 -136007 -146 -134831
rect -112 -136007 -106 -134831
rect -152 -136019 -106 -136007
rect 106 -134831 152 -134819
rect 106 -136007 112 -134831
rect 146 -136007 152 -134831
rect 106 -136019 152 -136007
rect -96 -136057 96 -136051
rect -96 -136091 -84 -136057
rect 84 -136091 96 -136057
rect -96 -136097 96 -136091
rect -96 -136165 96 -136159
rect -96 -136199 -84 -136165
rect 84 -136199 96 -136165
rect -96 -136205 96 -136199
rect -152 -136249 -106 -136237
rect -152 -137425 -146 -136249
rect -112 -137425 -106 -136249
rect -152 -137437 -106 -137425
rect 106 -136249 152 -136237
rect 106 -137425 112 -136249
rect 146 -137425 152 -136249
rect 106 -137437 152 -137425
rect -96 -137475 96 -137469
rect -96 -137509 -84 -137475
rect 84 -137509 96 -137475
rect -96 -137515 96 -137509
rect -96 -137583 96 -137577
rect -96 -137617 -84 -137583
rect 84 -137617 96 -137583
rect -96 -137623 96 -137617
rect -152 -137667 -106 -137655
rect -152 -138843 -146 -137667
rect -112 -138843 -106 -137667
rect -152 -138855 -106 -138843
rect 106 -137667 152 -137655
rect 106 -138843 112 -137667
rect 146 -138843 152 -137667
rect 106 -138855 152 -138843
rect -96 -138893 96 -138887
rect -96 -138927 -84 -138893
rect 84 -138927 96 -138893
rect -96 -138933 96 -138927
rect -96 -139001 96 -138995
rect -96 -139035 -84 -139001
rect 84 -139035 96 -139001
rect -96 -139041 96 -139035
rect -152 -139085 -106 -139073
rect -152 -140261 -146 -139085
rect -112 -140261 -106 -139085
rect -152 -140273 -106 -140261
rect 106 -139085 152 -139073
rect 106 -140261 112 -139085
rect 146 -140261 152 -139085
rect 106 -140273 152 -140261
rect -96 -140311 96 -140305
rect -96 -140345 -84 -140311
rect 84 -140345 96 -140311
rect -96 -140351 96 -140345
rect -96 -140419 96 -140413
rect -96 -140453 -84 -140419
rect 84 -140453 96 -140419
rect -96 -140459 96 -140453
rect -152 -140503 -106 -140491
rect -152 -141679 -146 -140503
rect -112 -141679 -106 -140503
rect -152 -141691 -106 -141679
rect 106 -140503 152 -140491
rect 106 -141679 112 -140503
rect 146 -141679 152 -140503
rect 106 -141691 152 -141679
rect -96 -141729 96 -141723
rect -96 -141763 -84 -141729
rect 84 -141763 96 -141729
rect -96 -141769 96 -141763
rect -96 -141837 96 -141831
rect -96 -141871 -84 -141837
rect 84 -141871 96 -141837
rect -96 -141877 96 -141871
rect -152 -141921 -106 -141909
rect -152 -143097 -146 -141921
rect -112 -143097 -106 -141921
rect -152 -143109 -106 -143097
rect 106 -141921 152 -141909
rect 106 -143097 112 -141921
rect 146 -143097 152 -141921
rect 106 -143109 152 -143097
rect -96 -143147 96 -143141
rect -96 -143181 -84 -143147
rect 84 -143181 96 -143147
rect -96 -143187 96 -143181
rect -96 -143255 96 -143249
rect -96 -143289 -84 -143255
rect 84 -143289 96 -143255
rect -96 -143295 96 -143289
rect -152 -143339 -106 -143327
rect -152 -144515 -146 -143339
rect -112 -144515 -106 -143339
rect -152 -144527 -106 -144515
rect 106 -143339 152 -143327
rect 106 -144515 112 -143339
rect 146 -144515 152 -143339
rect 106 -144527 152 -144515
rect -96 -144565 96 -144559
rect -96 -144599 -84 -144565
rect 84 -144599 96 -144565
rect -96 -144605 96 -144599
rect -96 -144673 96 -144667
rect -96 -144707 -84 -144673
rect 84 -144707 96 -144673
rect -96 -144713 96 -144707
rect -152 -144757 -106 -144745
rect -152 -145933 -146 -144757
rect -112 -145933 -106 -144757
rect -152 -145945 -106 -145933
rect 106 -144757 152 -144745
rect 106 -145933 112 -144757
rect 146 -145933 152 -144757
rect 106 -145945 152 -145933
rect -96 -145983 96 -145977
rect -96 -146017 -84 -145983
rect 84 -146017 96 -145983
rect -96 -146023 96 -146017
rect -96 -146091 96 -146085
rect -96 -146125 -84 -146091
rect 84 -146125 96 -146091
rect -96 -146131 96 -146125
rect -152 -146175 -106 -146163
rect -152 -147351 -146 -146175
rect -112 -147351 -106 -146175
rect -152 -147363 -106 -147351
rect 106 -146175 152 -146163
rect 106 -147351 112 -146175
rect 146 -147351 152 -146175
rect 106 -147363 152 -147351
rect -96 -147401 96 -147395
rect -96 -147435 -84 -147401
rect 84 -147435 96 -147401
rect -96 -147441 96 -147435
rect -96 -147509 96 -147503
rect -96 -147543 -84 -147509
rect 84 -147543 96 -147509
rect -96 -147549 96 -147543
rect -152 -147593 -106 -147581
rect -152 -148769 -146 -147593
rect -112 -148769 -106 -147593
rect -152 -148781 -106 -148769
rect 106 -147593 152 -147581
rect 106 -148769 112 -147593
rect 146 -148769 152 -147593
rect 106 -148781 152 -148769
rect -96 -148819 96 -148813
rect -96 -148853 -84 -148819
rect 84 -148853 96 -148819
rect -96 -148859 96 -148853
rect -96 -148927 96 -148921
rect -96 -148961 -84 -148927
rect 84 -148961 96 -148927
rect -96 -148967 96 -148961
rect -152 -149011 -106 -148999
rect -152 -150187 -146 -149011
rect -112 -150187 -106 -149011
rect -152 -150199 -106 -150187
rect 106 -149011 152 -148999
rect 106 -150187 112 -149011
rect 146 -150187 152 -149011
rect 106 -150199 152 -150187
rect -96 -150237 96 -150231
rect -96 -150271 -84 -150237
rect 84 -150271 96 -150237
rect -96 -150277 96 -150271
rect -96 -150345 96 -150339
rect -96 -150379 -84 -150345
rect 84 -150379 96 -150345
rect -96 -150385 96 -150379
rect -152 -150429 -106 -150417
rect -152 -151605 -146 -150429
rect -112 -151605 -106 -150429
rect -152 -151617 -106 -151605
rect 106 -150429 152 -150417
rect 106 -151605 112 -150429
rect 146 -151605 152 -150429
rect 106 -151617 152 -151605
rect -96 -151655 96 -151649
rect -96 -151689 -84 -151655
rect 84 -151689 96 -151655
rect -96 -151695 96 -151689
rect -96 -151763 96 -151757
rect -96 -151797 -84 -151763
rect 84 -151797 96 -151763
rect -96 -151803 96 -151797
rect -152 -151847 -106 -151835
rect -152 -153023 -146 -151847
rect -112 -153023 -106 -151847
rect -152 -153035 -106 -153023
rect 106 -151847 152 -151835
rect 106 -153023 112 -151847
rect 146 -153023 152 -151847
rect 106 -153035 152 -153023
rect -96 -153073 96 -153067
rect -96 -153107 -84 -153073
rect 84 -153107 96 -153073
rect -96 -153113 96 -153107
rect -96 -153181 96 -153175
rect -96 -153215 -84 -153181
rect 84 -153215 96 -153181
rect -96 -153221 96 -153215
rect -152 -153265 -106 -153253
rect -152 -154441 -146 -153265
rect -112 -154441 -106 -153265
rect -152 -154453 -106 -154441
rect 106 -153265 152 -153253
rect 106 -154441 112 -153265
rect 146 -154441 152 -153265
rect 106 -154453 152 -154441
rect -96 -154491 96 -154485
rect -96 -154525 -84 -154491
rect 84 -154525 96 -154491
rect -96 -154531 96 -154525
rect -96 -154599 96 -154593
rect -96 -154633 -84 -154599
rect 84 -154633 96 -154599
rect -96 -154639 96 -154633
rect -152 -154683 -106 -154671
rect -152 -155859 -146 -154683
rect -112 -155859 -106 -154683
rect -152 -155871 -106 -155859
rect 106 -154683 152 -154671
rect 106 -155859 112 -154683
rect 146 -155859 152 -154683
rect 106 -155871 152 -155859
rect -96 -155909 96 -155903
rect -96 -155943 -84 -155909
rect 84 -155943 96 -155909
rect -96 -155949 96 -155943
rect -96 -156017 96 -156011
rect -96 -156051 -84 -156017
rect 84 -156051 96 -156017
rect -96 -156057 96 -156051
rect -152 -156101 -106 -156089
rect -152 -157277 -146 -156101
rect -112 -157277 -106 -156101
rect -152 -157289 -106 -157277
rect 106 -156101 152 -156089
rect 106 -157277 112 -156101
rect 146 -157277 152 -156101
rect 106 -157289 152 -157277
rect -96 -157327 96 -157321
rect -96 -157361 -84 -157327
rect 84 -157361 96 -157327
rect -96 -157367 96 -157361
rect -96 -157435 96 -157429
rect -96 -157469 -84 -157435
rect 84 -157469 96 -157435
rect -96 -157475 96 -157469
rect -152 -157519 -106 -157507
rect -152 -158695 -146 -157519
rect -112 -158695 -106 -157519
rect -152 -158707 -106 -158695
rect 106 -157519 152 -157507
rect 106 -158695 112 -157519
rect 146 -158695 152 -157519
rect 106 -158707 152 -158695
rect -96 -158745 96 -158739
rect -96 -158779 -84 -158745
rect 84 -158779 96 -158745
rect -96 -158785 96 -158779
rect -96 -158853 96 -158847
rect -96 -158887 -84 -158853
rect 84 -158887 96 -158853
rect -96 -158893 96 -158887
rect -152 -158937 -106 -158925
rect -152 -160113 -146 -158937
rect -112 -160113 -106 -158937
rect -152 -160125 -106 -160113
rect 106 -158937 152 -158925
rect 106 -160113 112 -158937
rect 146 -160113 152 -158937
rect 106 -160125 152 -160113
rect -96 -160163 96 -160157
rect -96 -160197 -84 -160163
rect 84 -160197 96 -160163
rect -96 -160203 96 -160197
rect -96 -160271 96 -160265
rect -96 -160305 -84 -160271
rect 84 -160305 96 -160271
rect -96 -160311 96 -160305
rect -152 -160355 -106 -160343
rect -152 -161531 -146 -160355
rect -112 -161531 -106 -160355
rect -152 -161543 -106 -161531
rect 106 -160355 152 -160343
rect 106 -161531 112 -160355
rect 146 -161531 152 -160355
rect 106 -161543 152 -161531
rect -96 -161581 96 -161575
rect -96 -161615 -84 -161581
rect 84 -161615 96 -161581
rect -96 -161621 96 -161615
rect -96 -161689 96 -161683
rect -96 -161723 -84 -161689
rect 84 -161723 96 -161689
rect -96 -161729 96 -161723
rect -152 -161773 -106 -161761
rect -152 -162949 -146 -161773
rect -112 -162949 -106 -161773
rect -152 -162961 -106 -162949
rect 106 -161773 152 -161761
rect 106 -162949 112 -161773
rect 146 -162949 152 -161773
rect 106 -162961 152 -162949
rect -96 -162999 96 -162993
rect -96 -163033 -84 -162999
rect 84 -163033 96 -162999
rect -96 -163039 96 -163033
rect -96 -163107 96 -163101
rect -96 -163141 -84 -163107
rect 84 -163141 96 -163107
rect -96 -163147 96 -163141
rect -152 -163191 -106 -163179
rect -152 -164367 -146 -163191
rect -112 -164367 -106 -163191
rect -152 -164379 -106 -164367
rect 106 -163191 152 -163179
rect 106 -164367 112 -163191
rect 146 -164367 152 -163191
rect 106 -164379 152 -164367
rect -96 -164417 96 -164411
rect -96 -164451 -84 -164417
rect 84 -164451 96 -164417
rect -96 -164457 96 -164451
rect -96 -164525 96 -164519
rect -96 -164559 -84 -164525
rect 84 -164559 96 -164525
rect -96 -164565 96 -164559
rect -152 -164609 -106 -164597
rect -152 -165785 -146 -164609
rect -112 -165785 -106 -164609
rect -152 -165797 -106 -165785
rect 106 -164609 152 -164597
rect 106 -165785 112 -164609
rect 146 -165785 152 -164609
rect 106 -165797 152 -165785
rect -96 -165835 96 -165829
rect -96 -165869 -84 -165835
rect 84 -165869 96 -165835
rect -96 -165875 96 -165869
rect -96 -165943 96 -165937
rect -96 -165977 -84 -165943
rect 84 -165977 96 -165943
rect -96 -165983 96 -165977
rect -152 -166027 -106 -166015
rect -152 -167203 -146 -166027
rect -112 -167203 -106 -166027
rect -152 -167215 -106 -167203
rect 106 -166027 152 -166015
rect 106 -167203 112 -166027
rect 146 -167203 152 -166027
rect 106 -167215 152 -167203
rect -96 -167253 96 -167247
rect -96 -167287 -84 -167253
rect 84 -167287 96 -167253
rect -96 -167293 96 -167287
rect -96 -167361 96 -167355
rect -96 -167395 -84 -167361
rect 84 -167395 96 -167361
rect -96 -167401 96 -167395
rect -152 -167445 -106 -167433
rect -152 -168621 -146 -167445
rect -112 -168621 -106 -167445
rect -152 -168633 -106 -168621
rect 106 -167445 152 -167433
rect 106 -168621 112 -167445
rect 146 -168621 152 -167445
rect 106 -168633 152 -168621
rect -96 -168671 96 -168665
rect -96 -168705 -84 -168671
rect 84 -168705 96 -168671
rect -96 -168711 96 -168705
rect -96 -168779 96 -168773
rect -96 -168813 -84 -168779
rect 84 -168813 96 -168779
rect -96 -168819 96 -168813
rect -152 -168863 -106 -168851
rect -152 -170039 -146 -168863
rect -112 -170039 -106 -168863
rect -152 -170051 -106 -170039
rect 106 -168863 152 -168851
rect 106 -170039 112 -168863
rect 146 -170039 152 -168863
rect 106 -170051 152 -170039
rect -96 -170089 96 -170083
rect -96 -170123 -84 -170089
rect 84 -170123 96 -170089
rect -96 -170129 96 -170123
rect -96 -170197 96 -170191
rect -96 -170231 -84 -170197
rect 84 -170231 96 -170197
rect -96 -170237 96 -170231
rect -152 -170281 -106 -170269
rect -152 -171457 -146 -170281
rect -112 -171457 -106 -170281
rect -152 -171469 -106 -171457
rect 106 -170281 152 -170269
rect 106 -171457 112 -170281
rect 146 -171457 152 -170281
rect 106 -171469 152 -171457
rect -96 -171507 96 -171501
rect -96 -171541 -84 -171507
rect 84 -171541 96 -171507
rect -96 -171547 96 -171541
rect -96 -171615 96 -171609
rect -96 -171649 -84 -171615
rect 84 -171649 96 -171615
rect -96 -171655 96 -171649
rect -152 -171699 -106 -171687
rect -152 -172875 -146 -171699
rect -112 -172875 -106 -171699
rect -152 -172887 -106 -172875
rect 106 -171699 152 -171687
rect 106 -172875 112 -171699
rect 146 -172875 152 -171699
rect 106 -172887 152 -172875
rect -96 -172925 96 -172919
rect -96 -172959 -84 -172925
rect 84 -172959 96 -172925
rect -96 -172965 96 -172959
rect -96 -173033 96 -173027
rect -96 -173067 -84 -173033
rect 84 -173067 96 -173033
rect -96 -173073 96 -173067
rect -152 -173117 -106 -173105
rect -152 -174293 -146 -173117
rect -112 -174293 -106 -173117
rect -152 -174305 -106 -174293
rect 106 -173117 152 -173105
rect 106 -174293 112 -173117
rect 146 -174293 152 -173117
rect 106 -174305 152 -174293
rect -96 -174343 96 -174337
rect -96 -174377 -84 -174343
rect 84 -174377 96 -174343
rect -96 -174383 96 -174377
rect -96 -174451 96 -174445
rect -96 -174485 -84 -174451
rect 84 -174485 96 -174451
rect -96 -174491 96 -174485
rect -152 -174535 -106 -174523
rect -152 -175711 -146 -174535
rect -112 -175711 -106 -174535
rect -152 -175723 -106 -175711
rect 106 -174535 152 -174523
rect 106 -175711 112 -174535
rect 146 -175711 152 -174535
rect 106 -175723 152 -175711
rect -96 -175761 96 -175755
rect -96 -175795 -84 -175761
rect 84 -175795 96 -175761
rect -96 -175801 96 -175795
rect -96 -175869 96 -175863
rect -96 -175903 -84 -175869
rect 84 -175903 96 -175869
rect -96 -175909 96 -175903
rect -152 -175953 -106 -175941
rect -152 -177129 -146 -175953
rect -112 -177129 -106 -175953
rect -152 -177141 -106 -177129
rect 106 -175953 152 -175941
rect 106 -177129 112 -175953
rect 146 -177129 152 -175953
rect 106 -177141 152 -177129
rect -96 -177179 96 -177173
rect -96 -177213 -84 -177179
rect 84 -177213 96 -177179
rect -96 -177219 96 -177213
rect -96 -177287 96 -177281
rect -96 -177321 -84 -177287
rect 84 -177321 96 -177287
rect -96 -177327 96 -177321
rect -152 -177371 -106 -177359
rect -152 -178547 -146 -177371
rect -112 -178547 -106 -177371
rect -152 -178559 -106 -178547
rect 106 -177371 152 -177359
rect 106 -178547 112 -177371
rect 146 -178547 152 -177371
rect 106 -178559 152 -178547
rect -96 -178597 96 -178591
rect -96 -178631 -84 -178597
rect 84 -178631 96 -178597
rect -96 -178637 96 -178631
rect -96 -178705 96 -178699
rect -96 -178739 -84 -178705
rect 84 -178739 96 -178705
rect -96 -178745 96 -178739
rect -152 -178789 -106 -178777
rect -152 -179965 -146 -178789
rect -112 -179965 -106 -178789
rect -152 -179977 -106 -179965
rect 106 -178789 152 -178777
rect 106 -179965 112 -178789
rect 146 -179965 152 -178789
rect 106 -179977 152 -179965
rect -96 -180015 96 -180009
rect -96 -180049 -84 -180015
rect 84 -180049 96 -180015
rect -96 -180055 96 -180049
rect -96 -180123 96 -180117
rect -96 -180157 -84 -180123
rect 84 -180157 96 -180123
rect -96 -180163 96 -180157
rect -152 -180207 -106 -180195
rect -152 -181383 -146 -180207
rect -112 -181383 -106 -180207
rect -152 -181395 -106 -181383
rect 106 -180207 152 -180195
rect 106 -181383 112 -180207
rect 146 -181383 152 -180207
rect 106 -181395 152 -181383
rect -96 -181433 96 -181427
rect -96 -181467 -84 -181433
rect 84 -181467 96 -181433
rect -96 -181473 96 -181467
<< properties >>
string FIXED_BBOX -263 -181588 263 181588
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 6.0 l 1.0 m 256 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
