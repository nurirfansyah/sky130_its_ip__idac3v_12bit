magic
tech sky130A
magscale 1 2
timestamp 1717441772
<< metal1 >>
rect 121049 -18777 121247 -10275
rect 121279 -16560 121476 -7744
rect 121506 -18684 121703 -7927
rect 121733 -17865 121931 -7749
rect 121962 -16567 122160 -8461
rect 122191 -18092 122388 -9408
rect 122420 -18093 122615 -8975
rect 122650 -18313 122841 -10023
use icell64scs  x1
timestamp 1717439915
transform 1 0 0 0 1 0
box 4823 -12682 122844 2790
use icell64scs  x2
timestamp 1717439915
transform 1 0 1 0 1 -15044
box 4823 -12682 122844 2790
<< end >>
