magic
tech sky130A
timestamp 1717438951
<< metal1 >>
rect 2432 1181 2532 1281
rect 2432 -315 2532 -215
rect 4045 -657 4524 -557
use icell1scs  x1
timestamp 1717438951
transform 1 0 3663 0 1 129
box 584 -2709 2420 1266
use icell1scs  x2
timestamp 1717438951
transform 1 0 1848 0 1 129
box 584 -2709 2420 1266
<< labels >>
flabel metal1 s 2432 1229 2432 1229 3 FreeSans 800 0 0 0 iout
port 0 e
flabel metal1 2432 -265 2432 -265 3 FreeSans 800 0 0 0 avdd
port 1 e
flabel space 2432 1342 2432 1342 3 FreeSans 800 0 0 0 ioutn
port 3 e
flabel metal1 s 2609 -603 2609 -603 3 FreeSans 800 0 0 0 sw
port 4 e
flabel space 2433 -499 2433 -499 3 FreeSans 800 0 0 0 pcbias
port 5 e
flabel space 2431 -379 2431 -379 3 FreeSans 800 0 0 0 pbias
port 2 e
flabel space 2432 -1189 2432 -1189 3 FreeSans 800 0 0 0 idir_sel
port 6 e
flabel space 2433 -1301 2433 -1301 3 FreeSans 800 0 0 0 ncbias
port 7 e
flabel space 2432 -1409 2432 -1409 3 FreeSans 800 0 0 0 nbias
port 8 e
flabel space 2432 -1533 2432 -1533 3 FreeSans 800 0 0 0 avss
port 9 e
<< end >>
