magic
tech sky130A
magscale 1 2
timestamp 1717438773
<< nwell >>
rect 1148 -522 1212 -322
rect 1860 -522 1868 -322
rect 2576 -506 2642 -334
<< viali >>
rect 1598 1742 1966 1778
<< metal1 >>
rect 710 2382 3380 2388
rect 710 2200 1698 2382
rect 1866 2200 3380 2382
rect 710 2188 3380 2200
rect 710 2152 3380 2160
rect 710 1970 984 2152
rect 1152 1970 3380 2152
rect 710 1960 3380 1970
rect 710 1924 3380 1932
rect 710 1740 876 1924
rect 928 1778 3380 1924
rect 928 1742 1598 1778
rect 1966 1742 3380 1778
rect 928 1740 3380 1742
rect 710 1732 3380 1740
rect 1692 1658 1872 1664
rect 1692 1606 1698 1658
rect 1866 1606 1872 1658
rect 1692 1600 1872 1606
rect 978 458 1158 464
rect 978 406 984 458
rect 1152 406 1158 458
rect 978 400 1158 406
rect 2406 58 2586 64
rect 2406 6 2412 58
rect 2580 6 2586 58
rect 2406 0 2586 6
rect 2932 58 3112 64
rect 2932 6 2938 58
rect 3106 6 3112 58
rect 2932 0 3112 6
rect 904 -342 970 -336
rect 904 -502 910 -342
rect 964 -502 970 -342
rect 904 -508 970 -502
rect 1148 -340 1212 -322
rect 1148 -502 1154 -340
rect 1610 -342 1704 -322
rect 1610 -502 1636 -342
rect 1696 -502 1704 -342
rect 1148 -522 1212 -502
rect 1610 -522 1704 -502
rect 1868 -342 1934 -322
rect 2602 -334 2916 -42
rect 1928 -502 1934 -342
rect 1868 -522 1934 -502
rect 2576 -340 2916 -334
rect 2576 -500 2582 -340
rect 2642 -500 2916 -340
rect 2576 -506 2916 -500
rect 2332 -582 2396 -576
rect 2332 -742 2338 -582
rect 2390 -742 2396 -582
rect 2332 -748 2396 -742
rect 2602 -840 2916 -506
rect 3128 -340 3180 -40
rect 3128 -842 3180 -500
rect 710 -1068 3380 -1060
rect 710 -1252 2338 -1068
rect 2390 -1252 3380 -1068
rect 710 -1260 3380 -1252
rect 710 -1296 3380 -1288
rect 710 -1480 3128 -1296
rect 3180 -1480 3380 -1296
rect 710 -1488 3380 -1480
<< via1 >>
rect 1698 2200 1866 2382
rect 984 1970 1152 2152
rect 876 1740 928 1924
rect 1698 1606 1866 1658
rect 984 406 1152 458
rect 2412 6 2580 58
rect 2938 6 3106 58
rect 910 -502 964 -342
rect 1154 -502 1214 -340
rect 1636 -502 1696 -342
rect 1868 -502 1928 -342
rect 2582 -500 2642 -340
rect 2338 -742 2390 -582
rect 3128 -500 3180 -340
rect 2338 -1252 2390 -1068
rect 3128 -1480 3180 -1296
<< metal2 >>
rect 1692 2382 1872 2388
rect 1692 2200 1698 2382
rect 1866 2200 1872 2382
rect 978 2152 1158 2160
rect 978 1970 984 2152
rect 1152 1970 1158 2152
rect 870 1924 934 1932
rect 870 1740 876 1924
rect 928 1740 934 1924
rect 870 -336 934 1740
rect 978 458 1158 1970
rect 1692 1658 1872 2200
rect 1692 1606 1698 1658
rect 1866 1606 1872 1658
rect 1692 1600 1872 1606
rect 978 406 984 458
rect 1152 406 1158 458
rect 978 400 1158 406
rect 2406 6 2412 58
rect 2580 6 2586 58
rect 2406 0 2586 6
rect 2932 6 2938 58
rect 3106 6 3112 58
rect 2932 0 3112 6
rect 870 -342 970 -336
rect 870 -502 910 -342
rect 964 -502 970 -342
rect 870 -508 970 -502
rect 1148 -340 1704 -322
rect 1148 -502 1154 -340
rect 1214 -342 1704 -340
rect 1214 -502 1636 -342
rect 1696 -502 1704 -342
rect 1148 -522 1704 -502
rect 1860 -340 2654 -322
rect 1860 -342 2582 -340
rect 1860 -502 1868 -342
rect 1928 -500 2582 -342
rect 2642 -500 2654 -340
rect 1928 -502 2654 -500
rect 1860 -522 2654 -502
rect 3122 -340 3186 -334
rect 3122 -500 3128 -340
rect 3180 -500 3186 -340
rect 2332 -582 2396 -576
rect 2332 -742 2338 -582
rect 2390 -742 2396 -582
rect 2332 -1068 2396 -742
rect 2332 -1252 2338 -1068
rect 2390 -1252 2396 -1068
rect 2332 -1260 2396 -1252
rect 3122 -1296 3186 -500
rect 3122 -1480 3128 -1296
rect 3180 -1480 3186 -1296
rect 3122 -1488 3186 -1480
use sky130_fd_pr__pfet_g5v0d10v5_243UAW  sky130_fd_pr__pfet_g5v0d10v5_243UAW_0
timestamp 1717438773
transform 1 0 1782 0 1 359
box -358 -1497 358 1497
use sky130_fd_pr__pfet_g5v0d10v5_FGF6VM  sky130_fd_pr__pfet_g5v0d10v5_FGF6VM_0
timestamp 1717438773
transform 1 0 1068 0 1 -241
box -358 -897 358 897
use sky130_fd_pr__pfet_g5v0d10v5_FGR8VM  sky130_fd_pr__pfet_g5v0d10v5_FGR8VM_0
timestamp 1717417325
transform 1 0 3022 0 1 -441
box -358 -697 358 697
use sky130_fd_pr__pfet_g5v0d10v5_FGR8VM  sky130_fd_pr__pfet_g5v0d10v5_FGR8VM_1
timestamp 1717417325
transform 1 0 2496 0 1 -441
box -358 -697 358 697
<< labels >>
flabel metal1 s 710 1830 724 1834 3 FreeSans 800 0 0 0 avdd
port 0 e
flabel metal1 s 710 -1172 710 -1172 3 FreeSans 800 0 0 0 iout
port 6 e
flabel metal1 s 710 -1386 710 -1386 3 FreeSans 800 0 0 0 iout_n
port 5 e
flabel metal1 s 710 2280 710 2280 3 FreeSans 800 0 0 0 pcbias
port 2 e
flabel metal1 s 710 2072 710 2072 3 FreeSans 800 0 0 0 pbias
port 1 e
flabel metal1 s 2494 22 2494 22 0 FreeSans 800 0 0 0 sw_b
port 3 nsew
flabel metal1 s 3020 20 3020 20 0 FreeSans 800 0 0 0 sw_bn
port 4 nsew
<< end >>
