magic
tech sky130A
magscale 1 2
timestamp 1717434370
<< pwell >>
rect 149 -2436 805 -1930
rect 1239 -2272 1811 -2088
rect 149 -2472 806 -2436
rect 149 -2530 805 -2472
<< viali >>
rect 949 -2483 1317 -2448
<< metal1 >>
rect 149 -430 2514 -422
rect 149 -616 1496 -430
rect 1548 -616 2514 -430
rect 149 -622 2514 -616
rect 149 -658 2514 -650
rect 149 -844 2294 -658
rect 2348 -844 2514 -658
rect 149 -850 2514 -844
rect 307 -1500 371 -1488
rect 307 -1660 313 -1500
rect 365 -1660 371 -1500
rect 307 -1672 371 -1660
rect 583 -1672 1027 -1072
rect 1490 -1084 1553 -1072
rect 1490 -1244 1495 -1084
rect 1547 -1244 1553 -1084
rect 1490 -1256 1553 -1244
rect 382 -1710 573 -1704
rect 382 -1763 416 -1710
rect 536 -1763 573 -1710
rect 382 -1769 573 -1763
rect 1765 -2088 2079 -1072
rect 2291 -1084 2354 -1072
rect 2291 -1244 2297 -1084
rect 2349 -1244 2354 -1084
rect 2291 -1256 2354 -1244
rect 1239 -2100 1297 -2088
rect 1239 -2260 1245 -2100
rect 1239 -2272 1297 -2260
rect 1747 -2100 2079 -2088
rect 1747 -2260 1753 -2100
rect 1805 -2260 2079 -2100
rect 1747 -2271 2079 -2260
rect 1765 -2272 2079 -2271
rect 1036 -2357 1073 -2304
rect 1193 -2357 1229 -2304
rect 1036 -2363 1229 -2357
rect 149 -2448 2514 -2436
rect 149 -2470 949 -2448
rect 149 -2630 314 -2470
rect 366 -2483 949 -2470
rect 1317 -2483 2514 -2448
rect 366 -2630 2514 -2483
rect 149 -2636 2514 -2630
rect 149 -2805 2514 -2664
rect 149 -2858 417 -2805
rect 537 -2858 2514 -2805
rect 149 -2864 2514 -2858
rect 149 -3033 2514 -2892
rect 149 -3086 1074 -3033
rect 1194 -3086 2514 -3033
rect 149 -3092 2514 -3086
<< via1 >>
rect 1496 -616 1548 -430
rect 2294 -844 2348 -658
rect 313 -1660 365 -1500
rect 1495 -1244 1547 -1084
rect 416 -1763 536 -1710
rect 2297 -1244 2349 -1084
rect 1245 -2260 1297 -2100
rect 1753 -2260 1805 -2100
rect 1073 -2357 1193 -2304
rect 314 -2630 366 -2470
rect 417 -2858 537 -2805
rect 1074 -3086 1194 -3033
<< metal2 >>
rect 1490 -430 1553 -423
rect 1490 -616 1496 -430
rect 1548 -616 1553 -430
rect 1490 -1084 1553 -616
rect 1490 -1244 1495 -1084
rect 1547 -1244 1553 -1084
rect 1490 -1256 1553 -1244
rect 2291 -658 2354 -650
rect 2291 -844 2294 -658
rect 2348 -844 2354 -658
rect 2291 -1084 2354 -844
rect 2291 -1244 2297 -1084
rect 2349 -1244 2354 -1084
rect 2291 -1256 2354 -1244
rect 307 -1500 371 -1488
rect 307 -1660 313 -1500
rect 365 -1660 371 -1500
rect 307 -2470 371 -1660
rect 307 -2630 314 -2470
rect 366 -2630 371 -2470
rect 410 -1710 542 -1703
rect 410 -1763 416 -1710
rect 536 -1763 542 -1710
rect 410 -2436 542 -1763
rect 1239 -2100 1811 -2088
rect 1239 -2260 1245 -2100
rect 1297 -2260 1753 -2100
rect 1805 -2260 1811 -2100
rect 1239 -2270 1811 -2260
rect 1067 -2304 1199 -2298
rect 1067 -2357 1073 -2304
rect 1193 -2357 1199 -2304
rect 410 -2494 543 -2436
rect 307 -2636 371 -2630
rect 411 -2805 543 -2494
rect 411 -2858 417 -2805
rect 537 -2858 543 -2805
rect 411 -2864 543 -2858
rect 1067 -3033 1199 -2357
rect 1067 -3086 1074 -3033
rect 1194 -3086 1199 -3033
rect 1067 -3092 1199 -3086
use sky130_fd_pr__nfet_g5v0d10v5_BHMQGH  sky130_fd_pr__nfet_g5v0d10v5_BHMQGH_0
timestamp 1717401419
transform 1 0 1133 0 1 -1672
box -328 -858 328 858
use sky130_fd_pr__nfet_g5v0d10v5_D8TNYB  sky130_fd_pr__nfet_g5v0d10v5_D8TNYB_0
timestamp 1717401419
transform 1 0 477 0 1 -1372
box -328 -558 328 558
use sky130_fd_pr__nfet_g5v0d10v5_BHMQGH  XM1
timestamp 1717401419
transform 1 0 1659 0 1 -1672
box -328 -858 328 858
use sky130_fd_pr__nfet_g5v0d10v5_BHMQGH  XM2
timestamp 1717401419
transform 1 0 2185 0 1 -1672
box -328 -858 328 858
<< labels >>
flabel metal1 s 2184 -2328 2184 -2328 0 FreeSans 800 0 0 0 swn
port 7 nsew
flabel metal1 s 1658 -2328 1658 -2328 0 FreeSans 800 0 0 0 sw
port 3 nsew
flabel metal1 s 150 -2552 150 -2552 3 FreeSans 800 0 0 0 avss
port 6 e
flabel metal1 s 150 -2768 150 -2768 3 FreeSans 800 0 0 0 nbias
port 5 e
flabel metal1 s 150 -3006 150 -3006 3 FreeSans 800 0 0 0 ncbias
port 4 e
flabel metal1 s 150 -522 150 -522 3 FreeSans 800 0 0 0 iout
port 0 e
flabel metal1 s 150 -758 150 -758 3 FreeSans 800 0 0 0 ioutn
port 1 e
<< end >>
