magic
tech sky130A
magscale 1 2
timestamp 1717439915
<< metal1 >>
rect 120819 -438 121020 -430
rect 120819 -622 120838 -438
rect 121008 -622 121020 -438
rect 120819 -630 121020 -622
rect 121276 -438 121476 -430
rect 121276 -622 121290 -438
rect 121460 -622 121476 -438
rect 120332 -1122 121020 -1114
rect 120332 -1306 120838 -1122
rect 121008 -1306 121020 -1122
rect 120332 -1314 121020 -1306
rect 120986 -2270 121020 -2262
rect 121008 -2454 121020 -2270
rect 120986 -2462 121020 -2454
rect 120986 -2498 121020 -2490
rect 121008 -2682 121020 -2498
rect 120986 -2690 121020 -2682
rect 120986 -2726 121020 -2718
rect 121008 -2912 121020 -2726
rect 120986 -2918 121020 -2912
rect 120819 -2954 121020 -2946
rect 120819 -3140 120838 -2954
rect 121008 -3140 121020 -2954
rect 120819 -3146 121020 -3140
rect 121048 -2954 121248 -2946
rect 121048 -3140 121062 -2954
rect 121232 -3140 121248 -2954
rect 120442 -8644 121020 -8636
rect 120442 -8828 120840 -8644
rect 121010 -8828 121020 -8644
rect 120442 -8836 121020 -8828
rect 121000 -10474 121020 -10468
rect 121010 -10658 121020 -10474
rect 121000 -10668 121020 -10658
rect 121048 -10474 121248 -3140
rect 121276 -7960 121476 -622
rect 121276 -8144 121292 -7960
rect 121462 -8144 121476 -7960
rect 121276 -8152 121476 -8144
rect 121504 -666 121704 -658
rect 121504 -850 121520 -666
rect 121690 -850 121704 -666
rect 121504 -8188 121704 -850
rect 121504 -8372 121518 -8188
rect 121688 -8372 121704 -8188
rect 121504 -8380 121704 -8372
rect 121732 -892 121932 -886
rect 121732 -1076 121748 -892
rect 121918 -1076 121932 -892
rect 121732 -8414 121932 -1076
rect 121732 -8598 121746 -8414
rect 121916 -8598 121932 -8414
rect 121732 -8604 121932 -8598
rect 121960 -1124 122160 -1114
rect 121960 -1308 121976 -1124
rect 122146 -1308 122160 -1124
rect 121960 -8642 122160 -1308
rect 121960 -8826 121976 -8642
rect 122146 -8826 122160 -8642
rect 121960 -8836 122160 -8826
rect 122188 -2270 122388 -2262
rect 122188 -2454 122204 -2270
rect 122374 -2454 122388 -2270
rect 122188 -9792 122388 -2454
rect 122188 -9976 122204 -9792
rect 122374 -9976 122388 -9792
rect 122188 -9984 122388 -9976
rect 122416 -2496 122616 -2490
rect 122416 -2680 122432 -2496
rect 122602 -2680 122616 -2496
rect 122416 -10020 122616 -2680
rect 122416 -10204 122430 -10020
rect 122600 -10204 122616 -10020
rect 122416 -10212 122616 -10204
rect 122644 -2724 122844 -2718
rect 122644 -2908 122660 -2724
rect 122830 -2908 122844 -2724
rect 122644 -10248 122844 -2908
rect 122644 -10432 122660 -10248
rect 122830 -10432 122844 -10248
rect 122644 -10440 122844 -10432
rect 121048 -10658 121062 -10474
rect 121232 -10658 121248 -10474
rect 121048 -10668 121248 -10658
<< via1 >>
rect 120838 -622 121008 -438
rect 121290 -622 121460 -438
rect 120838 -850 121008 -666
rect 120838 -1078 121008 -894
rect 120838 -1306 121008 -1122
rect 120838 -2454 121008 -2270
rect 120838 -2682 121008 -2498
rect 120838 -2912 121008 -2726
rect 120838 -3140 121008 -2954
rect 121062 -3140 121232 -2954
rect 120840 -8144 121010 -7960
rect 120840 -8372 121010 -8188
rect 120840 -8598 121010 -8414
rect 120840 -8828 121010 -8644
rect 120840 -9976 121010 -9792
rect 120840 -10204 121010 -10020
rect 120840 -10432 121010 -10248
rect 120840 -10658 121010 -10474
rect 121292 -8144 121462 -7960
rect 121520 -850 121690 -666
rect 121518 -8372 121688 -8188
rect 121748 -1076 121918 -892
rect 121746 -8598 121916 -8414
rect 121976 -1308 122146 -1124
rect 121976 -8826 122146 -8642
rect 122204 -2454 122374 -2270
rect 122204 -9976 122374 -9792
rect 122432 -2680 122602 -2496
rect 122430 -10204 122600 -10020
rect 122660 -2908 122830 -2724
rect 122660 -10432 122830 -10248
rect 121062 -10658 121232 -10474
<< metal2 >>
rect 120832 -438 121476 -430
rect 120832 -622 120838 -438
rect 121008 -622 121290 -438
rect 121460 -622 121476 -438
rect 120832 -630 121476 -622
rect 120832 -666 121704 -658
rect 120832 -850 120838 -666
rect 121008 -850 121520 -666
rect 121690 -850 121704 -666
rect 120832 -858 121704 -850
rect 120832 -892 121932 -886
rect 120832 -894 121748 -892
rect 120832 -1078 120838 -894
rect 121008 -1076 121748 -894
rect 121918 -1076 121932 -892
rect 121008 -1078 121932 -1076
rect 120832 -1086 121932 -1078
rect 120832 -1122 122160 -1114
rect 120832 -1306 120838 -1122
rect 121008 -1124 122160 -1122
rect 121008 -1306 121976 -1124
rect 120832 -1308 121976 -1306
rect 122146 -1308 122160 -1124
rect 120832 -1314 122160 -1308
rect 120832 -2270 122388 -2262
rect 120832 -2454 120838 -2270
rect 121008 -2454 122204 -2270
rect 122374 -2454 122388 -2270
rect 120832 -2462 122388 -2454
rect 120832 -2496 122616 -2490
rect 120832 -2498 122432 -2496
rect 120832 -2682 120838 -2498
rect 121008 -2680 122432 -2498
rect 122602 -2680 122616 -2496
rect 121008 -2682 122616 -2680
rect 120832 -2690 122616 -2682
rect 120832 -2724 122844 -2718
rect 120832 -2726 122660 -2724
rect 120832 -2912 120838 -2726
rect 121008 -2908 122660 -2726
rect 122830 -2908 122844 -2724
rect 121008 -2912 122844 -2908
rect 120832 -2918 122844 -2912
rect 120818 -2954 121248 -2946
rect 120818 -3140 120838 -2954
rect 121008 -3140 121062 -2954
rect 121232 -3140 121248 -2954
rect 120818 -3146 121248 -3140
rect 120834 -7960 121476 -7952
rect 120834 -8144 120840 -7960
rect 121010 -8144 121292 -7960
rect 121462 -8144 121476 -7960
rect 120834 -8152 121476 -8144
rect 120834 -8188 121704 -8180
rect 120834 -8372 120840 -8188
rect 121010 -8372 121518 -8188
rect 121688 -8372 121704 -8188
rect 120834 -8380 121704 -8372
rect 120834 -8414 121932 -8408
rect 120834 -8598 120840 -8414
rect 121010 -8598 121746 -8414
rect 121916 -8598 121932 -8414
rect 120834 -8608 121932 -8598
rect 120834 -8642 122160 -8636
rect 120834 -8644 121976 -8642
rect 120834 -8828 120840 -8644
rect 121010 -8826 121976 -8644
rect 122146 -8826 122160 -8642
rect 121010 -8828 122160 -8826
rect 120834 -8836 122160 -8828
rect 120834 -9792 122388 -9784
rect 120834 -9976 120840 -9792
rect 121010 -9976 122204 -9792
rect 122374 -9976 122388 -9792
rect 120834 -9984 122388 -9976
rect 120834 -10020 122616 -10012
rect 120834 -10204 120840 -10020
rect 121010 -10204 122430 -10020
rect 122600 -10204 122616 -10020
rect 120834 -10212 122616 -10204
rect 120834 -10248 122844 -10240
rect 120834 -10432 120840 -10248
rect 121010 -10432 122660 -10248
rect 122830 -10432 122844 -10248
rect 120834 -10440 122844 -10432
rect 120834 -10474 121248 -10468
rect 120834 -10658 120840 -10474
rect 121010 -10658 121062 -10474
rect 121232 -10658 121248 -10474
rect 120834 -10668 121248 -10658
use icell32scs  x1
timestamp 1717438951
transform 1 0 0 0 1 0
box 4862 -5160 121061 2790
use icell32scs  x2
timestamp 1717438951
transform -1 0 125884 0 1 -7522
box 4862 -5160 121061 2790
<< end >>
