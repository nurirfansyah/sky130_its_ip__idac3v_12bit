magic
tech sky130A
magscale 1 2
timestamp 1717438951
<< nwell >>
rect 1168 -1632 1216 -1630
rect 1168 -1780 1202 -1632
rect 1820 -1772 1980 -1636
rect 2972 -1922 3030 -1866
rect 2138 -2058 2210 -1986
rect 2366 -1992 2424 -1942
<< pwell >>
rect 1654 -2182 1726 -2180
rect 1168 -2512 4798 -2182
rect 1654 -3532 1944 -3466
<< locali >>
rect 2378 -2102 2412 -1982
rect 2984 -2104 3018 -1912
<< viali >>
rect 2984 -1912 3018 -1878
rect 2378 -1982 2412 -1948
rect 1288 -2144 1322 -2110
rect 2154 -2136 2188 -2102
rect 2258 -2136 2292 -2102
rect 2378 -2136 2412 -2102
rect 2496 -2136 2530 -2102
rect 2708 -2152 2742 -2118
rect 2864 -2148 2898 -2114
rect 2984 -2138 3018 -2104
rect 3114 -2138 3148 -2104
rect 3288 -2136 3322 -2102
rect 3542 -2136 3576 -2102
rect 3900 -2146 3934 -2112
rect 4128 -2146 4162 -2112
rect 4328 -2164 4362 -2130
rect 4710 -2152 4744 -2118
rect 1840 -2228 1876 -2194
rect 3284 -2246 3318 -2212
rect 3810 -2226 3844 -2192
rect 1480 -2300 1514 -2266
<< metal1 >>
rect 3590 2522 4798 2532
rect 3590 2340 3972 2522
rect 4140 2340 4798 2522
rect 3590 2332 4798 2340
rect 3374 2294 4798 2304
rect 3374 2112 4254 2294
rect 4422 2112 4798 2294
rect 3374 2104 4798 2112
rect 1956 348 2146 354
rect 3792 348 3864 354
rect 1956 276 1962 348
rect 2140 276 2146 348
rect 3180 276 3186 348
rect 3258 276 3792 348
rect 1956 270 2146 276
rect 3792 270 3864 276
rect 1430 236 1620 242
rect 1430 164 1436 236
rect 1614 164 1620 236
rect 1430 158 1620 164
rect 3194 -888 4798 -688
rect 3614 -1114 3636 -916
rect 3638 -1114 4798 -916
rect 3614 -1116 4798 -1114
rect 2550 -1336 2602 -1152
rect 3638 -1344 4798 -1144
rect 1522 -1380 4442 -1372
rect 1522 -1564 2148 -1380
rect 2200 -1564 4442 -1380
rect 1522 -1572 4442 -1564
rect 1168 -1636 4798 -1630
rect 1168 -1772 1820 -1636
rect 1980 -1772 4798 -1636
rect 1168 -1780 4798 -1772
rect 1930 -1864 2002 -1858
rect 1930 -1872 1936 -1864
rect 1283 -1914 1936 -1872
rect 1283 -2104 1325 -1914
rect 1930 -1924 1936 -1914
rect 1996 -1872 2002 -1864
rect 2972 -1872 3030 -1866
rect 1996 -1878 3030 -1872
rect 1996 -1912 2984 -1878
rect 3018 -1880 3030 -1878
rect 3018 -1912 4366 -1880
rect 1996 -1914 4366 -1912
rect 1996 -1924 2002 -1914
rect 2972 -1922 4366 -1914
rect 1930 -1930 2002 -1924
rect 2366 -1948 2424 -1942
rect 2366 -1982 2378 -1948
rect 2412 -1950 2424 -1948
rect 2412 -1982 4166 -1950
rect 2138 -1992 2210 -1986
rect 2366 -1992 4166 -1982
rect 2138 -2052 2144 -1992
rect 2204 -2020 2210 -1992
rect 2204 -2052 3938 -2020
rect 2138 -2058 3938 -2052
rect 2150 -2062 3938 -2058
rect 2150 -2090 2192 -2062
rect 2142 -2102 2200 -2090
rect 1276 -2110 1334 -2104
rect 1276 -2144 1288 -2110
rect 1322 -2144 1334 -2110
rect 1276 -2156 1334 -2144
rect 2142 -2136 2154 -2102
rect 2188 -2136 2200 -2102
rect 2142 -2148 2200 -2136
rect 2246 -2098 2298 -2090
rect 2372 -2098 2418 -2096
rect 2490 -2098 2542 -2090
rect 2246 -2102 2542 -2098
rect 2246 -2136 2258 -2102
rect 2292 -2136 2378 -2102
rect 2412 -2136 2496 -2102
rect 2530 -2136 2542 -2102
rect 2246 -2140 2542 -2136
rect 2246 -2148 2298 -2140
rect 2372 -2142 2418 -2140
rect 2490 -2148 2542 -2140
rect 1654 -2240 1660 -2180
rect 1720 -2182 1726 -2180
rect 1720 -2194 1888 -2182
rect 1720 -2228 1840 -2194
rect 1876 -2228 1888 -2194
rect 1720 -2240 1888 -2228
rect 1472 -2266 1526 -2254
rect 1472 -2300 1480 -2266
rect 1514 -2274 1526 -2266
rect 2150 -2274 2192 -2148
rect 2690 -2166 2696 -2106
rect 2756 -2166 2762 -2106
rect 2854 -2114 2906 -2100
rect 2854 -2148 2864 -2114
rect 2898 -2148 2906 -2114
rect 2854 -2158 2906 -2148
rect 2954 -2104 3170 -2090
rect 2954 -2138 2984 -2104
rect 3018 -2138 3114 -2104
rect 3148 -2138 3170 -2104
rect 2954 -2150 3170 -2138
rect 3278 -2098 3330 -2090
rect 3536 -2098 3588 -2090
rect 3278 -2102 3588 -2098
rect 3896 -2100 3938 -2062
rect 3278 -2136 3288 -2102
rect 3322 -2136 3542 -2102
rect 3576 -2136 3588 -2102
rect 3278 -2140 3588 -2136
rect 3278 -2148 3330 -2140
rect 3536 -2148 3588 -2140
rect 3890 -2112 3942 -2100
rect 4124 -2106 4166 -1992
rect 3890 -2146 3900 -2112
rect 3934 -2146 3942 -2112
rect 3890 -2158 3942 -2146
rect 4116 -2112 4174 -2106
rect 4116 -2146 4128 -2112
rect 4162 -2146 4174 -2112
rect 4324 -2124 4366 -1922
rect 4702 -2106 4762 -2100
rect 4116 -2158 4174 -2146
rect 4316 -2130 4374 -2124
rect 2858 -2208 2900 -2158
rect 4316 -2164 4328 -2130
rect 4362 -2164 4374 -2130
rect 3798 -2180 3858 -2174
rect 4316 -2176 4374 -2164
rect 4702 -2172 4762 -2166
rect 3278 -2208 3330 -2200
rect 2858 -2212 3330 -2208
rect 2858 -2246 3284 -2212
rect 3318 -2246 3330 -2212
rect 3798 -2246 3858 -2240
rect 2858 -2250 3330 -2246
rect 3278 -2258 3330 -2250
rect 1514 -2300 2192 -2274
rect 1472 -2316 2192 -2300
rect 1168 -2350 4798 -2344
rect 1168 -2486 3618 -2350
rect 3778 -2486 4798 -2350
rect 1168 -2492 4798 -2486
rect 1168 -2528 4798 -2520
rect 1168 -2712 1940 -2528
rect 1992 -2712 4798 -2528
rect 1168 -2720 4798 -2712
rect 3333 -2948 4798 -2748
rect 1490 -3096 1562 -3024
rect 1664 -3104 1716 -2984
rect 1654 -3176 1726 -3104
rect 3333 -3176 4798 -2976
rect 2978 -3210 4798 -3204
rect 2978 -3398 3618 -3210
rect 3778 -3398 4798 -3210
rect 2978 -3404 4798 -3398
rect 1932 -3472 2112 -3466
rect 1932 -3526 1938 -3472
rect 2106 -3526 2112 -3472
rect 1932 -3532 2112 -3526
rect 1448 -4400 1540 -4384
rect 1448 -4460 1464 -4400
rect 1524 -4460 1540 -4400
rect 1448 -4840 1540 -4460
rect 3842 -4394 3914 -4388
rect 3914 -4466 4464 -4394
rect 4536 -4466 4542 -4394
rect 3842 -4472 3914 -4466
rect 3242 -4998 4798 -4990
rect 3242 -5180 3972 -4998
rect 4140 -5180 4798 -4998
rect 3242 -5190 4798 -5180
rect 3222 -5228 4798 -5218
rect 3222 -5410 4254 -5228
rect 4422 -5410 4798 -5228
rect 3222 -5418 4798 -5410
<< via1 >>
rect 3972 2340 4140 2522
rect 4254 2112 4422 2294
rect 1962 276 2140 348
rect 3186 276 3258 348
rect 3792 276 3864 348
rect 1436 164 1614 236
rect 1818 -880 1984 -698
rect 2148 -1564 2200 -1380
rect 1820 -1772 1980 -1636
rect 1936 -1924 1996 -1864
rect 2144 -2052 2204 -1992
rect 1660 -2240 1720 -2180
rect 2696 -2118 2756 -2106
rect 2696 -2152 2708 -2118
rect 2708 -2152 2742 -2118
rect 2742 -2152 2756 -2118
rect 2696 -2166 2756 -2152
rect 4702 -2118 4762 -2106
rect 4702 -2152 4710 -2118
rect 4710 -2152 4744 -2118
rect 4744 -2152 4762 -2118
rect 4702 -2166 4762 -2152
rect 3798 -2192 3858 -2180
rect 3798 -2226 3810 -2192
rect 3810 -2226 3844 -2192
rect 3844 -2226 3858 -2192
rect 3798 -2240 3858 -2226
rect 3618 -2486 3778 -2350
rect 1940 -2712 1992 -2528
rect 3618 -3398 3778 -3210
rect 1938 -3526 2106 -3472
rect 1464 -4460 1524 -4400
rect 3842 -4466 3914 -4394
rect 4464 -4466 4536 -4394
rect 3972 -5180 4140 -4998
rect 4254 -5410 4422 -5228
<< metal2 >>
rect 3966 2522 4146 2532
rect 3966 2340 3972 2522
rect 4140 2340 4146 2522
rect 1436 242 1614 1044
rect 1962 354 2140 1044
rect 1956 348 2146 354
rect 3186 348 3258 354
rect 1956 276 1962 348
rect 2140 276 3186 348
rect 3786 276 3792 348
rect 3864 276 3870 348
rect 1956 270 2146 276
rect 3186 270 3258 276
rect 1430 236 1620 242
rect 1430 164 1436 236
rect 1614 164 2378 236
rect 1430 158 1620 164
rect 1810 -698 1990 -688
rect 1810 -880 1818 -698
rect 1984 -880 1990 -698
rect 1810 -1636 1990 -880
rect 1810 -1772 1820 -1636
rect 1980 -1772 1990 -1636
rect 1810 -1780 1990 -1772
rect 2138 -1380 2210 -1372
rect 2138 -1564 2148 -1380
rect 2200 -1564 2210 -1380
rect 1930 -1864 2002 -1858
rect 1930 -1924 1936 -1864
rect 1996 -1924 2002 -1864
rect 1654 -2180 1726 -2174
rect 1654 -2240 1660 -2180
rect 1720 -2240 1726 -2180
rect 1654 -3466 1726 -2240
rect 1930 -2528 2002 -1924
rect 2138 -1992 2210 -1564
rect 2138 -2052 2144 -1992
rect 2204 -2052 2210 -1992
rect 2138 -2058 2210 -2052
rect 2306 -2100 2378 164
rect 2306 -2106 2762 -2100
rect 2306 -2166 2696 -2106
rect 2756 -2166 2762 -2106
rect 2306 -2172 2762 -2166
rect 3792 -2180 3864 276
rect 3792 -2240 3798 -2180
rect 3858 -2240 3864 -2180
rect 3792 -2246 3864 -2240
rect 1930 -2712 1940 -2528
rect 1992 -2712 2002 -2528
rect 1930 -2720 2002 -2712
rect 3612 -2350 3784 -2344
rect 3612 -2486 3618 -2350
rect 3778 -2486 3784 -2350
rect 3612 -3210 3784 -2486
rect 3612 -3398 3618 -3210
rect 3778 -3398 3784 -3210
rect 3612 -3404 3784 -3398
rect 1654 -3472 2112 -3466
rect 1654 -3526 1938 -3472
rect 2106 -3526 2112 -3472
rect 1654 -3532 2112 -3526
rect 1458 -4400 3842 -4394
rect 1458 -4460 1464 -4400
rect 1524 -4460 3842 -4400
rect 1458 -4466 3842 -4460
rect 3914 -4466 3920 -4394
rect 3966 -4998 4146 2340
rect 3966 -5180 3972 -4998
rect 4140 -5180 4146 -4998
rect 3966 -5190 4146 -5180
rect 4248 2294 4428 2304
rect 4248 2112 4254 2294
rect 4422 2112 4428 2294
rect 4248 -5228 4428 2112
rect 4464 -2106 4768 -2100
rect 4464 -2166 4702 -2106
rect 4762 -2166 4768 -2106
rect 4464 -4394 4536 -2166
rect 4464 -4472 4536 -4466
rect 4248 -5410 4254 -5228
rect 4422 -5410 4428 -5228
rect 4248 -5418 4428 -5410
use pcell1scs  x1
timestamp 1717438773
transform -1 0 4548 0 -1 1044
box 710 -1488 3380 2388
use ncell1scs  x2
timestamp 1717434370
transform -1 0 3682 0 -1 -5840
box 149 -3092 2514 -422
use sky130_fd_sc_hvl__nand2_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 3490 0 1 -2469
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 3070 0 1 -2469
box -66 -43 354 897
use sky130_fd_sc_hvl__and2_1  x5 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 1234 0 1 -2469
box -66 -43 738 897
use sky130_fd_sc_hvl__inv_1  x6
timestamp 1710522493
transform 1 0 2038 0 1 -2469
box -66 -43 354 897
use sky130_fd_sc_hvl__nand2_1  x7
timestamp 1710522493
transform 1 0 2458 0 1 -2469
box -66 -43 546 897
use sky130_fd_sc_hvl__and2_1  x8
timestamp 1710522493
transform 1 0 4102 0 1 -2469
box -66 -43 738 897
<< labels >>
flabel metal1 s 1168 -1016 1168 -1016 3 FreeSans 800 0 0 0 pbias
port 2 e
flabel metal1 s 1168 -1256 1168 -1256 3 FreeSans 800 0 0 0 pcbias
port 5 e
flabel metal1 s 1168 -2636 1168 -2636 3 FreeSans 800 0 0 0 idir_sel
port 6 e
flabel metal1 s 1168 -2860 1168 -2860 3 FreeSans 800 0 0 0 ncbias
port 7 e
flabel metal1 s 1168 -3080 1168 -3080 3 FreeSans 800 0 0 0 nbias
port 8 e
flabel metal1 s 1168 -796 1168 -796 3 FreeSans 800 0 0 0 avdd
port 1 e
flabel metal1 s 1168 2426 1168 2426 3 FreeSans 800 0 0 0 ioutn
port 3 e
flabel metal1 s 1168 -3310 1168 -3310 3 FreeSans 800 0 0 0 avss
port 9 e
flabel metal1 s 1564 -1474 1564 -1474 3 FreeSans 800 0 0 0 sw
port 4 e
flabel metal1 s 1168 2204 1168 2204 3 FreeSans 800 0 0 0 iout
port 0 e
<< end >>
