magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
rect 0 -8800 200 -8600
rect 0 -9200 200 -9000
rect 0 -9600 200 -9400
rect 0 -10000 200 -9800
use sky130_fd_sc_hvl__and3_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 738 0 1 -10043
box -66 -43 834 897
use sky130_fd_sc_hvl__or2_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 2310 0 1 -10129
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x3
timestamp 1710522493
transform 1 0 3048 0 1 -10172
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1710522493
transform 1 0 3882 0 1 -10215
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x5
timestamp 1710522493
transform 1 0 0 0 1 -10000
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x6
timestamp 1710522493
transform 1 0 4620 0 1 -10258
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x7
timestamp 1710522493
transform 1 0 5358 0 1 -10301
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x8
timestamp 1710522493
transform 1 0 6192 0 1 -10344
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x9
timestamp 1710522493
transform 1 0 6930 0 1 -10387
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x10
timestamp 1710522493
transform 1 0 7668 0 1 -10430
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x11
timestamp 1710522493
transform 1 0 8502 0 1 -10473
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x12
timestamp 1710522493
transform 1 0 9240 0 1 -10516
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x13
timestamp 1710522493
transform 1 0 9978 0 1 -10559
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x14
timestamp 1710522493
transform 1 0 10812 0 1 -10602
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x15
timestamp 1710522493
transform 1 0 11550 0 1 -10645
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x16
timestamp 1710522493
transform 1 0 12288 0 1 -10688
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x17
timestamp 1710522493
transform 1 0 13122 0 1 -10731
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x18
timestamp 1710522493
transform 1 0 13860 0 1 -10774
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x19
timestamp 1710522493
transform 1 0 14598 0 1 -10817
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x20
timestamp 1710522493
transform 1 0 15432 0 1 -10860
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x21
timestamp 1710522493
transform 1 0 16170 0 1 -10903
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x22
timestamp 1710522493
transform 1 0 16908 0 1 -10946
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x23
timestamp 1710522493
transform 1 0 17742 0 1 -10989
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x24
timestamp 1710522493
transform 1 0 18480 0 1 -11032
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x25
timestamp 1710522493
transform 1 0 19218 0 1 -11075
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x26
timestamp 1710522493
transform 1 0 20052 0 1 -11118
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x27
timestamp 1710522493
transform 1 0 20790 0 1 -11161
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x28
timestamp 1710522493
transform 1 0 21528 0 1 -11204
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x29
timestamp 1710522493
transform 1 0 22362 0 1 -11247
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x30
timestamp 1710522493
transform 1 0 23100 0 1 -11290
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x31
timestamp 1710522493
transform 1 0 23838 0 1 -11333
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x32
timestamp 1710522493
transform 1 0 1572 0 1 -10086
box -66 -43 738 897
use sky130_fd_sc_hvl__and2_1  x33
timestamp 1710522493
transform 1 0 24672 0 1 -11376
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x34
timestamp 1710522493
transform 1 0 25410 0 1 -11419
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x35
timestamp 1710522493
transform 1 0 26148 0 1 -11462
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x36
timestamp 1710522493
transform 1 0 26982 0 1 -11505
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x41
timestamp 1710522493
transform 1 0 27720 0 1 -11548
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x42
timestamp 1710522493
transform 1 0 28554 0 1 -11591
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x43
timestamp 1710522493
transform 1 0 29292 0 1 -11634
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x44
timestamp 1710522493
transform 1 0 30030 0 1 -11677
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x45
timestamp 1710522493
transform 1 0 30864 0 1 -11720
box -66 -43 738 897
use sky130_fd_sc_hvl__or2_1  x46
timestamp 1710522493
transform 1 0 31602 0 1 -11763
box -66 -43 738 897
use sky130_fd_sc_hvl__and3_1  x47
timestamp 1710522493
transform 1 0 32340 0 1 -11806
box -66 -43 834 897
use sky130_fd_sc_hvl__and2_1  x48
timestamp 1710522493
transform 1 0 33174 0 1 -11849
box -66 -43 738 897
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avss
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 din0
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 t0
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 din1
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 t1
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 din2
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 t2
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 t3
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 din3
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 t4
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 t5
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 t6
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 t7
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 din0_n
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 din1_n
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 t8
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 t9
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 din2_n
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 din3_n
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 t10
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 256 0 0 0 t11
port 21 nsew
flabel metal1 0 -8800 200 -8600 0 FreeSans 256 0 0 0 t12
port 22 nsew
flabel metal1 0 -9200 200 -9000 0 FreeSans 256 0 0 0 {}
port 23 nsew
flabel metal1 0 -9600 200 -9400 0 FreeSans 256 0 0 0 t13
port 24 nsew
flabel metal1 0 -10000 200 -9800 0 FreeSans 256 0 0 0 t14
port 25 nsew
<< end >>
