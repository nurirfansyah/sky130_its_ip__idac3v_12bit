magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 217375 -8565 217491 -8499
rect 220719 -8565 220835 -8499
rect 224063 -8565 224179 -8499
rect 227407 -8565 227523 -8499
rect 230751 -8565 230867 -8499
rect 234095 -8565 234211 -8499
rect 237439 -8565 237555 -8499
rect 240783 -8565 240899 -8499
rect 244127 -8565 244243 -8499
rect 247471 -8565 247587 -8499
rect 250815 -8565 250931 -8499
rect 254159 -8565 254275 -8499
rect 257503 -8565 257619 -8499
rect 260847 -8565 260963 -8499
rect 264191 -8565 264307 -8499
rect 267535 -8565 267651 -8499
rect 270879 -8565 270995 -8499
rect 274223 -8565 274339 -8499
rect 277567 -8565 277683 -8499
rect 280911 -8565 281027 -8499
rect 284255 -8565 284371 -8499
rect 287599 -8565 287715 -8499
rect 290943 -8565 291059 -8499
rect 294287 -8565 294403 -8499
rect 297631 -8565 297747 -8499
rect 300975 -8565 301091 -8499
rect 304319 -8565 304435 -8499
rect 307663 -8565 307779 -8499
rect 311007 -8565 311123 -8499
rect 314351 -8565 314467 -8499
rect 317695 -8565 317811 -8499
rect 321039 -8565 321155 -8499
rect 324383 -8565 324499 -8499
rect 327727 -8565 327843 -8499
rect 331071 -8565 331187 -8499
rect 334415 -8565 334531 -8499
rect 337759 -8565 337875 -8499
rect 341103 -8565 341219 -8499
rect 344447 -8565 344563 -8499
rect 347791 -8565 347907 -8499
rect 351135 -8565 351251 -8499
rect 354479 -8565 354595 -8499
rect 357823 -8565 357939 -8499
rect 361167 -8565 361283 -8499
rect 364511 -8565 364627 -8499
rect 367855 -8565 367971 -8499
rect 371199 -8565 371315 -8499
rect 374543 -8565 374659 -8499
rect 377887 -8565 378003 -8499
rect 381231 -8565 381347 -8499
rect 384575 -8565 384691 -8499
rect 387919 -8565 388035 -8499
rect 391263 -8565 391379 -8499
rect 394607 -8565 394723 -8499
rect 397951 -8565 398067 -8499
rect 401295 -8565 401411 -8499
rect 404639 -8565 404755 -8499
rect 407983 -8565 408099 -8499
rect 411327 -8565 411443 -8499
rect 414671 -8565 414787 -8499
rect 418015 -8565 418131 -8499
rect 421359 -8565 421475 -8499
rect 424703 -8565 424819 -8499
rect 217227 -8832 217237 -8819
rect 217161 -8874 217237 -8832
rect 217289 -8874 217491 -8819
rect 217305 -8877 217491 -8874
rect 220835 -8819 221221 -8753
rect 224179 -8819 224565 -8753
rect 227523 -8819 227909 -8753
rect 230867 -8819 231253 -8753
rect 234211 -8819 234597 -8753
rect 237555 -8819 237941 -8753
rect 240899 -8819 241285 -8753
rect 244243 -8819 244629 -8753
rect 247587 -8819 247973 -8753
rect 250931 -8819 251317 -8753
rect 254275 -8819 254661 -8753
rect 257619 -8819 258005 -8753
rect 260963 -8819 261349 -8753
rect 264307 -8819 264693 -8753
rect 267651 -8819 268037 -8753
rect 270995 -8819 271381 -8753
rect 274339 -8819 274725 -8753
rect 277683 -8819 278069 -8753
rect 281027 -8819 281413 -8753
rect 284371 -8819 284757 -8753
rect 287715 -8819 288101 -8753
rect 291059 -8819 291445 -8753
rect 294403 -8819 294789 -8753
rect 297747 -8819 298133 -8753
rect 301091 -8819 301477 -8753
rect 304435 -8819 304821 -8753
rect 307779 -8819 308165 -8753
rect 311123 -8819 311509 -8753
rect 314467 -8819 314853 -8753
rect 317811 -8819 318197 -8753
rect 321155 -8819 321541 -8753
rect 324499 -8819 324885 -8753
rect 327843 -8819 328229 -8753
rect 331187 -8819 331573 -8753
rect 334531 -8819 334917 -8753
rect 337875 -8819 338261 -8753
rect 341219 -8819 341605 -8753
rect 344563 -8819 344949 -8753
rect 347907 -8819 348293 -8753
rect 351251 -8819 351637 -8753
rect 354595 -8819 354981 -8753
rect 357939 -8819 358325 -8753
rect 361283 -8819 361669 -8753
rect 364627 -8819 365013 -8753
rect 367971 -8819 368357 -8753
rect 371315 -8819 371701 -8753
rect 374659 -8819 375045 -8753
rect 378003 -8819 378389 -8753
rect 381347 -8819 381733 -8753
rect 384691 -8819 385077 -8753
rect 388035 -8819 388421 -8753
rect 391379 -8819 391765 -8753
rect 394723 -8819 395109 -8753
rect 398067 -8819 398453 -8753
rect 401411 -8819 401797 -8753
rect 404755 -8819 405141 -8753
rect 408099 -8819 408485 -8753
rect 411443 -8819 411829 -8753
rect 414787 -8819 415173 -8753
rect 418131 -8819 418517 -8753
rect 421475 -8819 421861 -8753
rect 424819 -8819 425205 -8753
rect 220571 -8832 220581 -8819
rect 220505 -8874 220581 -8832
rect 220633 -8874 221221 -8819
rect 223915 -8832 223925 -8819
rect 220505 -8877 221221 -8874
rect 217419 -8993 217619 -8985
rect 217435 -8997 217603 -8993
rect 217361 -9174 217461 -9050
rect 220505 -9114 220649 -8877
rect 220835 -8899 221221 -8877
rect 220759 -8985 221221 -8899
rect 223849 -8874 223925 -8832
rect 223977 -8874 224565 -8819
rect 227259 -8832 227269 -8819
rect 223849 -8877 224565 -8874
rect 220763 -8993 220963 -8985
rect 220779 -8997 220947 -8993
rect 217361 -9228 217363 -9174
rect 220505 -9200 220679 -9114
rect 220705 -9174 220805 -9050
rect 223849 -9114 223993 -8877
rect 224179 -8899 224565 -8877
rect 224103 -8985 224565 -8899
rect 227193 -8874 227269 -8832
rect 227321 -8874 227909 -8819
rect 230603 -8832 230613 -8819
rect 227193 -8877 227909 -8874
rect 224107 -8993 224307 -8985
rect 224123 -8997 224291 -8993
rect 220705 -9228 220707 -9174
rect 223849 -9200 224023 -9114
rect 224049 -9174 224149 -9050
rect 227193 -9114 227337 -8877
rect 227523 -8899 227909 -8877
rect 227447 -8985 227909 -8899
rect 230537 -8874 230613 -8832
rect 230665 -8874 231253 -8819
rect 233947 -8832 233957 -8819
rect 230537 -8877 231253 -8874
rect 227451 -8993 227651 -8985
rect 227467 -8997 227635 -8993
rect 224049 -9228 224051 -9174
rect 227193 -9200 227367 -9114
rect 227393 -9174 227493 -9050
rect 230537 -9114 230681 -8877
rect 230867 -8899 231253 -8877
rect 230791 -8985 231253 -8899
rect 233881 -8874 233957 -8832
rect 234009 -8874 234597 -8819
rect 237291 -8832 237301 -8819
rect 233881 -8877 234597 -8874
rect 230795 -8993 230995 -8985
rect 230811 -8997 230979 -8993
rect 227393 -9228 227395 -9174
rect 230537 -9200 230711 -9114
rect 230737 -9174 230837 -9050
rect 233881 -9114 234025 -8877
rect 234211 -8899 234597 -8877
rect 234135 -8985 234597 -8899
rect 237225 -8874 237301 -8832
rect 237353 -8874 237941 -8819
rect 240635 -8832 240645 -8819
rect 237225 -8877 237941 -8874
rect 234139 -8993 234339 -8985
rect 234155 -8997 234323 -8993
rect 230737 -9228 230739 -9174
rect 233881 -9200 234055 -9114
rect 234081 -9174 234181 -9050
rect 237225 -9114 237369 -8877
rect 237555 -8899 237941 -8877
rect 237479 -8985 237941 -8899
rect 240569 -8874 240645 -8832
rect 240697 -8874 241285 -8819
rect 243979 -8832 243989 -8819
rect 240569 -8877 241285 -8874
rect 237483 -8993 237683 -8985
rect 237499 -8997 237667 -8993
rect 234081 -9228 234083 -9174
rect 237225 -9200 237399 -9114
rect 237425 -9174 237525 -9050
rect 240569 -9114 240713 -8877
rect 240899 -8899 241285 -8877
rect 240823 -8985 241285 -8899
rect 243913 -8874 243989 -8832
rect 244041 -8874 244629 -8819
rect 247323 -8832 247333 -8819
rect 243913 -8877 244629 -8874
rect 240827 -8993 241027 -8985
rect 240843 -8997 241011 -8993
rect 237425 -9228 237427 -9174
rect 240569 -9200 240743 -9114
rect 240769 -9174 240869 -9050
rect 243913 -9114 244057 -8877
rect 244243 -8899 244629 -8877
rect 244167 -8985 244629 -8899
rect 247257 -8874 247333 -8832
rect 247385 -8874 247973 -8819
rect 250667 -8832 250677 -8819
rect 247257 -8877 247973 -8874
rect 244171 -8993 244371 -8985
rect 244187 -8997 244355 -8993
rect 240769 -9228 240771 -9174
rect 243913 -9200 244087 -9114
rect 244113 -9174 244213 -9050
rect 247257 -9114 247401 -8877
rect 247587 -8899 247973 -8877
rect 247511 -8985 247973 -8899
rect 250601 -8874 250677 -8832
rect 250729 -8874 251317 -8819
rect 254011 -8832 254021 -8819
rect 250601 -8877 251317 -8874
rect 247515 -8993 247715 -8985
rect 247531 -8997 247699 -8993
rect 244113 -9228 244115 -9174
rect 247257 -9200 247431 -9114
rect 247457 -9174 247557 -9050
rect 250601 -9114 250745 -8877
rect 250931 -8899 251317 -8877
rect 250855 -8985 251317 -8899
rect 253945 -8874 254021 -8832
rect 254073 -8874 254661 -8819
rect 257355 -8832 257365 -8819
rect 253945 -8877 254661 -8874
rect 250859 -8993 251059 -8985
rect 250875 -8997 251043 -8993
rect 247457 -9228 247459 -9174
rect 250601 -9200 250775 -9114
rect 250801 -9174 250901 -9050
rect 253945 -9114 254089 -8877
rect 254275 -8899 254661 -8877
rect 254199 -8985 254661 -8899
rect 257289 -8874 257365 -8832
rect 257417 -8874 258005 -8819
rect 260699 -8832 260709 -8819
rect 257289 -8877 258005 -8874
rect 254203 -8993 254403 -8985
rect 254219 -8997 254387 -8993
rect 250801 -9228 250803 -9174
rect 253945 -9200 254119 -9114
rect 254145 -9174 254245 -9050
rect 257289 -9114 257433 -8877
rect 257619 -8899 258005 -8877
rect 257543 -8985 258005 -8899
rect 260633 -8874 260709 -8832
rect 260761 -8874 261349 -8819
rect 264043 -8832 264053 -8819
rect 260633 -8877 261349 -8874
rect 257547 -8993 257747 -8985
rect 257563 -8997 257731 -8993
rect 254145 -9228 254147 -9174
rect 257289 -9200 257463 -9114
rect 257489 -9174 257589 -9050
rect 260633 -9114 260777 -8877
rect 260963 -8899 261349 -8877
rect 260887 -8985 261349 -8899
rect 263977 -8874 264053 -8832
rect 264105 -8874 264693 -8819
rect 267387 -8832 267397 -8819
rect 263977 -8877 264693 -8874
rect 260891 -8993 261091 -8985
rect 260907 -8997 261075 -8993
rect 257489 -9228 257491 -9174
rect 260633 -9200 260807 -9114
rect 260833 -9174 260933 -9050
rect 263977 -9114 264121 -8877
rect 264307 -8899 264693 -8877
rect 264231 -8985 264693 -8899
rect 267321 -8874 267397 -8832
rect 267449 -8874 268037 -8819
rect 270731 -8832 270741 -8819
rect 267321 -8877 268037 -8874
rect 264235 -8993 264435 -8985
rect 264251 -8997 264419 -8993
rect 260833 -9228 260835 -9174
rect 263977 -9200 264151 -9114
rect 264177 -9174 264277 -9050
rect 267321 -9114 267465 -8877
rect 267651 -8899 268037 -8877
rect 267575 -8985 268037 -8899
rect 270665 -8874 270741 -8832
rect 270793 -8874 271381 -8819
rect 274075 -8832 274085 -8819
rect 270665 -8877 271381 -8874
rect 267579 -8993 267779 -8985
rect 267595 -8997 267763 -8993
rect 264177 -9228 264179 -9174
rect 267321 -9200 267495 -9114
rect 267521 -9174 267621 -9050
rect 270665 -9114 270809 -8877
rect 270995 -8899 271381 -8877
rect 270919 -8985 271381 -8899
rect 274009 -8874 274085 -8832
rect 274137 -8874 274725 -8819
rect 277419 -8832 277429 -8819
rect 274009 -8877 274725 -8874
rect 270923 -8993 271123 -8985
rect 270939 -8997 271107 -8993
rect 267521 -9228 267523 -9174
rect 270665 -9200 270839 -9114
rect 270865 -9174 270965 -9050
rect 274009 -9114 274153 -8877
rect 274339 -8899 274725 -8877
rect 274263 -8985 274725 -8899
rect 277353 -8874 277429 -8832
rect 277481 -8874 278069 -8819
rect 280763 -8832 280773 -8819
rect 277353 -8877 278069 -8874
rect 274267 -8993 274467 -8985
rect 274283 -8997 274451 -8993
rect 270865 -9228 270867 -9174
rect 274009 -9200 274183 -9114
rect 274209 -9174 274309 -9050
rect 277353 -9114 277497 -8877
rect 277683 -8899 278069 -8877
rect 277607 -8985 278069 -8899
rect 280697 -8874 280773 -8832
rect 280825 -8874 281413 -8819
rect 284107 -8832 284117 -8819
rect 280697 -8877 281413 -8874
rect 277611 -8993 277811 -8985
rect 277627 -8997 277795 -8993
rect 274209 -9228 274211 -9174
rect 277353 -9200 277527 -9114
rect 277553 -9174 277653 -9050
rect 280697 -9114 280841 -8877
rect 281027 -8899 281413 -8877
rect 280951 -8985 281413 -8899
rect 284041 -8874 284117 -8832
rect 284169 -8874 284757 -8819
rect 287451 -8832 287461 -8819
rect 284041 -8877 284757 -8874
rect 280955 -8993 281155 -8985
rect 280971 -8997 281139 -8993
rect 277553 -9228 277555 -9174
rect 280697 -9200 280871 -9114
rect 280897 -9174 280997 -9050
rect 284041 -9114 284185 -8877
rect 284371 -8899 284757 -8877
rect 284295 -8985 284757 -8899
rect 287385 -8874 287461 -8832
rect 287513 -8874 288101 -8819
rect 290795 -8832 290805 -8819
rect 287385 -8877 288101 -8874
rect 284299 -8993 284499 -8985
rect 284315 -8997 284483 -8993
rect 280897 -9228 280899 -9174
rect 284041 -9200 284215 -9114
rect 284241 -9174 284341 -9050
rect 287385 -9114 287529 -8877
rect 287715 -8899 288101 -8877
rect 287639 -8985 288101 -8899
rect 290729 -8874 290805 -8832
rect 290857 -8874 291445 -8819
rect 294139 -8832 294149 -8819
rect 290729 -8877 291445 -8874
rect 287643 -8993 287843 -8985
rect 287659 -8997 287827 -8993
rect 284241 -9228 284243 -9174
rect 287385 -9200 287559 -9114
rect 287585 -9174 287685 -9050
rect 290729 -9114 290873 -8877
rect 291059 -8899 291445 -8877
rect 290983 -8985 291445 -8899
rect 294073 -8874 294149 -8832
rect 294201 -8874 294789 -8819
rect 297483 -8832 297493 -8819
rect 294073 -8877 294789 -8874
rect 290987 -8993 291187 -8985
rect 291003 -8997 291171 -8993
rect 287585 -9228 287587 -9174
rect 290729 -9200 290903 -9114
rect 290929 -9174 291029 -9050
rect 294073 -9114 294217 -8877
rect 294403 -8899 294789 -8877
rect 294327 -8985 294789 -8899
rect 297417 -8874 297493 -8832
rect 297545 -8874 298133 -8819
rect 300827 -8832 300837 -8819
rect 297417 -8877 298133 -8874
rect 294331 -8993 294531 -8985
rect 294347 -8997 294515 -8993
rect 290929 -9228 290931 -9174
rect 294073 -9200 294247 -9114
rect 294273 -9174 294373 -9050
rect 297417 -9114 297561 -8877
rect 297747 -8899 298133 -8877
rect 297671 -8985 298133 -8899
rect 300761 -8874 300837 -8832
rect 300889 -8874 301477 -8819
rect 304171 -8832 304181 -8819
rect 300761 -8877 301477 -8874
rect 297675 -8993 297875 -8985
rect 297691 -8997 297859 -8993
rect 294273 -9228 294275 -9174
rect 297417 -9200 297591 -9114
rect 297617 -9174 297717 -9050
rect 300761 -9114 300905 -8877
rect 301091 -8899 301477 -8877
rect 301015 -8985 301477 -8899
rect 304105 -8874 304181 -8832
rect 304233 -8874 304821 -8819
rect 307515 -8832 307525 -8819
rect 304105 -8877 304821 -8874
rect 301019 -8993 301219 -8985
rect 301035 -8997 301203 -8993
rect 297617 -9228 297619 -9174
rect 300761 -9200 300935 -9114
rect 300961 -9174 301061 -9050
rect 304105 -9114 304249 -8877
rect 304435 -8899 304821 -8877
rect 304359 -8985 304821 -8899
rect 307449 -8874 307525 -8832
rect 307577 -8874 308165 -8819
rect 310859 -8832 310869 -8819
rect 307449 -8877 308165 -8874
rect 304363 -8993 304563 -8985
rect 304379 -8997 304547 -8993
rect 300961 -9228 300963 -9174
rect 304105 -9200 304279 -9114
rect 304305 -9174 304405 -9050
rect 307449 -9114 307593 -8877
rect 307779 -8899 308165 -8877
rect 307703 -8985 308165 -8899
rect 310793 -8874 310869 -8832
rect 310921 -8874 311509 -8819
rect 314203 -8832 314213 -8819
rect 310793 -8877 311509 -8874
rect 307707 -8993 307907 -8985
rect 307723 -8997 307891 -8993
rect 304305 -9228 304307 -9174
rect 307449 -9200 307623 -9114
rect 307649 -9174 307749 -9050
rect 310793 -9114 310937 -8877
rect 311123 -8899 311509 -8877
rect 311047 -8985 311509 -8899
rect 314137 -8874 314213 -8832
rect 314265 -8874 314853 -8819
rect 317547 -8832 317557 -8819
rect 314137 -8877 314853 -8874
rect 311051 -8993 311251 -8985
rect 311067 -8997 311235 -8993
rect 307649 -9228 307651 -9174
rect 310793 -9200 310967 -9114
rect 310993 -9174 311093 -9050
rect 314137 -9114 314281 -8877
rect 314467 -8899 314853 -8877
rect 314391 -8985 314853 -8899
rect 317481 -8874 317557 -8832
rect 317609 -8874 318197 -8819
rect 320891 -8832 320901 -8819
rect 317481 -8877 318197 -8874
rect 314395 -8993 314595 -8985
rect 314411 -8997 314579 -8993
rect 310993 -9228 310995 -9174
rect 314137 -9200 314311 -9114
rect 314337 -9174 314437 -9050
rect 317481 -9114 317625 -8877
rect 317811 -8899 318197 -8877
rect 317735 -8985 318197 -8899
rect 320825 -8874 320901 -8832
rect 320953 -8874 321541 -8819
rect 324235 -8832 324245 -8819
rect 320825 -8877 321541 -8874
rect 317739 -8993 317939 -8985
rect 317755 -8997 317923 -8993
rect 314337 -9228 314339 -9174
rect 317481 -9200 317655 -9114
rect 317681 -9174 317781 -9050
rect 320825 -9114 320969 -8877
rect 321155 -8899 321541 -8877
rect 321079 -8985 321541 -8899
rect 324169 -8874 324245 -8832
rect 324297 -8874 324885 -8819
rect 327579 -8832 327589 -8819
rect 324169 -8877 324885 -8874
rect 321083 -8993 321283 -8985
rect 321099 -8997 321267 -8993
rect 317681 -9228 317683 -9174
rect 320825 -9200 320999 -9114
rect 321025 -9174 321125 -9050
rect 324169 -9114 324313 -8877
rect 324499 -8899 324885 -8877
rect 324423 -8985 324885 -8899
rect 327513 -8874 327589 -8832
rect 327641 -8874 328229 -8819
rect 330923 -8832 330933 -8819
rect 327513 -8877 328229 -8874
rect 324427 -8993 324627 -8985
rect 324443 -8997 324611 -8993
rect 321025 -9228 321027 -9174
rect 324169 -9200 324343 -9114
rect 324369 -9174 324469 -9050
rect 327513 -9114 327657 -8877
rect 327843 -8899 328229 -8877
rect 327767 -8985 328229 -8899
rect 330857 -8874 330933 -8832
rect 330985 -8874 331573 -8819
rect 334267 -8832 334277 -8819
rect 330857 -8877 331573 -8874
rect 327771 -8993 327971 -8985
rect 327787 -8997 327955 -8993
rect 324369 -9228 324371 -9174
rect 327513 -9200 327687 -9114
rect 327713 -9174 327813 -9050
rect 330857 -9114 331001 -8877
rect 331187 -8899 331573 -8877
rect 331111 -8985 331573 -8899
rect 334201 -8874 334277 -8832
rect 334329 -8874 334917 -8819
rect 337611 -8832 337621 -8819
rect 334201 -8877 334917 -8874
rect 331115 -8993 331315 -8985
rect 331131 -8997 331299 -8993
rect 327713 -9228 327715 -9174
rect 330857 -9200 331031 -9114
rect 331057 -9174 331157 -9050
rect 334201 -9114 334345 -8877
rect 334531 -8899 334917 -8877
rect 334455 -8985 334917 -8899
rect 337545 -8874 337621 -8832
rect 337673 -8874 338261 -8819
rect 340955 -8832 340965 -8819
rect 337545 -8877 338261 -8874
rect 334459 -8993 334659 -8985
rect 334475 -8997 334643 -8993
rect 331057 -9228 331059 -9174
rect 334201 -9200 334375 -9114
rect 334401 -9174 334501 -9050
rect 337545 -9114 337689 -8877
rect 337875 -8899 338261 -8877
rect 337799 -8985 338261 -8899
rect 340889 -8874 340965 -8832
rect 341017 -8874 341605 -8819
rect 344299 -8832 344309 -8819
rect 340889 -8877 341605 -8874
rect 337803 -8993 338003 -8985
rect 337819 -8997 337987 -8993
rect 334401 -9228 334403 -9174
rect 337545 -9200 337719 -9114
rect 337745 -9174 337845 -9050
rect 340889 -9114 341033 -8877
rect 341219 -8899 341605 -8877
rect 341143 -8985 341605 -8899
rect 344233 -8874 344309 -8832
rect 344361 -8874 344949 -8819
rect 347643 -8832 347653 -8819
rect 344233 -8877 344949 -8874
rect 341147 -8993 341347 -8985
rect 341163 -8997 341331 -8993
rect 337745 -9228 337747 -9174
rect 340889 -9200 341063 -9114
rect 341089 -9174 341189 -9050
rect 344233 -9114 344377 -8877
rect 344563 -8899 344949 -8877
rect 344487 -8985 344949 -8899
rect 347577 -8874 347653 -8832
rect 347705 -8874 348293 -8819
rect 350987 -8832 350997 -8819
rect 347577 -8877 348293 -8874
rect 344491 -8993 344691 -8985
rect 344507 -8997 344675 -8993
rect 341089 -9228 341091 -9174
rect 344233 -9200 344407 -9114
rect 344433 -9174 344533 -9050
rect 347577 -9114 347721 -8877
rect 347907 -8899 348293 -8877
rect 347831 -8985 348293 -8899
rect 350921 -8874 350997 -8832
rect 351049 -8874 351637 -8819
rect 354331 -8832 354341 -8819
rect 350921 -8877 351637 -8874
rect 347835 -8993 348035 -8985
rect 347851 -8997 348019 -8993
rect 344433 -9228 344435 -9174
rect 347577 -9200 347751 -9114
rect 347777 -9174 347877 -9050
rect 350921 -9114 351065 -8877
rect 351251 -8899 351637 -8877
rect 351175 -8985 351637 -8899
rect 354265 -8874 354341 -8832
rect 354393 -8874 354981 -8819
rect 357675 -8832 357685 -8819
rect 354265 -8877 354981 -8874
rect 351179 -8993 351379 -8985
rect 351195 -8997 351363 -8993
rect 347777 -9228 347779 -9174
rect 350921 -9200 351095 -9114
rect 351121 -9174 351221 -9050
rect 354265 -9114 354409 -8877
rect 354595 -8899 354981 -8877
rect 354519 -8985 354981 -8899
rect 357609 -8874 357685 -8832
rect 357737 -8874 358325 -8819
rect 361019 -8832 361029 -8819
rect 357609 -8877 358325 -8874
rect 354523 -8993 354723 -8985
rect 354539 -8997 354707 -8993
rect 351121 -9228 351123 -9174
rect 354265 -9200 354439 -9114
rect 354465 -9174 354565 -9050
rect 357609 -9114 357753 -8877
rect 357939 -8899 358325 -8877
rect 357863 -8985 358325 -8899
rect 360953 -8874 361029 -8832
rect 361081 -8874 361669 -8819
rect 364363 -8832 364373 -8819
rect 360953 -8877 361669 -8874
rect 357867 -8993 358067 -8985
rect 357883 -8997 358051 -8993
rect 354465 -9228 354467 -9174
rect 357609 -9200 357783 -9114
rect 357809 -9174 357909 -9050
rect 360953 -9114 361097 -8877
rect 361283 -8899 361669 -8877
rect 361207 -8985 361669 -8899
rect 364297 -8874 364373 -8832
rect 364425 -8874 365013 -8819
rect 367707 -8832 367717 -8819
rect 364297 -8877 365013 -8874
rect 361211 -8993 361411 -8985
rect 361227 -8997 361395 -8993
rect 357809 -9228 357811 -9174
rect 360953 -9200 361127 -9114
rect 361153 -9174 361253 -9050
rect 364297 -9114 364441 -8877
rect 364627 -8899 365013 -8877
rect 364551 -8985 365013 -8899
rect 367641 -8874 367717 -8832
rect 367769 -8874 368357 -8819
rect 371051 -8832 371061 -8819
rect 367641 -8877 368357 -8874
rect 364555 -8993 364755 -8985
rect 364571 -8997 364739 -8993
rect 361153 -9228 361155 -9174
rect 364297 -9200 364471 -9114
rect 364497 -9174 364597 -9050
rect 367641 -9114 367785 -8877
rect 367971 -8899 368357 -8877
rect 367895 -8985 368357 -8899
rect 370985 -8874 371061 -8832
rect 371113 -8874 371701 -8819
rect 374395 -8832 374405 -8819
rect 370985 -8877 371701 -8874
rect 367899 -8993 368099 -8985
rect 367915 -8997 368083 -8993
rect 364497 -9228 364499 -9174
rect 367641 -9200 367815 -9114
rect 367841 -9174 367941 -9050
rect 370985 -9114 371129 -8877
rect 371315 -8899 371701 -8877
rect 371239 -8985 371701 -8899
rect 374329 -8874 374405 -8832
rect 374457 -8874 375045 -8819
rect 377739 -8832 377749 -8819
rect 374329 -8877 375045 -8874
rect 371243 -8993 371443 -8985
rect 371259 -8997 371427 -8993
rect 367841 -9228 367843 -9174
rect 370985 -9200 371159 -9114
rect 371185 -9174 371285 -9050
rect 374329 -9114 374473 -8877
rect 374659 -8899 375045 -8877
rect 374583 -8985 375045 -8899
rect 377673 -8874 377749 -8832
rect 377801 -8874 378389 -8819
rect 381083 -8832 381093 -8819
rect 377673 -8877 378389 -8874
rect 374587 -8993 374787 -8985
rect 374603 -8997 374771 -8993
rect 371185 -9228 371187 -9174
rect 374329 -9200 374503 -9114
rect 374529 -9174 374629 -9050
rect 377673 -9114 377817 -8877
rect 378003 -8899 378389 -8877
rect 377927 -8985 378389 -8899
rect 381017 -8874 381093 -8832
rect 381145 -8874 381733 -8819
rect 384427 -8832 384437 -8819
rect 381017 -8877 381733 -8874
rect 377931 -8993 378131 -8985
rect 377947 -8997 378115 -8993
rect 374529 -9228 374531 -9174
rect 377673 -9200 377847 -9114
rect 377873 -9174 377973 -9050
rect 381017 -9114 381161 -8877
rect 381347 -8899 381733 -8877
rect 381271 -8985 381733 -8899
rect 384361 -8874 384437 -8832
rect 384489 -8874 385077 -8819
rect 387771 -8832 387781 -8819
rect 384361 -8877 385077 -8874
rect 381275 -8993 381475 -8985
rect 381291 -8997 381459 -8993
rect 377873 -9228 377875 -9174
rect 381017 -9200 381191 -9114
rect 381217 -9174 381317 -9050
rect 384361 -9114 384505 -8877
rect 384691 -8899 385077 -8877
rect 384615 -8985 385077 -8899
rect 387705 -8874 387781 -8832
rect 387833 -8874 388421 -8819
rect 391115 -8832 391125 -8819
rect 387705 -8877 388421 -8874
rect 384619 -8993 384819 -8985
rect 384635 -8997 384803 -8993
rect 381217 -9228 381219 -9174
rect 384361 -9200 384535 -9114
rect 384561 -9174 384661 -9050
rect 387705 -9114 387849 -8877
rect 388035 -8899 388421 -8877
rect 387959 -8985 388421 -8899
rect 391049 -8874 391125 -8832
rect 391177 -8874 391765 -8819
rect 394459 -8832 394469 -8819
rect 391049 -8877 391765 -8874
rect 387963 -8993 388163 -8985
rect 387979 -8997 388147 -8993
rect 384561 -9228 384563 -9174
rect 387705 -9200 387879 -9114
rect 387905 -9174 388005 -9050
rect 391049 -9114 391193 -8877
rect 391379 -8899 391765 -8877
rect 391303 -8985 391765 -8899
rect 394393 -8874 394469 -8832
rect 394521 -8874 395109 -8819
rect 397803 -8832 397813 -8819
rect 394393 -8877 395109 -8874
rect 391307 -8993 391507 -8985
rect 391323 -8997 391491 -8993
rect 387905 -9228 387907 -9174
rect 391049 -9200 391223 -9114
rect 391249 -9174 391349 -9050
rect 394393 -9114 394537 -8877
rect 394723 -8899 395109 -8877
rect 394647 -8985 395109 -8899
rect 397737 -8874 397813 -8832
rect 397865 -8874 398453 -8819
rect 401147 -8832 401157 -8819
rect 397737 -8877 398453 -8874
rect 394651 -8993 394851 -8985
rect 394667 -8997 394835 -8993
rect 391249 -9228 391251 -9174
rect 394393 -9200 394567 -9114
rect 394593 -9174 394693 -9050
rect 397737 -9114 397881 -8877
rect 398067 -8899 398453 -8877
rect 397991 -8985 398453 -8899
rect 401081 -8874 401157 -8832
rect 401209 -8874 401797 -8819
rect 404491 -8832 404501 -8819
rect 401081 -8877 401797 -8874
rect 397995 -8993 398195 -8985
rect 398011 -8997 398179 -8993
rect 394593 -9228 394595 -9174
rect 397737 -9200 397911 -9114
rect 397937 -9174 398037 -9050
rect 401081 -9114 401225 -8877
rect 401411 -8899 401797 -8877
rect 401335 -8985 401797 -8899
rect 404425 -8874 404501 -8832
rect 404553 -8874 405141 -8819
rect 407835 -8832 407845 -8819
rect 404425 -8877 405141 -8874
rect 401339 -8993 401539 -8985
rect 401355 -8997 401523 -8993
rect 397937 -9228 397939 -9174
rect 401081 -9200 401255 -9114
rect 401281 -9174 401381 -9050
rect 404425 -9114 404569 -8877
rect 404755 -8899 405141 -8877
rect 404679 -8985 405141 -8899
rect 407769 -8874 407845 -8832
rect 407897 -8874 408485 -8819
rect 411179 -8832 411189 -8819
rect 407769 -8877 408485 -8874
rect 404683 -8993 404883 -8985
rect 404699 -8997 404867 -8993
rect 401281 -9228 401283 -9174
rect 404425 -9200 404599 -9114
rect 404625 -9174 404725 -9050
rect 407769 -9114 407913 -8877
rect 408099 -8899 408485 -8877
rect 408023 -8985 408485 -8899
rect 411113 -8874 411189 -8832
rect 411241 -8874 411829 -8819
rect 414523 -8832 414533 -8819
rect 411113 -8877 411829 -8874
rect 408027 -8993 408227 -8985
rect 408043 -8997 408211 -8993
rect 404625 -9228 404627 -9174
rect 407769 -9200 407943 -9114
rect 407969 -9174 408069 -9050
rect 411113 -9114 411257 -8877
rect 411443 -8899 411829 -8877
rect 411367 -8985 411829 -8899
rect 414457 -8874 414533 -8832
rect 414585 -8874 415173 -8819
rect 417867 -8832 417877 -8819
rect 414457 -8877 415173 -8874
rect 411371 -8993 411571 -8985
rect 411387 -8997 411555 -8993
rect 407969 -9228 407971 -9174
rect 411113 -9200 411287 -9114
rect 411313 -9174 411413 -9050
rect 414457 -9114 414601 -8877
rect 414787 -8899 415173 -8877
rect 414711 -8985 415173 -8899
rect 417801 -8874 417877 -8832
rect 417929 -8874 418517 -8819
rect 421211 -8832 421221 -8819
rect 417801 -8877 418517 -8874
rect 414715 -8993 414915 -8985
rect 414731 -8997 414899 -8993
rect 411313 -9228 411315 -9174
rect 414457 -9200 414631 -9114
rect 414657 -9174 414757 -9050
rect 417801 -9114 417945 -8877
rect 418131 -8899 418517 -8877
rect 418055 -8985 418517 -8899
rect 421145 -8874 421221 -8832
rect 421273 -8874 421861 -8819
rect 424555 -8832 424565 -8819
rect 421145 -8877 421861 -8874
rect 418059 -8993 418259 -8985
rect 418075 -8997 418243 -8993
rect 414657 -9228 414659 -9174
rect 417801 -9200 417975 -9114
rect 418001 -9174 418101 -9050
rect 421145 -9114 421289 -8877
rect 421475 -8899 421861 -8877
rect 421399 -8985 421861 -8899
rect 424489 -8874 424565 -8832
rect 424617 -8874 425205 -8819
rect 427899 -8832 427909 -8819
rect 424489 -8877 425205 -8874
rect 421403 -8993 421603 -8985
rect 421419 -8997 421587 -8993
rect 418001 -9228 418003 -9174
rect 421145 -9200 421319 -9114
rect 421345 -9174 421445 -9050
rect 424489 -9114 424633 -8877
rect 424819 -8899 425205 -8877
rect 424743 -8985 425205 -8899
rect 427833 -8874 427909 -8832
rect 424747 -8993 424947 -8985
rect 424763 -8997 424931 -8993
rect 421345 -9228 421347 -9174
rect 424489 -9200 424663 -9114
rect 424689 -9174 424789 -9050
rect 427833 -9114 427977 -8874
rect 424689 -9228 424691 -9174
rect 427833 -9200 428007 -9114
rect 428033 -9174 428133 -9050
rect 428033 -9228 428035 -9174
rect 217046 -9971 217190 -9924
rect 217227 -9971 217244 -9870
rect 220390 -9971 220534 -9924
rect 220571 -9971 220588 -9870
rect 223734 -9971 223878 -9924
rect 223915 -9971 223932 -9870
rect 227078 -9971 227222 -9924
rect 227259 -9971 227276 -9870
rect 230422 -9971 230566 -9924
rect 230603 -9971 230620 -9870
rect 233766 -9971 233910 -9924
rect 233947 -9971 233964 -9870
rect 237110 -9971 237254 -9924
rect 237291 -9971 237308 -9870
rect 240454 -9971 240598 -9924
rect 240635 -9971 240652 -9870
rect 243798 -9971 243942 -9924
rect 243979 -9971 243996 -9870
rect 247142 -9971 247286 -9924
rect 247323 -9971 247340 -9870
rect 250486 -9971 250630 -9924
rect 250667 -9971 250684 -9870
rect 253830 -9971 253974 -9924
rect 254011 -9971 254028 -9870
rect 257174 -9971 257318 -9924
rect 257355 -9971 257372 -9870
rect 260518 -9971 260662 -9924
rect 260699 -9971 260716 -9870
rect 263862 -9971 264006 -9924
rect 264043 -9971 264060 -9870
rect 267206 -9971 267350 -9924
rect 267387 -9971 267404 -9870
rect 270550 -9971 270694 -9924
rect 270731 -9971 270748 -9870
rect 273894 -9971 274038 -9924
rect 274075 -9971 274092 -9870
rect 277238 -9971 277382 -9924
rect 277419 -9971 277436 -9870
rect 280582 -9971 280726 -9924
rect 280763 -9971 280780 -9870
rect 283926 -9971 284070 -9924
rect 284107 -9971 284124 -9870
rect 287270 -9971 287414 -9924
rect 287451 -9971 287468 -9870
rect 290614 -9971 290758 -9924
rect 290795 -9971 290812 -9870
rect 293958 -9971 294102 -9924
rect 294139 -9971 294156 -9870
rect 297302 -9971 297446 -9924
rect 297483 -9971 297500 -9870
rect 300646 -9971 300790 -9924
rect 300827 -9971 300844 -9870
rect 303990 -9971 304134 -9924
rect 304171 -9971 304188 -9870
rect 307334 -9971 307478 -9924
rect 307515 -9971 307532 -9870
rect 310678 -9971 310822 -9924
rect 310859 -9971 310876 -9870
rect 314022 -9971 314166 -9924
rect 314203 -9971 314220 -9870
rect 317366 -9971 317510 -9924
rect 317547 -9971 317564 -9870
rect 320710 -9971 320854 -9924
rect 320891 -9971 320908 -9870
rect 324054 -9971 324198 -9924
rect 324235 -9971 324252 -9870
rect 327398 -9971 327542 -9924
rect 327579 -9971 327596 -9870
rect 330742 -9971 330886 -9924
rect 330923 -9971 330940 -9870
rect 334086 -9971 334230 -9924
rect 334267 -9971 334284 -9870
rect 337430 -9971 337574 -9924
rect 337611 -9971 337628 -9870
rect 340774 -9971 340918 -9924
rect 340955 -9971 340972 -9870
rect 344118 -9971 344262 -9924
rect 344299 -9971 344316 -9870
rect 347462 -9971 347606 -9924
rect 347643 -9971 347660 -9870
rect 350806 -9971 350950 -9924
rect 350987 -9971 351004 -9870
rect 354150 -9971 354294 -9924
rect 354331 -9971 354348 -9870
rect 357494 -9971 357638 -9924
rect 357675 -9971 357692 -9870
rect 360838 -9971 360982 -9924
rect 361019 -9971 361036 -9870
rect 364182 -9971 364326 -9924
rect 364363 -9971 364380 -9870
rect 367526 -9971 367670 -9924
rect 367707 -9971 367724 -9870
rect 370870 -9971 371014 -9924
rect 371051 -9971 371068 -9870
rect 374214 -9971 374358 -9924
rect 374395 -9971 374412 -9870
rect 377558 -9971 377702 -9924
rect 377739 -9971 377756 -9870
rect 380902 -9971 381046 -9924
rect 381083 -9971 381100 -9870
rect 384246 -9971 384390 -9924
rect 384427 -9971 384444 -9870
rect 387590 -9971 387734 -9924
rect 387771 -9971 387788 -9870
rect 390934 -9971 391078 -9924
rect 391115 -9971 391132 -9870
rect 394278 -9971 394422 -9924
rect 394459 -9971 394476 -9870
rect 397622 -9971 397766 -9924
rect 397803 -9971 397820 -9870
rect 400966 -9971 401110 -9924
rect 401147 -9971 401164 -9870
rect 404310 -9971 404454 -9924
rect 404491 -9971 404508 -9870
rect 407654 -9971 407798 -9924
rect 407835 -9971 407852 -9870
rect 410998 -9971 411142 -9924
rect 411179 -9971 411196 -9870
rect 414342 -9971 414486 -9924
rect 414523 -9971 414540 -9870
rect 417686 -9971 417830 -9924
rect 417867 -9971 417884 -9870
rect 421030 -9971 421174 -9924
rect 421211 -9971 421228 -9870
rect 424374 -9971 424518 -9924
rect 424555 -9971 424572 -9870
rect 427718 -9971 427862 -9924
rect 427899 -9971 427916 -9870
rect 217046 -9982 217162 -9971
rect 217132 -10007 217162 -9982
rect 217144 -10506 217162 -10007
rect 220390 -9982 221162 -9971
rect 223734 -9982 224506 -9971
rect 227078 -9982 227850 -9971
rect 230422 -9982 231194 -9971
rect 233766 -9982 234538 -9971
rect 237110 -9982 237882 -9971
rect 240454 -9982 241226 -9971
rect 243798 -9982 244570 -9971
rect 247142 -9982 247914 -9971
rect 250486 -9982 251258 -9971
rect 253830 -9982 254602 -9971
rect 257174 -9982 257946 -9971
rect 260518 -9982 261290 -9971
rect 263862 -9982 264634 -9971
rect 267206 -9982 267978 -9971
rect 270550 -9982 271322 -9971
rect 273894 -9982 274666 -9971
rect 277238 -9982 278010 -9971
rect 280582 -9982 281354 -9971
rect 283926 -9982 284698 -9971
rect 287270 -9982 288042 -9971
rect 290614 -9982 291386 -9971
rect 293958 -9982 294730 -9971
rect 297302 -9982 298074 -9971
rect 300646 -9982 301418 -9971
rect 303990 -9982 304762 -9971
rect 307334 -9982 308106 -9971
rect 310678 -9982 311450 -9971
rect 314022 -9982 314794 -9971
rect 317366 -9982 318138 -9971
rect 320710 -9982 321482 -9971
rect 324054 -9982 324826 -9971
rect 327398 -9982 328170 -9971
rect 330742 -9982 331514 -9971
rect 334086 -9982 334858 -9971
rect 337430 -9982 338202 -9971
rect 340774 -9982 341546 -9971
rect 344118 -9982 344890 -9971
rect 347462 -9982 348234 -9971
rect 350806 -9982 351578 -9971
rect 354150 -9982 354922 -9971
rect 357494 -9982 358266 -9971
rect 360838 -9982 361610 -9971
rect 364182 -9982 364954 -9971
rect 367526 -9982 368298 -9971
rect 370870 -9982 371642 -9971
rect 374214 -9982 374986 -9971
rect 377558 -9982 378330 -9971
rect 380902 -9982 381674 -9971
rect 384246 -9982 385018 -9971
rect 387590 -9982 388362 -9971
rect 390934 -9982 391706 -9971
rect 394278 -9982 395050 -9971
rect 397622 -9982 398394 -9971
rect 400966 -9982 401738 -9971
rect 404310 -9982 405082 -9971
rect 407654 -9982 408426 -9971
rect 410998 -9982 411770 -9971
rect 414342 -9982 415114 -9971
rect 417686 -9982 418458 -9971
rect 421030 -9982 421802 -9971
rect 424374 -9982 425146 -9971
rect 427718 -9982 428490 -9971
rect 220476 -10007 221162 -9982
rect 223820 -10007 224506 -9982
rect 227164 -10007 227850 -9982
rect 230508 -10007 231194 -9982
rect 233852 -10007 234538 -9982
rect 237196 -10007 237882 -9982
rect 240540 -10007 241226 -9982
rect 243884 -10007 244570 -9982
rect 247228 -10007 247914 -9982
rect 250572 -10007 251258 -9982
rect 253916 -10007 254602 -9982
rect 257260 -10007 257946 -9982
rect 260604 -10007 261290 -9982
rect 263948 -10007 264634 -9982
rect 267292 -10007 267978 -9982
rect 270636 -10007 271322 -9982
rect 273980 -10007 274666 -9982
rect 277324 -10007 278010 -9982
rect 280668 -10007 281354 -9982
rect 284012 -10007 284698 -9982
rect 287356 -10007 288042 -9982
rect 290700 -10007 291386 -9982
rect 294044 -10007 294730 -9982
rect 297388 -10007 298074 -9982
rect 300732 -10007 301418 -9982
rect 304076 -10007 304762 -9982
rect 307420 -10007 308106 -9982
rect 310764 -10007 311450 -9982
rect 314108 -10007 314794 -9982
rect 317452 -10007 318138 -9982
rect 320796 -10007 321482 -9982
rect 324140 -10007 324826 -9982
rect 327484 -10007 328170 -9982
rect 330828 -10007 331514 -9982
rect 334172 -10007 334858 -9982
rect 337516 -10007 338202 -9982
rect 340860 -10007 341546 -9982
rect 344204 -10007 344890 -9982
rect 347548 -10007 348234 -9982
rect 350892 -10007 351578 -9982
rect 354236 -10007 354922 -9982
rect 357580 -10007 358266 -9982
rect 360924 -10007 361610 -9982
rect 364268 -10007 364954 -9982
rect 367612 -10007 368298 -9982
rect 370956 -10007 371642 -9982
rect 374300 -10007 374986 -9982
rect 377644 -10007 378330 -9982
rect 380988 -10007 381674 -9982
rect 384332 -10007 385018 -9982
rect 387676 -10007 388362 -9982
rect 391020 -10007 391706 -9982
rect 394364 -10007 395050 -9982
rect 397708 -10007 398394 -9982
rect 401052 -10007 401738 -9982
rect 404396 -10007 405082 -9982
rect 407740 -10007 408426 -9982
rect 411084 -10007 411770 -9982
rect 414428 -10007 415114 -9982
rect 417772 -10007 418458 -9982
rect 421116 -10007 421802 -9982
rect 424460 -10007 425146 -9982
rect 427804 -10007 428490 -9982
rect 220488 -10036 221162 -10007
rect 223832 -10036 224506 -10007
rect 227176 -10036 227850 -10007
rect 230520 -10036 231194 -10007
rect 233864 -10036 234538 -10007
rect 237208 -10036 237882 -10007
rect 240552 -10036 241226 -10007
rect 243896 -10036 244570 -10007
rect 247240 -10036 247914 -10007
rect 250584 -10036 251258 -10007
rect 253928 -10036 254602 -10007
rect 257272 -10036 257946 -10007
rect 260616 -10036 261290 -10007
rect 263960 -10036 264634 -10007
rect 267304 -10036 267978 -10007
rect 270648 -10036 271322 -10007
rect 273992 -10036 274666 -10007
rect 277336 -10036 278010 -10007
rect 280680 -10036 281354 -10007
rect 284024 -10036 284698 -10007
rect 287368 -10036 288042 -10007
rect 290712 -10036 291386 -10007
rect 294056 -10036 294730 -10007
rect 297400 -10036 298074 -10007
rect 300744 -10036 301418 -10007
rect 304088 -10036 304762 -10007
rect 307432 -10036 308106 -10007
rect 310776 -10036 311450 -10007
rect 314120 -10036 314794 -10007
rect 317464 -10036 318138 -10007
rect 320808 -10036 321482 -10007
rect 324152 -10036 324826 -10007
rect 327496 -10036 328170 -10007
rect 330840 -10036 331514 -10007
rect 334184 -10036 334858 -10007
rect 337528 -10036 338202 -10007
rect 340872 -10036 341546 -10007
rect 344216 -10036 344890 -10007
rect 347560 -10036 348234 -10007
rect 350904 -10036 351578 -10007
rect 354248 -10036 354922 -10007
rect 357592 -10036 358266 -10007
rect 360936 -10036 361610 -10007
rect 364280 -10036 364954 -10007
rect 367624 -10036 368298 -10007
rect 370968 -10036 371642 -10007
rect 374312 -10036 374986 -10007
rect 377656 -10036 378330 -10007
rect 381000 -10036 381674 -10007
rect 384344 -10036 385018 -10007
rect 387688 -10036 388362 -10007
rect 391032 -10036 391706 -10007
rect 394376 -10036 395050 -10007
rect 397720 -10036 398394 -10007
rect 401064 -10036 401738 -10007
rect 404408 -10036 405082 -10007
rect 407752 -10036 408426 -10007
rect 411096 -10036 411770 -10007
rect 414440 -10036 415114 -10007
rect 417784 -10036 418458 -10007
rect 421128 -10036 421802 -10007
rect 424472 -10036 425146 -10007
rect 427816 -10036 428490 -10007
rect 218326 -10448 218373 -10083
rect 218380 -10448 218427 -10137
rect 220488 -10448 221221 -10036
rect 221670 -10448 221717 -10083
rect 221724 -10448 221771 -10137
rect 223832 -10448 224565 -10036
rect 225014 -10448 225061 -10083
rect 225068 -10448 225115 -10137
rect 227176 -10448 227909 -10036
rect 228358 -10448 228405 -10083
rect 228412 -10448 228459 -10137
rect 230520 -10448 231253 -10036
rect 231702 -10448 231749 -10083
rect 231756 -10448 231803 -10137
rect 233864 -10448 234597 -10036
rect 235046 -10448 235093 -10083
rect 235100 -10448 235147 -10137
rect 237208 -10448 237941 -10036
rect 238390 -10448 238437 -10083
rect 238444 -10448 238491 -10137
rect 240552 -10448 241285 -10036
rect 241734 -10448 241781 -10083
rect 241788 -10448 241835 -10137
rect 243896 -10448 244629 -10036
rect 245078 -10448 245125 -10083
rect 245132 -10448 245179 -10137
rect 247240 -10448 247973 -10036
rect 248422 -10448 248469 -10083
rect 248476 -10448 248523 -10137
rect 250584 -10448 251317 -10036
rect 251766 -10448 251813 -10083
rect 251820 -10448 251867 -10137
rect 253928 -10448 254661 -10036
rect 255110 -10448 255157 -10083
rect 255164 -10448 255211 -10137
rect 257272 -10448 258005 -10036
rect 258454 -10448 258501 -10083
rect 258508 -10448 258555 -10137
rect 260616 -10448 261349 -10036
rect 261798 -10448 261845 -10083
rect 261852 -10448 261899 -10137
rect 263960 -10448 264693 -10036
rect 265142 -10448 265189 -10083
rect 265196 -10448 265243 -10137
rect 267304 -10448 268037 -10036
rect 268486 -10448 268533 -10083
rect 268540 -10448 268587 -10137
rect 270648 -10448 271381 -10036
rect 271830 -10448 271877 -10083
rect 271884 -10448 271931 -10137
rect 273992 -10448 274725 -10036
rect 275174 -10448 275221 -10083
rect 275228 -10448 275275 -10137
rect 277336 -10448 278069 -10036
rect 278518 -10448 278565 -10083
rect 278572 -10448 278619 -10137
rect 280680 -10448 281413 -10036
rect 281862 -10448 281909 -10083
rect 281916 -10448 281963 -10137
rect 284024 -10448 284757 -10036
rect 285206 -10448 285253 -10083
rect 285260 -10448 285307 -10137
rect 287368 -10448 288101 -10036
rect 288550 -10448 288597 -10083
rect 288604 -10448 288651 -10137
rect 290712 -10448 291445 -10036
rect 291894 -10448 291941 -10083
rect 291948 -10448 291995 -10137
rect 294056 -10448 294789 -10036
rect 295238 -10448 295285 -10083
rect 295292 -10448 295339 -10137
rect 297400 -10448 298133 -10036
rect 298582 -10448 298629 -10083
rect 298636 -10448 298683 -10137
rect 300744 -10448 301477 -10036
rect 301926 -10448 301973 -10083
rect 301980 -10448 302027 -10137
rect 304088 -10448 304821 -10036
rect 305270 -10448 305317 -10083
rect 305324 -10448 305371 -10137
rect 307432 -10448 308165 -10036
rect 308614 -10448 308661 -10083
rect 308668 -10448 308715 -10137
rect 310776 -10448 311509 -10036
rect 311958 -10448 312005 -10083
rect 312012 -10448 312059 -10137
rect 314120 -10448 314853 -10036
rect 315302 -10448 315349 -10083
rect 315356 -10448 315403 -10137
rect 317464 -10448 318197 -10036
rect 318646 -10448 318693 -10083
rect 318700 -10448 318747 -10137
rect 320808 -10448 321541 -10036
rect 321990 -10448 322037 -10083
rect 322044 -10448 322091 -10137
rect 324152 -10448 324885 -10036
rect 325334 -10448 325381 -10083
rect 325388 -10448 325435 -10137
rect 327496 -10448 328229 -10036
rect 328678 -10448 328725 -10083
rect 328732 -10448 328779 -10137
rect 330840 -10448 331573 -10036
rect 332022 -10448 332069 -10083
rect 332076 -10448 332123 -10137
rect 334184 -10448 334917 -10036
rect 335366 -10448 335413 -10083
rect 335420 -10448 335467 -10137
rect 337528 -10448 338261 -10036
rect 338710 -10448 338757 -10083
rect 338764 -10448 338811 -10137
rect 340872 -10448 341605 -10036
rect 342054 -10448 342101 -10083
rect 342108 -10448 342155 -10137
rect 344216 -10448 344949 -10036
rect 345398 -10448 345445 -10083
rect 345452 -10448 345499 -10137
rect 347560 -10448 348293 -10036
rect 348742 -10448 348789 -10083
rect 348796 -10448 348843 -10137
rect 350904 -10448 351637 -10036
rect 352086 -10448 352133 -10083
rect 352140 -10448 352187 -10137
rect 354248 -10448 354981 -10036
rect 355430 -10448 355477 -10083
rect 355484 -10448 355531 -10137
rect 357592 -10448 358325 -10036
rect 358774 -10448 358821 -10083
rect 358828 -10448 358875 -10137
rect 360936 -10448 361669 -10036
rect 362118 -10448 362165 -10083
rect 362172 -10448 362219 -10137
rect 364280 -10448 365013 -10036
rect 365462 -10448 365509 -10083
rect 365516 -10448 365563 -10137
rect 367624 -10448 368357 -10036
rect 368806 -10448 368853 -10083
rect 368860 -10448 368907 -10137
rect 370968 -10448 371701 -10036
rect 372150 -10448 372197 -10083
rect 372204 -10448 372251 -10137
rect 374312 -10448 375045 -10036
rect 375494 -10448 375541 -10083
rect 375548 -10448 375595 -10137
rect 377656 -10448 378389 -10036
rect 378838 -10448 378885 -10083
rect 378892 -10448 378939 -10137
rect 381000 -10448 381733 -10036
rect 382182 -10448 382229 -10083
rect 382236 -10448 382283 -10137
rect 384344 -10448 385077 -10036
rect 385526 -10448 385573 -10083
rect 385580 -10448 385627 -10137
rect 387688 -10448 388421 -10036
rect 388870 -10448 388917 -10083
rect 388924 -10448 388971 -10137
rect 391032 -10448 391765 -10036
rect 392214 -10448 392261 -10083
rect 392268 -10448 392315 -10137
rect 394376 -10448 395109 -10036
rect 395558 -10448 395605 -10083
rect 395612 -10448 395659 -10137
rect 397720 -10448 398453 -10036
rect 398902 -10448 398949 -10083
rect 398956 -10448 399003 -10137
rect 401064 -10448 401797 -10036
rect 402246 -10448 402293 -10083
rect 402300 -10448 402347 -10137
rect 404408 -10448 405141 -10036
rect 405590 -10448 405637 -10083
rect 405644 -10448 405691 -10137
rect 407752 -10448 408485 -10036
rect 408934 -10448 408981 -10083
rect 408988 -10448 409035 -10137
rect 411096 -10448 411829 -10036
rect 412278 -10448 412325 -10083
rect 412332 -10448 412379 -10137
rect 414440 -10448 415173 -10036
rect 415622 -10448 415669 -10083
rect 415676 -10448 415723 -10137
rect 417784 -10448 418517 -10036
rect 418966 -10448 419013 -10083
rect 419020 -10448 419067 -10137
rect 421128 -10448 421861 -10036
rect 422310 -10448 422357 -10083
rect 422364 -10448 422411 -10137
rect 424472 -10448 425205 -10036
rect 425654 -10448 425701 -10083
rect 425708 -10448 425755 -10137
rect 427816 -10448 428549 -10036
rect 428998 -10448 429045 -10083
rect 429052 -10448 429099 -10137
rect 218294 -10543 218498 -10448
rect 220488 -10506 221842 -10448
rect 223832 -10506 225186 -10448
rect 227176 -10506 228530 -10448
rect 230520 -10506 231874 -10448
rect 233864 -10506 235218 -10448
rect 237208 -10506 238562 -10448
rect 240552 -10506 241906 -10448
rect 243896 -10506 245250 -10448
rect 247240 -10506 248594 -10448
rect 250584 -10506 251938 -10448
rect 253928 -10506 255282 -10448
rect 257272 -10506 258626 -10448
rect 260616 -10506 261970 -10448
rect 263960 -10506 265314 -10448
rect 267304 -10506 268658 -10448
rect 270648 -10506 272002 -10448
rect 273992 -10506 275346 -10448
rect 277336 -10506 278690 -10448
rect 280680 -10506 282034 -10448
rect 284024 -10506 285378 -10448
rect 287368 -10506 288722 -10448
rect 290712 -10506 292066 -10448
rect 294056 -10506 295410 -10448
rect 297400 -10506 298754 -10448
rect 300744 -10506 302098 -10448
rect 304088 -10506 305442 -10448
rect 307432 -10506 308786 -10448
rect 310776 -10506 312130 -10448
rect 314120 -10506 315474 -10448
rect 317464 -10506 318818 -10448
rect 320808 -10506 322162 -10448
rect 324152 -10506 325506 -10448
rect 327496 -10506 328850 -10448
rect 330840 -10506 332194 -10448
rect 334184 -10506 335538 -10448
rect 337528 -10506 338882 -10448
rect 340872 -10506 342226 -10448
rect 344216 -10506 345570 -10448
rect 347560 -10506 348914 -10448
rect 350904 -10506 352258 -10448
rect 354248 -10506 355602 -10448
rect 357592 -10506 358946 -10448
rect 360936 -10506 362290 -10448
rect 364280 -10506 365634 -10448
rect 367624 -10506 368978 -10448
rect 370968 -10506 372322 -10448
rect 374312 -10506 375666 -10448
rect 377656 -10506 379010 -10448
rect 381000 -10506 382354 -10448
rect 384344 -10506 385698 -10448
rect 387688 -10506 389042 -10448
rect 391032 -10506 392386 -10448
rect 394376 -10506 395730 -10448
rect 397720 -10506 399074 -10448
rect 401064 -10506 402418 -10448
rect 404408 -10506 405762 -10448
rect 407752 -10506 409106 -10448
rect 411096 -10506 412450 -10448
rect 414440 -10506 415794 -10448
rect 417784 -10506 419138 -10448
rect 421128 -10506 422482 -10448
rect 424472 -10506 425826 -10448
rect 427816 -10506 429170 -10448
rect 219915 -10543 221842 -10506
rect 223259 -10543 225186 -10506
rect 226603 -10543 228530 -10506
rect 229947 -10543 231874 -10506
rect 233291 -10543 235218 -10506
rect 236635 -10543 238562 -10506
rect 239979 -10543 241906 -10506
rect 243323 -10543 245250 -10506
rect 246667 -10543 248594 -10506
rect 250011 -10543 251938 -10506
rect 253355 -10543 255282 -10506
rect 256699 -10543 258626 -10506
rect 260043 -10543 261970 -10506
rect 263387 -10543 265314 -10506
rect 266731 -10543 268658 -10506
rect 270075 -10543 272002 -10506
rect 273419 -10543 275346 -10506
rect 276763 -10543 278690 -10506
rect 280107 -10543 282034 -10506
rect 283451 -10543 285378 -10506
rect 286795 -10543 288722 -10506
rect 290139 -10543 292066 -10506
rect 293483 -10543 295410 -10506
rect 296827 -10543 298754 -10506
rect 300171 -10543 302098 -10506
rect 303515 -10543 305442 -10506
rect 306859 -10543 308786 -10506
rect 310203 -10543 312130 -10506
rect 313547 -10543 315474 -10506
rect 316891 -10543 318818 -10506
rect 320235 -10543 322162 -10506
rect 323579 -10543 325506 -10506
rect 326923 -10543 328850 -10506
rect 330267 -10543 332194 -10506
rect 333611 -10543 335538 -10506
rect 336955 -10543 338882 -10506
rect 340299 -10543 342226 -10506
rect 343643 -10543 345570 -10506
rect 346987 -10543 348914 -10506
rect 350331 -10543 352258 -10506
rect 353675 -10543 355602 -10506
rect 357019 -10543 358946 -10506
rect 360363 -10543 362290 -10506
rect 363707 -10543 365634 -10506
rect 367051 -10543 368978 -10506
rect 370395 -10543 372322 -10506
rect 373739 -10543 375666 -10506
rect 377083 -10543 379010 -10506
rect 380427 -10543 382354 -10506
rect 383771 -10543 385698 -10506
rect 387115 -10543 389042 -10506
rect 390459 -10543 392386 -10506
rect 393803 -10543 395730 -10506
rect 397147 -10543 399074 -10506
rect 400491 -10543 402418 -10506
rect 403835 -10543 405762 -10506
rect 407179 -10543 409106 -10506
rect 410523 -10543 412450 -10506
rect 413867 -10543 415794 -10506
rect 417211 -10543 419138 -10506
rect 420555 -10543 422482 -10506
rect 423899 -10543 425826 -10506
rect 427243 -10543 429170 -10506
rect 218294 -10667 219000 -10543
rect 219915 -10667 222344 -10543
rect 223259 -10667 225688 -10543
rect 226603 -10667 229032 -10543
rect 229947 -10667 232376 -10543
rect 233291 -10667 235720 -10543
rect 236635 -10667 239064 -10543
rect 239979 -10667 242408 -10543
rect 243323 -10667 245752 -10543
rect 246667 -10667 249096 -10543
rect 250011 -10667 252440 -10543
rect 253355 -10667 255784 -10543
rect 256699 -10667 259128 -10543
rect 260043 -10667 262472 -10543
rect 263387 -10667 265816 -10543
rect 266731 -10667 269160 -10543
rect 270075 -10667 272504 -10543
rect 273419 -10667 275848 -10543
rect 276763 -10667 279192 -10543
rect 280107 -10667 282536 -10543
rect 283451 -10667 285880 -10543
rect 286795 -10667 289224 -10543
rect 290139 -10667 292568 -10543
rect 293483 -10667 295912 -10543
rect 296827 -10667 299256 -10543
rect 300171 -10667 302600 -10543
rect 303515 -10667 305944 -10543
rect 306859 -10667 309288 -10543
rect 310203 -10667 312632 -10543
rect 313547 -10667 315976 -10543
rect 316891 -10667 319320 -10543
rect 320235 -10667 322664 -10543
rect 323579 -10667 326008 -10543
rect 326923 -10667 329352 -10543
rect 330267 -10667 332696 -10543
rect 333611 -10667 336040 -10543
rect 336955 -10667 339384 -10543
rect 340299 -10667 342728 -10543
rect 343643 -10667 346072 -10543
rect 346987 -10667 349416 -10543
rect 350331 -10667 352760 -10543
rect 353675 -10667 356104 -10543
rect 357019 -10667 359448 -10543
rect 360363 -10667 362792 -10543
rect 363707 -10667 366136 -10543
rect 367051 -10667 369480 -10543
rect 370395 -10667 372824 -10543
rect 373739 -10667 376168 -10543
rect 377083 -10667 379512 -10543
rect 380427 -10667 382856 -10543
rect 383771 -10667 386200 -10543
rect 387115 -10667 389544 -10543
rect 390459 -10667 392888 -10543
rect 393803 -10667 396232 -10543
rect 397147 -10667 399576 -10543
rect 400491 -10667 402920 -10543
rect 403835 -10667 406264 -10543
rect 407179 -10667 409608 -10543
rect 410523 -10667 412952 -10543
rect 413867 -10667 416296 -10543
rect 417211 -10667 419640 -10543
rect 420555 -10667 422984 -10543
rect 423899 -10667 426328 -10543
rect 427243 -10667 429672 -10543
rect 218294 -11752 219053 -10667
rect 219915 -11622 222397 -10667
rect 223259 -11622 225741 -10667
rect 226603 -11622 229085 -10667
rect 229947 -11622 232429 -10667
rect 233291 -11622 235773 -10667
rect 236635 -11622 239117 -10667
rect 239979 -11622 242461 -10667
rect 243323 -11622 245805 -10667
rect 246667 -11622 249149 -10667
rect 250011 -11622 252493 -10667
rect 253355 -11622 255837 -10667
rect 256699 -11622 259181 -10667
rect 260043 -11622 262525 -10667
rect 263387 -11622 265869 -10667
rect 266731 -11622 269213 -10667
rect 270075 -11622 272557 -10667
rect 273419 -11622 275901 -10667
rect 276763 -11622 279245 -10667
rect 280107 -11622 282589 -10667
rect 283451 -11622 285933 -10667
rect 286795 -11622 289277 -10667
rect 290139 -11622 292621 -10667
rect 293483 -11622 295965 -10667
rect 296827 -11622 299309 -10667
rect 300171 -11622 302653 -10667
rect 303515 -11622 305997 -10667
rect 306859 -11622 309341 -10667
rect 310203 -11622 312685 -10667
rect 313547 -11622 316029 -10667
rect 316891 -11622 319373 -10667
rect 320235 -11622 322717 -10667
rect 323579 -11622 326061 -10667
rect 326923 -11622 329405 -10667
rect 330267 -11622 332749 -10667
rect 333611 -11622 336093 -10667
rect 336955 -11622 339437 -10667
rect 340299 -11622 342781 -10667
rect 343643 -11622 346125 -10667
rect 346987 -11622 349469 -10667
rect 350331 -11622 352813 -10667
rect 353675 -11622 356157 -10667
rect 357019 -11622 359501 -10667
rect 360363 -11622 362845 -10667
rect 363707 -11622 366189 -10667
rect 367051 -11622 369533 -10667
rect 370395 -11622 372877 -10667
rect 373739 -11622 376221 -10667
rect 377083 -11622 379565 -10667
rect 380427 -11622 382909 -10667
rect 383771 -11622 386253 -10667
rect 387115 -11622 389597 -10667
rect 390459 -11622 392941 -10667
rect 393803 -11622 396285 -10667
rect 397147 -11622 399629 -10667
rect 400491 -11622 402973 -10667
rect 403835 -11622 406317 -10667
rect 407179 -11622 409661 -10667
rect 410523 -11622 413005 -10667
rect 413867 -11622 416349 -10667
rect 417211 -11622 419693 -10667
rect 420555 -11622 423037 -10667
rect 423899 -11622 426381 -10667
rect 427243 -11622 429725 -10667
rect 220506 -11687 222397 -11622
rect 223850 -11687 225741 -11622
rect 227194 -11687 229085 -11622
rect 230538 -11687 232429 -11622
rect 233882 -11687 235773 -11622
rect 237226 -11687 239117 -11622
rect 240570 -11687 242461 -11622
rect 243914 -11687 245805 -11622
rect 247258 -11687 249149 -11622
rect 250602 -11687 252493 -11622
rect 253946 -11687 255837 -11622
rect 257290 -11687 259181 -11622
rect 260634 -11687 262525 -11622
rect 263978 -11687 265869 -11622
rect 267322 -11687 269213 -11622
rect 270666 -11687 272557 -11622
rect 274010 -11687 275901 -11622
rect 277354 -11687 279245 -11622
rect 280698 -11687 282589 -11622
rect 284042 -11687 285933 -11622
rect 287386 -11687 289277 -11622
rect 290730 -11687 292621 -11622
rect 294074 -11687 295965 -11622
rect 297418 -11687 299309 -11622
rect 300762 -11687 302653 -11622
rect 304106 -11687 305997 -11622
rect 307450 -11687 309341 -11622
rect 310794 -11687 312685 -11622
rect 314138 -11687 316029 -11622
rect 317482 -11687 319373 -11622
rect 320826 -11687 322717 -11622
rect 324170 -11687 326061 -11622
rect 327514 -11687 329405 -11622
rect 330858 -11687 332749 -11622
rect 334202 -11687 336093 -11622
rect 337546 -11687 339437 -11622
rect 340890 -11687 342781 -11622
rect 344234 -11687 346125 -11622
rect 347578 -11687 349469 -11622
rect 350922 -11687 352813 -11622
rect 354266 -11687 356157 -11622
rect 357610 -11687 359501 -11622
rect 360954 -11687 362845 -11622
rect 364298 -11687 366189 -11622
rect 367642 -11687 369533 -11622
rect 370986 -11687 372877 -11622
rect 374330 -11687 376221 -11622
rect 377674 -11687 379565 -11622
rect 381018 -11687 382909 -11622
rect 384362 -11687 386253 -11622
rect 387706 -11687 389597 -11622
rect 391050 -11687 392941 -11622
rect 394394 -11687 396285 -11622
rect 397738 -11687 399629 -11622
rect 401082 -11687 402973 -11622
rect 404426 -11687 406317 -11622
rect 407770 -11687 409661 -11622
rect 411114 -11687 413005 -11622
rect 414458 -11687 416349 -11622
rect 417802 -11687 419693 -11622
rect 421146 -11687 423037 -11622
rect 424490 -11687 426381 -11622
rect 427834 -11687 429725 -11622
rect 221097 -11747 222397 -11687
rect 224441 -11747 225741 -11687
rect 227785 -11747 229085 -11687
rect 231129 -11747 232429 -11687
rect 234473 -11747 235773 -11687
rect 237817 -11747 239117 -11687
rect 241161 -11747 242461 -11687
rect 244505 -11747 245805 -11687
rect 247849 -11747 249149 -11687
rect 251193 -11747 252493 -11687
rect 254537 -11747 255837 -11687
rect 257881 -11747 259181 -11687
rect 261225 -11747 262525 -11687
rect 264569 -11747 265869 -11687
rect 267913 -11747 269213 -11687
rect 271257 -11747 272557 -11687
rect 274601 -11747 275901 -11687
rect 277945 -11747 279245 -11687
rect 281289 -11747 282589 -11687
rect 284633 -11747 285933 -11687
rect 287977 -11747 289277 -11687
rect 291321 -11747 292621 -11687
rect 294665 -11747 295965 -11687
rect 298009 -11747 299309 -11687
rect 301353 -11747 302653 -11687
rect 304697 -11747 305997 -11687
rect 308041 -11747 309341 -11687
rect 311385 -11747 312685 -11687
rect 314729 -11747 316029 -11687
rect 318073 -11747 319373 -11687
rect 321417 -11747 322717 -11687
rect 324761 -11747 326061 -11687
rect 328105 -11747 329405 -11687
rect 331449 -11747 332749 -11687
rect 334793 -11747 336093 -11687
rect 338137 -11747 339437 -11687
rect 341481 -11747 342781 -11687
rect 344825 -11747 346125 -11687
rect 348169 -11747 349469 -11687
rect 351513 -11747 352813 -11687
rect 354857 -11747 356157 -11687
rect 358201 -11747 359501 -11687
rect 361545 -11747 362845 -11687
rect 364889 -11747 366189 -11687
rect 368233 -11747 369533 -11687
rect 371577 -11747 372877 -11687
rect 374921 -11747 376221 -11687
rect 378265 -11747 379565 -11687
rect 381609 -11747 382909 -11687
rect 384953 -11747 386253 -11687
rect 388297 -11747 389597 -11687
rect 391641 -11747 392941 -11687
rect 394985 -11747 396285 -11687
rect 398329 -11747 399629 -11687
rect 401673 -11747 402973 -11687
rect 405017 -11747 406317 -11687
rect 408361 -11747 409661 -11687
rect 411705 -11747 413005 -11687
rect 415049 -11747 416349 -11687
rect 418393 -11747 419693 -11687
rect 421737 -11747 423037 -11687
rect 425081 -11747 426381 -11687
rect 428425 -11747 429725 -11687
rect 221126 -11752 222397 -11747
rect 224470 -11752 225741 -11747
rect 227814 -11752 229085 -11747
rect 231158 -11752 232429 -11747
rect 234502 -11752 235773 -11747
rect 237846 -11752 239117 -11747
rect 241190 -11752 242461 -11747
rect 244534 -11752 245805 -11747
rect 247878 -11752 249149 -11747
rect 251222 -11752 252493 -11747
rect 254566 -11752 255837 -11747
rect 257910 -11752 259181 -11747
rect 261254 -11752 262525 -11747
rect 264598 -11752 265869 -11747
rect 267942 -11752 269213 -11747
rect 271286 -11752 272557 -11747
rect 274630 -11752 275901 -11747
rect 277974 -11752 279245 -11747
rect 281318 -11752 282589 -11747
rect 284662 -11752 285933 -11747
rect 288006 -11752 289277 -11747
rect 291350 -11752 292621 -11747
rect 294694 -11752 295965 -11747
rect 298038 -11752 299309 -11747
rect 301382 -11752 302653 -11747
rect 304726 -11752 305997 -11747
rect 308070 -11752 309341 -11747
rect 311414 -11752 312685 -11747
rect 314758 -11752 316029 -11747
rect 318102 -11752 319373 -11747
rect 321446 -11752 322717 -11747
rect 324790 -11752 326061 -11747
rect 328134 -11752 329405 -11747
rect 331478 -11752 332749 -11747
rect 334822 -11752 336093 -11747
rect 338166 -11752 339437 -11747
rect 341510 -11752 342781 -11747
rect 344854 -11752 346125 -11747
rect 348198 -11752 349469 -11747
rect 351542 -11752 352813 -11747
rect 354886 -11752 356157 -11747
rect 358230 -11752 359501 -11747
rect 361574 -11752 362845 -11747
rect 364918 -11752 366189 -11747
rect 368262 -11752 369533 -11747
rect 371606 -11752 372877 -11747
rect 374950 -11752 376221 -11747
rect 378294 -11752 379565 -11747
rect 381638 -11752 382909 -11747
rect 384982 -11752 386253 -11747
rect 388326 -11752 389597 -11747
rect 391670 -11752 392941 -11747
rect 395014 -11752 396285 -11747
rect 398358 -11752 399629 -11747
rect 401702 -11752 402973 -11747
rect 405046 -11752 406317 -11747
rect 408390 -11752 409661 -11747
rect 411734 -11752 413005 -11747
rect 415078 -11752 416349 -11747
rect 418422 -11752 419693 -11747
rect 421766 -11752 423037 -11747
rect 425110 -11752 426381 -11747
rect 428454 -11752 429725 -11747
rect 217906 -11770 219053 -11752
rect 221250 -11770 222397 -11752
rect 224594 -11770 225741 -11752
rect 227938 -11770 229085 -11752
rect 231282 -11770 232429 -11752
rect 234626 -11770 235773 -11752
rect 237970 -11770 239117 -11752
rect 241314 -11770 242461 -11752
rect 244658 -11770 245805 -11752
rect 248002 -11770 249149 -11752
rect 251346 -11770 252493 -11752
rect 254690 -11770 255837 -11752
rect 258034 -11770 259181 -11752
rect 261378 -11770 262525 -11752
rect 264722 -11770 265869 -11752
rect 268066 -11770 269213 -11752
rect 271410 -11770 272557 -11752
rect 274754 -11770 275901 -11752
rect 278098 -11770 279245 -11752
rect 281442 -11770 282589 -11752
rect 284786 -11770 285933 -11752
rect 288130 -11770 289277 -11752
rect 291474 -11770 292621 -11752
rect 294818 -11770 295965 -11752
rect 298162 -11770 299309 -11752
rect 301506 -11770 302653 -11752
rect 304850 -11770 305997 -11752
rect 308194 -11770 309341 -11752
rect 311538 -11770 312685 -11752
rect 314882 -11770 316029 -11752
rect 318226 -11770 319373 -11752
rect 321570 -11770 322717 -11752
rect 324914 -11770 326061 -11752
rect 328258 -11770 329405 -11752
rect 331602 -11770 332749 -11752
rect 334946 -11770 336093 -11752
rect 338290 -11770 339437 -11752
rect 341634 -11770 342781 -11752
rect 344978 -11770 346125 -11752
rect 348322 -11770 349469 -11752
rect 351666 -11770 352813 -11752
rect 355010 -11770 356157 -11752
rect 358354 -11770 359501 -11752
rect 361698 -11770 362845 -11752
rect 365042 -11770 366189 -11752
rect 368386 -11770 369533 -11752
rect 371730 -11770 372877 -11752
rect 375074 -11770 376221 -11752
rect 378418 -11770 379565 -11752
rect 381762 -11770 382909 -11752
rect 385106 -11770 386253 -11752
rect 388450 -11770 389597 -11752
rect 391794 -11770 392941 -11752
rect 395138 -11770 396285 -11752
rect 398482 -11770 399629 -11752
rect 401826 -11770 402973 -11752
rect 405170 -11770 406317 -11752
rect 408514 -11770 409661 -11752
rect 411858 -11770 413005 -11752
rect 415202 -11770 416349 -11752
rect 418546 -11770 419693 -11752
rect 421890 -11770 423037 -11752
rect 425234 -11770 426381 -11752
rect 428578 -11770 429725 -11752
rect 218344 -11781 219053 -11770
rect 221688 -11781 222397 -11770
rect 225032 -11781 225741 -11770
rect 228376 -11781 229085 -11770
rect 231720 -11781 232429 -11770
rect 235064 -11781 235773 -11770
rect 238408 -11781 239117 -11770
rect 241752 -11781 242461 -11770
rect 245096 -11781 245805 -11770
rect 248440 -11781 249149 -11770
rect 251784 -11781 252493 -11770
rect 255128 -11781 255837 -11770
rect 258472 -11781 259181 -11770
rect 261816 -11781 262525 -11770
rect 265160 -11781 265869 -11770
rect 268504 -11781 269213 -11770
rect 271848 -11781 272557 -11770
rect 275192 -11781 275901 -11770
rect 278536 -11781 279245 -11770
rect 281880 -11781 282589 -11770
rect 285224 -11781 285933 -11770
rect 288568 -11781 289277 -11770
rect 291912 -11781 292621 -11770
rect 295256 -11781 295965 -11770
rect 298600 -11781 299309 -11770
rect 301944 -11781 302653 -11770
rect 305288 -11781 305997 -11770
rect 308632 -11781 309341 -11770
rect 311976 -11781 312685 -11770
rect 315320 -11781 316029 -11770
rect 318664 -11781 319373 -11770
rect 322008 -11781 322717 -11770
rect 325352 -11781 326061 -11770
rect 328696 -11781 329405 -11770
rect 332040 -11781 332749 -11770
rect 335384 -11781 336093 -11770
rect 338728 -11781 339437 -11770
rect 342072 -11781 342781 -11770
rect 345416 -11781 346125 -11770
rect 348760 -11781 349469 -11770
rect 352104 -11781 352813 -11770
rect 355448 -11781 356157 -11770
rect 358792 -11781 359501 -11770
rect 362136 -11781 362845 -11770
rect 365480 -11781 366189 -11770
rect 368824 -11781 369533 -11770
rect 372168 -11781 372877 -11770
rect 375512 -11781 376221 -11770
rect 378856 -11781 379565 -11770
rect 382200 -11781 382909 -11770
rect 385544 -11781 386253 -11770
rect 388888 -11781 389597 -11770
rect 392232 -11781 392941 -11770
rect 395576 -11781 396285 -11770
rect 398920 -11781 399629 -11770
rect 402264 -11781 402973 -11770
rect 405608 -11781 406317 -11770
rect 408952 -11781 409661 -11770
rect 412296 -11781 413005 -11770
rect 415640 -11781 416349 -11770
rect 418984 -11781 419693 -11770
rect 422328 -11781 423037 -11770
rect 425672 -11781 426381 -11770
rect 429016 -11781 429725 -11770
rect 218344 -11817 219018 -11781
rect 221688 -11817 222362 -11781
rect 225032 -11817 225706 -11781
rect 228376 -11817 229050 -11781
rect 231720 -11817 232394 -11781
rect 235064 -11817 235738 -11781
rect 238408 -11817 239082 -11781
rect 241752 -11817 242426 -11781
rect 245096 -11817 245770 -11781
rect 248440 -11817 249114 -11781
rect 251784 -11817 252458 -11781
rect 255128 -11817 255802 -11781
rect 258472 -11817 259146 -11781
rect 261816 -11817 262490 -11781
rect 265160 -11817 265834 -11781
rect 268504 -11817 269178 -11781
rect 271848 -11817 272522 -11781
rect 275192 -11817 275866 -11781
rect 278536 -11817 279210 -11781
rect 281880 -11817 282554 -11781
rect 285224 -11817 285898 -11781
rect 288568 -11817 289242 -11781
rect 291912 -11817 292586 -11781
rect 295256 -11817 295930 -11781
rect 298600 -11817 299274 -11781
rect 301944 -11817 302618 -11781
rect 305288 -11817 305962 -11781
rect 308632 -11817 309306 -11781
rect 311976 -11817 312650 -11781
rect 315320 -11817 315994 -11781
rect 318664 -11817 319338 -11781
rect 322008 -11817 322682 -11781
rect 325352 -11817 326026 -11781
rect 328696 -11817 329370 -11781
rect 332040 -11817 332714 -11781
rect 335384 -11817 336058 -11781
rect 338728 -11817 339402 -11781
rect 342072 -11817 342746 -11781
rect 345416 -11817 346090 -11781
rect 348760 -11817 349434 -11781
rect 352104 -11817 352778 -11781
rect 355448 -11817 356122 -11781
rect 358792 -11817 359466 -11781
rect 362136 -11817 362810 -11781
rect 365480 -11817 366154 -11781
rect 368824 -11817 369498 -11781
rect 372168 -11817 372842 -11781
rect 375512 -11817 376186 -11781
rect 378856 -11817 379530 -11781
rect 382200 -11817 382874 -11781
rect 385544 -11817 386218 -11781
rect 388888 -11817 389562 -11781
rect 392232 -11817 392906 -11781
rect 395576 -11817 396250 -11781
rect 398920 -11817 399594 -11781
rect 402264 -11817 402938 -11781
rect 405608 -11817 406282 -11781
rect 408952 -11817 409626 -11781
rect 412296 -11817 412970 -11781
rect 415640 -11817 416314 -11781
rect 418984 -11817 419658 -11781
rect 422328 -11817 423002 -11781
rect 425672 -11817 426346 -11781
rect 429016 -11817 429690 -11781
rect 218527 -11835 219018 -11817
rect 221871 -11835 222362 -11817
rect 225215 -11835 225706 -11817
rect 228559 -11835 229050 -11817
rect 231903 -11835 232394 -11817
rect 235247 -11835 235738 -11817
rect 238591 -11835 239082 -11817
rect 241935 -11835 242426 -11817
rect 245279 -11835 245770 -11817
rect 248623 -11835 249114 -11817
rect 251967 -11835 252458 -11817
rect 255311 -11835 255802 -11817
rect 258655 -11835 259146 -11817
rect 261999 -11835 262490 -11817
rect 265343 -11835 265834 -11817
rect 268687 -11835 269178 -11817
rect 272031 -11835 272522 -11817
rect 275375 -11835 275866 -11817
rect 278719 -11835 279210 -11817
rect 282063 -11835 282554 -11817
rect 285407 -11835 285898 -11817
rect 288751 -11835 289242 -11817
rect 292095 -11835 292586 -11817
rect 295439 -11835 295930 -11817
rect 298783 -11835 299274 -11817
rect 302127 -11835 302618 -11817
rect 305471 -11835 305962 -11817
rect 308815 -11835 309306 -11817
rect 312159 -11835 312650 -11817
rect 315503 -11835 315994 -11817
rect 318847 -11835 319338 -11817
rect 322191 -11835 322682 -11817
rect 325535 -11835 326026 -11817
rect 328879 -11835 329370 -11817
rect 332223 -11835 332714 -11817
rect 335567 -11835 336058 -11817
rect 338911 -11835 339402 -11817
rect 342255 -11835 342746 -11817
rect 345599 -11835 346090 -11817
rect 348943 -11835 349434 -11817
rect 352287 -11835 352778 -11817
rect 355631 -11835 356122 -11817
rect 358975 -11835 359466 -11817
rect 362319 -11835 362810 -11817
rect 365663 -11835 366154 -11817
rect 369007 -11835 369498 -11817
rect 372351 -11835 372842 -11817
rect 375695 -11835 376186 -11817
rect 379039 -11835 379530 -11817
rect 382383 -11835 382874 -11817
rect 385727 -11835 386218 -11817
rect 389071 -11835 389562 -11817
rect 392415 -11835 392906 -11817
rect 395759 -11835 396250 -11817
rect 399103 -11835 399594 -11817
rect 402447 -11835 402938 -11817
rect 405791 -11835 406282 -11817
rect 409135 -11835 409626 -11817
rect 412479 -11835 412970 -11817
rect 415823 -11835 416314 -11817
rect 419167 -11835 419658 -11817
rect 422511 -11835 423002 -11817
rect 425855 -11835 426346 -11817
rect 429199 -11835 429690 -11817
<< error_s >>
rect 0 -5275 33 -3275
rect 121 -5179 437 -5167
rect 525 -5179 559 -3275
rect 3564 -4879 3707 -4788
rect 1135 -5179 2838 -5101
rect 121 -5213 2838 -5179
rect 121 -5225 437 -5213
rect 0 -5529 34 -5275
rect 133 -5342 167 -5225
rect 391 -5301 437 -5270
rect 525 -5279 559 -5213
rect 525 -5290 563 -5279
rect 379 -5317 437 -5301
rect 133 -5385 173 -5342
rect 180 -5351 437 -5317
rect 184 -5357 201 -5351
rect 133 -5410 167 -5385
rect 379 -5398 437 -5351
rect 513 -5301 524 -5290
rect 525 -5301 571 -5290
rect 133 -5529 168 -5410
rect 391 -5521 425 -5398
rect 381 -5529 425 -5521
rect 513 -5529 571 -5301
rect 1135 -5529 2838 -5213
rect -26 -5596 2838 -5529
rect 3364 -5462 3707 -4879
rect 3834 -5462 3868 -5440
rect 3364 -5474 3880 -5462
rect 3968 -5474 4002 -4665
rect 3364 -5508 4038 -5474
rect 3364 -5520 3880 -5508
rect 3968 -5518 4002 -5508
rect 3968 -5520 4088 -5518
rect 3364 -5596 3707 -5520
rect 3834 -5596 3880 -5565
rect -26 -5615 3707 -5596
rect 3822 -5612 3880 -5596
rect 0 -5623 34 -5615
rect 0 -5628 70 -5623
rect 0 -6149 34 -5628
rect 127 -5798 128 -5772
rect 133 -5786 168 -5615
rect 325 -5657 3707 -5615
rect 3770 -5646 3880 -5612
rect 3934 -5646 3954 -5612
rect 323 -5691 3707 -5657
rect 99 -5826 128 -5800
rect 134 -5971 168 -5786
rect 325 -5694 3707 -5691
rect 3822 -5693 3880 -5646
rect 325 -5705 3742 -5694
rect 325 -5798 3707 -5705
rect 179 -5845 180 -5798
rect 317 -5845 3707 -5798
rect 179 -5879 3707 -5845
rect 179 -5895 180 -5879
rect 325 -5971 3707 -5879
rect 122 -5983 3707 -5971
rect 100 -6017 3707 -5983
rect 122 -6029 3707 -6017
rect 544 -6070 3707 -6029
rect 542 -6117 3707 -6070
rect 544 -6138 3707 -6117
rect 542 -6149 3707 -6138
rect -47 -6421 3707 -6149
rect 3708 -6421 3742 -5705
rect -47 -6455 3742 -6421
rect 3834 -6421 3868 -5693
rect 3834 -6455 3892 -6421
rect 3956 -6455 4014 -5520
rect 4129 -5570 4146 -5508
rect 4654 -5518 4688 -4825
rect 5168 -5230 5226 -5078
rect 4642 -5557 4700 -5518
rect 4100 -5634 4146 -5570
rect 4183 -5634 4200 -5557
rect 4241 -5615 4767 -5557
rect 4642 -5634 4700 -5615
rect 4015 -6455 4700 -5634
rect -47 -6489 4700 -6455
rect -47 -6517 3707 -6489
rect 3708 -6517 3742 -6489
rect -47 -6586 3642 -6517
rect 3696 -6543 3753 -6517
rect 3708 -6544 3753 -6543
rect 3834 -6527 3868 -6489
rect 3956 -6517 4014 -6489
rect 3708 -6557 3809 -6544
rect 3834 -6557 3879 -6527
rect 3954 -6543 4014 -6517
rect -47 -6597 3653 -6586
rect 3679 -6589 3809 -6557
rect 3679 -6591 3798 -6589
rect 3823 -6591 3879 -6557
rect 3956 -6557 4014 -6543
rect 4015 -6557 4700 -6489
rect 3956 -6586 4700 -6557
rect -47 -6631 3658 -6597
rect -47 -6654 3642 -6631
rect 3645 -6654 3658 -6631
rect -47 -6699 3658 -6654
rect -47 -6722 3642 -6699
rect 3645 -6722 3658 -6699
rect -47 -6767 3658 -6722
rect -47 -6790 3642 -6767
rect 3645 -6790 3658 -6767
rect -47 -6835 3658 -6790
rect 3679 -6809 3692 -6591
rect 3708 -6612 3753 -6591
rect 3708 -6657 3809 -6612
rect 3708 -6680 3753 -6657
rect 3708 -6725 3809 -6680
rect 3708 -6748 3753 -6725
rect 3708 -6793 3809 -6748
rect 3708 -6809 3753 -6793
rect 3834 -6809 3879 -6591
rect 3954 -6591 4700 -6586
rect 3954 -6597 4014 -6591
rect 3891 -6654 3904 -6597
rect 3907 -6631 4014 -6597
rect 3956 -6654 4014 -6631
rect 3891 -6665 4014 -6654
rect 3891 -6722 3904 -6665
rect 3907 -6699 4014 -6665
rect 3956 -6722 4014 -6699
rect 3891 -6733 4014 -6722
rect 3891 -6790 3904 -6733
rect 3907 -6767 4014 -6733
rect 3956 -6790 4014 -6767
rect 3891 -6801 4014 -6790
rect -47 -6876 3642 -6835
rect 3645 -6843 3658 -6835
rect 3708 -6843 3742 -6809
rect 3696 -6873 3753 -6843
rect 3834 -6845 3868 -6809
rect 3891 -6843 3904 -6801
rect 3907 -6835 4014 -6801
rect 3956 -6843 4014 -6835
rect 3891 -6845 3902 -6843
rect 3696 -6876 3754 -6873
rect 3834 -6876 3879 -6845
rect 3954 -6876 4014 -6843
rect -47 -6923 3660 -6876
rect 3681 -6923 3796 -6876
rect 3817 -6879 3879 -6876
rect 3817 -6889 3868 -6879
rect 3804 -6923 3868 -6889
rect 3885 -6923 3932 -6876
rect 3953 -6923 4014 -6876
rect 4015 -6923 4700 -6591
rect -47 -6957 4700 -6923
rect -47 -6969 3642 -6957
rect 3696 -6969 3754 -6957
rect 3834 -6969 3879 -6957
rect 3954 -6969 4700 -6957
rect -47 -7265 4700 -6969
rect 544 -7295 4700 -7265
rect 1171 -7348 1218 -7295
rect 2743 -7301 4700 -7295
rect 2124 -7314 4700 -7301
rect 2743 -7329 4700 -7314
rect 2743 -7359 3620 -7329
rect 2743 -7373 3609 -7359
rect 3997 -7366 4014 -7329
rect 2743 -7378 3906 -7373
rect 4015 -7378 4700 -7329
rect 2743 -7390 4700 -7378
rect 3364 -7395 4700 -7390
rect 3488 -7407 4700 -7395
rect 3488 -7413 3609 -7407
rect 3670 -7412 4700 -7407
rect 4015 -7461 4700 -7412
rect 4709 -7461 4767 -5615
rect 4776 -7348 4821 -5503
rect 4788 -7352 4789 -7348
rect 4015 -7471 4688 -7461
rect 4721 -7467 4722 -7461
rect 4015 -7490 4671 -7471
rect 4687 -7473 4688 -7471
rect 4117 -7550 4671 -7490
rect 4700 -7499 4767 -7467
rect 4688 -7507 4767 -7499
rect 4700 -7519 4767 -7507
rect 4700 -7533 4821 -7521
rect 4688 -7541 4821 -7533
rect 4700 -7573 4821 -7541
rect 5209 -7579 5226 -5230
rect 5227 -5230 5292 -5194
rect 5227 -5288 5378 -5230
rect 5227 -7579 5321 -5288
rect 6445 -5754 6590 -5743
rect 6445 -5788 6553 -5754
rect 6445 -5800 6590 -5788
rect 5227 -7645 5292 -7579
rect 5800 -7674 5847 -5841
rect 6445 -5859 6503 -5800
rect 5854 -7728 5901 -5895
rect 6379 -7739 6503 -5859
rect 6579 -7573 6590 -5973
rect 6693 -7600 6759 -7586
rect 6665 -7628 6759 -7614
rect 6379 -7775 6492 -7739
rect 6445 -7791 6492 -7775
rect 6439 -7870 7095 -7791
rect 101 -8145 146 -8111
rect 197 -8145 242 -8111
rect 293 -8145 338 -8111
rect 389 -8145 434 -8111
rect 485 -8145 530 -8111
rect 3445 -8145 3490 -8111
rect 3541 -8145 3586 -8111
rect 3637 -8145 3682 -8111
rect 3733 -8145 3778 -8111
rect 3829 -8145 3874 -8111
rect 6790 -8145 6834 -8111
rect 6886 -8145 6930 -8111
rect 6982 -8145 7026 -8111
rect 7078 -8145 7122 -8111
rect 7174 -8145 7218 -8111
rect 10134 -8145 10178 -8111
rect 10230 -8145 10274 -8111
rect 10326 -8145 10370 -8111
rect 10422 -8145 10466 -8111
rect 10518 -8145 10562 -8111
rect 13479 -8145 13522 -8111
rect 13575 -8145 13618 -8111
rect 13671 -8145 13714 -8111
rect 13767 -8145 13810 -8111
rect 13863 -8145 13906 -8111
rect 16823 -8145 16866 -8111
rect 16919 -8145 16962 -8111
rect 17015 -8145 17058 -8111
rect 17111 -8145 17154 -8111
rect 17207 -8145 17250 -8111
rect 20167 -8145 20210 -8111
rect 20263 -8145 20306 -8111
rect 20359 -8145 20402 -8111
rect 20455 -8145 20498 -8111
rect 20551 -8145 20594 -8111
rect 23511 -8145 23554 -8111
rect 23607 -8145 23650 -8111
rect 23703 -8145 23746 -8111
rect 23799 -8145 23842 -8111
rect 23895 -8145 23938 -8111
rect 26856 -8145 26898 -8111
rect 26952 -8145 26994 -8111
rect 27048 -8145 27090 -8111
rect 27144 -8145 27186 -8111
rect 27240 -8145 27282 -8111
rect 30200 -8145 30242 -8111
rect 30296 -8145 30338 -8111
rect 30392 -8145 30434 -8111
rect 30488 -8145 30530 -8111
rect 30584 -8145 30626 -8111
rect 33544 -8145 33586 -8111
rect 33640 -8145 33682 -8111
rect 33736 -8145 33778 -8111
rect 33832 -8145 33874 -8111
rect 33928 -8145 33970 -8111
rect 36888 -8145 36930 -8111
rect 36984 -8145 37026 -8111
rect 37080 -8145 37122 -8111
rect 37176 -8145 37218 -8111
rect 37272 -8145 37314 -8111
rect 40232 -8145 40274 -8111
rect 40328 -8145 40370 -8111
rect 40424 -8145 40466 -8111
rect 40520 -8145 40562 -8111
rect 40616 -8145 40658 -8111
rect 43576 -8145 43618 -8111
rect 43672 -8145 43714 -8111
rect 43768 -8145 43810 -8111
rect 43864 -8145 43906 -8111
rect 43960 -8145 44002 -8111
rect 46920 -8145 46962 -8111
rect 47016 -8145 47058 -8111
rect 47112 -8145 47154 -8111
rect 47208 -8145 47250 -8111
rect 47304 -8145 47346 -8111
rect 50264 -8145 50306 -8111
rect 50360 -8145 50402 -8111
rect 50456 -8145 50498 -8111
rect 50552 -8145 50594 -8111
rect 50648 -8145 50690 -8111
rect 53609 -8145 53650 -8111
rect 53705 -8145 53746 -8111
rect 53801 -8145 53842 -8111
rect 53897 -8145 53938 -8111
rect 53993 -8145 54034 -8111
rect 56953 -8145 56994 -8111
rect 57049 -8145 57090 -8111
rect 57145 -8145 57186 -8111
rect 57241 -8145 57282 -8111
rect 57337 -8145 57378 -8111
rect 60297 -8145 60338 -8111
rect 60393 -8145 60434 -8111
rect 60489 -8145 60530 -8111
rect 60585 -8145 60626 -8111
rect 60681 -8145 60722 -8111
rect 63641 -8145 63682 -8111
rect 63737 -8145 63778 -8111
rect 63833 -8145 63874 -8111
rect 63929 -8145 63970 -8111
rect 64025 -8145 64066 -8111
rect 66985 -8145 67026 -8111
rect 67081 -8145 67122 -8111
rect 67177 -8145 67218 -8111
rect 67273 -8145 67314 -8111
rect 67369 -8145 67410 -8111
rect 70329 -8145 70370 -8111
rect 70425 -8145 70466 -8111
rect 70521 -8145 70562 -8111
rect 70617 -8145 70658 -8111
rect 70713 -8145 70754 -8111
rect 73673 -8145 73714 -8111
rect 73769 -8145 73810 -8111
rect 73865 -8145 73906 -8111
rect 73961 -8145 74002 -8111
rect 74057 -8145 74098 -8111
rect 77017 -8145 77058 -8111
rect 77113 -8145 77154 -8111
rect 77209 -8145 77250 -8111
rect 77305 -8145 77346 -8111
rect 77401 -8145 77442 -8111
rect 80361 -8145 80402 -8111
rect 80457 -8145 80498 -8111
rect 80553 -8145 80594 -8111
rect 80649 -8145 80690 -8111
rect 80745 -8145 80786 -8111
rect 83705 -8145 83746 -8111
rect 83801 -8145 83842 -8111
rect 83897 -8145 83938 -8111
rect 83993 -8145 84034 -8111
rect 84089 -8145 84130 -8111
rect 87049 -8145 87090 -8111
rect 87145 -8145 87186 -8111
rect 87241 -8145 87282 -8111
rect 87337 -8145 87378 -8111
rect 87433 -8145 87474 -8111
rect 90393 -8145 90434 -8111
rect 90489 -8145 90530 -8111
rect 90585 -8145 90626 -8111
rect 90681 -8145 90722 -8111
rect 90777 -8145 90818 -8111
rect 93737 -8145 93778 -8111
rect 93833 -8145 93874 -8111
rect 93929 -8145 93970 -8111
rect 94025 -8145 94066 -8111
rect 94121 -8145 94162 -8111
rect 97081 -8145 97122 -8111
rect 97177 -8145 97218 -8111
rect 97273 -8145 97314 -8111
rect 97369 -8145 97410 -8111
rect 97465 -8145 97506 -8111
rect 100425 -8145 100466 -8111
rect 100521 -8145 100562 -8111
rect 100617 -8145 100658 -8111
rect 100713 -8145 100754 -8111
rect 100809 -8145 100850 -8111
rect 103769 -8145 103810 -8111
rect 103865 -8145 103906 -8111
rect 103961 -8145 104002 -8111
rect 104057 -8145 104098 -8111
rect 104153 -8145 104194 -8111
rect 107119 -8145 107154 -8111
rect 107215 -8145 107250 -8111
rect 107311 -8145 107346 -8111
rect 107407 -8145 107442 -8111
rect 107503 -8145 107538 -8111
rect 110463 -8145 110498 -8111
rect 110559 -8145 110594 -8111
rect 110655 -8145 110690 -8111
rect 110751 -8145 110786 -8111
rect 110847 -8145 110882 -8111
rect 113807 -8145 113842 -8111
rect 113903 -8145 113938 -8111
rect 113999 -8145 114034 -8111
rect 114095 -8145 114130 -8111
rect 114191 -8145 114226 -8111
rect 117151 -8145 117186 -8111
rect 117247 -8145 117282 -8111
rect 117343 -8145 117378 -8111
rect 117439 -8145 117474 -8111
rect 117535 -8145 117570 -8111
rect 120495 -8145 120530 -8111
rect 120591 -8145 120626 -8111
rect 120687 -8145 120722 -8111
rect 120783 -8145 120818 -8111
rect 120879 -8145 120914 -8111
rect 123839 -8145 123874 -8111
rect 123935 -8145 123970 -8111
rect 124031 -8145 124066 -8111
rect 124127 -8145 124162 -8111
rect 124223 -8145 124258 -8111
rect 127183 -8145 127218 -8111
rect 127279 -8145 127314 -8111
rect 127375 -8145 127410 -8111
rect 127471 -8145 127506 -8111
rect 127567 -8145 127602 -8111
rect 130527 -8145 130562 -8111
rect 130623 -8145 130658 -8111
rect 130719 -8145 130754 -8111
rect 130815 -8145 130850 -8111
rect 130911 -8145 130946 -8111
rect 133871 -8145 133906 -8111
rect 133967 -8145 134002 -8111
rect 134063 -8145 134098 -8111
rect 134159 -8145 134194 -8111
rect 134255 -8145 134290 -8111
rect 137215 -8145 137250 -8111
rect 137311 -8145 137346 -8111
rect 137407 -8145 137442 -8111
rect 137503 -8145 137538 -8111
rect 137599 -8145 137634 -8111
rect 140559 -8145 140594 -8111
rect 140655 -8145 140690 -8111
rect 140751 -8145 140786 -8111
rect 140847 -8145 140882 -8111
rect 140943 -8145 140978 -8111
rect 143903 -8145 143938 -8111
rect 143999 -8145 144034 -8111
rect 144095 -8145 144130 -8111
rect 144191 -8145 144226 -8111
rect 144287 -8145 144322 -8111
rect 147247 -8145 147282 -8111
rect 147343 -8145 147378 -8111
rect 147439 -8145 147474 -8111
rect 147535 -8145 147570 -8111
rect 147631 -8145 147666 -8111
rect 150591 -8145 150626 -8111
rect 150687 -8145 150722 -8111
rect 150783 -8145 150818 -8111
rect 150879 -8145 150914 -8111
rect 150975 -8145 151010 -8111
rect 153935 -8145 153970 -8111
rect 154031 -8145 154066 -8111
rect 154127 -8145 154162 -8111
rect 154223 -8145 154258 -8111
rect 154319 -8145 154354 -8111
rect 157279 -8145 157314 -8111
rect 157375 -8145 157410 -8111
rect 157471 -8145 157506 -8111
rect 157567 -8145 157602 -8111
rect 157663 -8145 157698 -8111
rect 160623 -8145 160658 -8111
rect 160719 -8145 160754 -8111
rect 160815 -8145 160850 -8111
rect 160911 -8145 160946 -8111
rect 161007 -8145 161042 -8111
rect 163967 -8145 164002 -8111
rect 164063 -8145 164098 -8111
rect 164159 -8145 164194 -8111
rect 164255 -8145 164290 -8111
rect 164351 -8145 164386 -8111
rect 167311 -8145 167346 -8111
rect 167407 -8145 167442 -8111
rect 167503 -8145 167538 -8111
rect 167599 -8145 167634 -8111
rect 167695 -8145 167730 -8111
rect 170655 -8145 170690 -8111
rect 170751 -8145 170786 -8111
rect 170847 -8145 170882 -8111
rect 170943 -8145 170978 -8111
rect 171039 -8145 171074 -8111
rect 173999 -8145 174034 -8111
rect 174095 -8145 174130 -8111
rect 174191 -8145 174226 -8111
rect 174287 -8145 174322 -8111
rect 174383 -8145 174418 -8111
rect 177343 -8145 177378 -8111
rect 177439 -8145 177474 -8111
rect 177535 -8145 177570 -8111
rect 177631 -8145 177666 -8111
rect 177727 -8145 177762 -8111
rect 180687 -8145 180722 -8111
rect 180783 -8145 180818 -8111
rect 180879 -8145 180914 -8111
rect 180975 -8145 181010 -8111
rect 181071 -8145 181106 -8111
rect 184031 -8145 184066 -8111
rect 184127 -8145 184162 -8111
rect 184223 -8145 184258 -8111
rect 184319 -8145 184354 -8111
rect 184415 -8145 184450 -8111
rect 187375 -8145 187410 -8111
rect 187471 -8145 187506 -8111
rect 187567 -8145 187602 -8111
rect 187663 -8145 187698 -8111
rect 187759 -8145 187794 -8111
rect 190719 -8145 190754 -8111
rect 190815 -8145 190850 -8111
rect 190911 -8145 190946 -8111
rect 191007 -8145 191042 -8111
rect 191103 -8145 191138 -8111
rect 194063 -8145 194098 -8111
rect 194159 -8145 194194 -8111
rect 194255 -8145 194290 -8111
rect 194351 -8145 194386 -8111
rect 194447 -8145 194482 -8111
rect 197407 -8145 197442 -8111
rect 197503 -8145 197538 -8111
rect 197599 -8145 197634 -8111
rect 197695 -8145 197730 -8111
rect 197791 -8145 197826 -8111
rect 200751 -8145 200786 -8111
rect 200847 -8145 200882 -8111
rect 200943 -8145 200978 -8111
rect 201039 -8145 201074 -8111
rect 201135 -8145 201170 -8111
rect 204095 -8145 204130 -8111
rect 204191 -8145 204226 -8111
rect 204287 -8145 204322 -8111
rect 204383 -8145 204418 -8111
rect 204479 -8145 204514 -8111
rect 207439 -8145 207474 -8111
rect 207535 -8145 207570 -8111
rect 207631 -8145 207666 -8111
rect 207727 -8145 207762 -8111
rect 207823 -8145 207858 -8111
rect 210783 -8145 210818 -8111
rect 210879 -8145 210914 -8111
rect 210975 -8145 211010 -8111
rect 211071 -8145 211106 -8111
rect 211167 -8145 211202 -8111
rect 647 -8188 692 -8154
rect 743 -8188 788 -8154
rect 839 -8188 884 -8154
rect 935 -8188 980 -8154
rect 1031 -8188 1076 -8154
rect 1127 -8188 1172 -8154
rect 1223 -8188 1268 -8154
rect 3991 -8188 4036 -8154
rect 4087 -8188 4132 -8154
rect 4183 -8188 4228 -8154
rect 4279 -8188 4324 -8154
rect 4375 -8188 4420 -8154
rect 4471 -8188 4516 -8154
rect 4567 -8188 4612 -8154
rect 7336 -8188 7380 -8154
rect 7432 -8188 7476 -8154
rect 7528 -8188 7572 -8154
rect 7624 -8188 7668 -8154
rect 7720 -8188 7764 -8154
rect 7816 -8188 7860 -8154
rect 7912 -8188 7956 -8154
rect 10680 -8188 10724 -8154
rect 10776 -8188 10820 -8154
rect 10872 -8188 10916 -8154
rect 10968 -8188 11012 -8154
rect 11064 -8188 11108 -8154
rect 11160 -8188 11204 -8154
rect 11256 -8188 11300 -8154
rect 14025 -8188 14068 -8154
rect 14121 -8188 14164 -8154
rect 14217 -8188 14260 -8154
rect 14313 -8188 14356 -8154
rect 14409 -8188 14452 -8154
rect 14505 -8188 14548 -8154
rect 14601 -8188 14644 -8154
rect 17369 -8188 17412 -8154
rect 17465 -8188 17508 -8154
rect 17561 -8188 17604 -8154
rect 17657 -8188 17700 -8154
rect 17753 -8188 17796 -8154
rect 17849 -8188 17892 -8154
rect 17945 -8188 17988 -8154
rect 20713 -8188 20756 -8154
rect 20809 -8188 20852 -8154
rect 20905 -8188 20948 -8154
rect 21001 -8188 21044 -8154
rect 21097 -8188 21140 -8154
rect 21193 -8188 21236 -8154
rect 21289 -8188 21332 -8154
rect 24057 -8188 24100 -8154
rect 24153 -8188 24196 -8154
rect 24249 -8188 24292 -8154
rect 24345 -8188 24388 -8154
rect 24441 -8188 24484 -8154
rect 24537 -8188 24580 -8154
rect 24633 -8188 24676 -8154
rect 27402 -8188 27444 -8154
rect 27498 -8188 27540 -8154
rect 27594 -8188 27636 -8154
rect 27690 -8188 27732 -8154
rect 27786 -8188 27828 -8154
rect 27882 -8188 27924 -8154
rect 27978 -8188 28020 -8154
rect 30746 -8188 30788 -8154
rect 30842 -8188 30884 -8154
rect 30938 -8188 30980 -8154
rect 31034 -8188 31076 -8154
rect 31130 -8188 31172 -8154
rect 31226 -8188 31268 -8154
rect 31322 -8188 31364 -8154
rect 34090 -8188 34132 -8154
rect 34186 -8188 34228 -8154
rect 34282 -8188 34324 -8154
rect 34378 -8188 34420 -8154
rect 34474 -8188 34516 -8154
rect 34570 -8188 34612 -8154
rect 34666 -8188 34708 -8154
rect 37434 -8188 37476 -8154
rect 37530 -8188 37572 -8154
rect 37626 -8188 37668 -8154
rect 37722 -8188 37764 -8154
rect 37818 -8188 37860 -8154
rect 37914 -8188 37956 -8154
rect 38010 -8188 38052 -8154
rect 40778 -8188 40820 -8154
rect 40874 -8188 40916 -8154
rect 40970 -8188 41012 -8154
rect 41066 -8188 41108 -8154
rect 41162 -8188 41204 -8154
rect 41258 -8188 41300 -8154
rect 41354 -8188 41396 -8154
rect 44122 -8188 44164 -8154
rect 44218 -8188 44260 -8154
rect 44314 -8188 44356 -8154
rect 44410 -8188 44452 -8154
rect 44506 -8188 44548 -8154
rect 44602 -8188 44644 -8154
rect 44698 -8188 44740 -8154
rect 47466 -8188 47508 -8154
rect 47562 -8188 47604 -8154
rect 47658 -8188 47700 -8154
rect 47754 -8188 47796 -8154
rect 47850 -8188 47892 -8154
rect 47946 -8188 47988 -8154
rect 48042 -8188 48084 -8154
rect 50810 -8188 50852 -8154
rect 50906 -8188 50948 -8154
rect 51002 -8188 51044 -8154
rect 51098 -8188 51140 -8154
rect 51194 -8188 51236 -8154
rect 51290 -8188 51332 -8154
rect 51386 -8188 51428 -8154
rect 54155 -8188 54196 -8154
rect 54251 -8188 54292 -8154
rect 54347 -8188 54388 -8154
rect 54443 -8188 54484 -8154
rect 54539 -8188 54580 -8154
rect 54635 -8188 54676 -8154
rect 54731 -8188 54772 -8154
rect 57499 -8188 57540 -8154
rect 57595 -8188 57636 -8154
rect 57691 -8188 57732 -8154
rect 57787 -8188 57828 -8154
rect 57883 -8188 57924 -8154
rect 57979 -8188 58020 -8154
rect 58075 -8188 58116 -8154
rect 60843 -8188 60884 -8154
rect 60939 -8188 60980 -8154
rect 61035 -8188 61076 -8154
rect 61131 -8188 61172 -8154
rect 61227 -8188 61268 -8154
rect 61323 -8188 61364 -8154
rect 61419 -8188 61460 -8154
rect 64187 -8188 64228 -8154
rect 64283 -8188 64324 -8154
rect 64379 -8188 64420 -8154
rect 64475 -8188 64516 -8154
rect 64571 -8188 64612 -8154
rect 64667 -8188 64708 -8154
rect 64763 -8188 64804 -8154
rect 67531 -8188 67572 -8154
rect 67627 -8188 67668 -8154
rect 67723 -8188 67764 -8154
rect 67819 -8188 67860 -8154
rect 67915 -8188 67956 -8154
rect 68011 -8188 68052 -8154
rect 68107 -8188 68148 -8154
rect 70875 -8188 70916 -8154
rect 70971 -8188 71012 -8154
rect 71067 -8188 71108 -8154
rect 71163 -8188 71204 -8154
rect 71259 -8188 71300 -8154
rect 71355 -8188 71396 -8154
rect 71451 -8188 71492 -8154
rect 74219 -8188 74260 -8154
rect 74315 -8188 74356 -8154
rect 74411 -8188 74452 -8154
rect 74507 -8188 74548 -8154
rect 74603 -8188 74644 -8154
rect 74699 -8188 74740 -8154
rect 74795 -8188 74836 -8154
rect 77563 -8188 77604 -8154
rect 77659 -8188 77700 -8154
rect 77755 -8188 77796 -8154
rect 77851 -8188 77892 -8154
rect 77947 -8188 77988 -8154
rect 78043 -8188 78084 -8154
rect 78139 -8188 78180 -8154
rect 80907 -8188 80948 -8154
rect 81003 -8188 81044 -8154
rect 81099 -8188 81140 -8154
rect 81195 -8188 81236 -8154
rect 81291 -8188 81332 -8154
rect 81387 -8188 81428 -8154
rect 81483 -8188 81524 -8154
rect 84251 -8188 84292 -8154
rect 84347 -8188 84388 -8154
rect 84443 -8188 84484 -8154
rect 84539 -8188 84580 -8154
rect 84635 -8188 84676 -8154
rect 84731 -8188 84772 -8154
rect 84827 -8188 84868 -8154
rect 87595 -8188 87636 -8154
rect 87691 -8188 87732 -8154
rect 87787 -8188 87828 -8154
rect 87883 -8188 87924 -8154
rect 87979 -8188 88020 -8154
rect 88075 -8188 88116 -8154
rect 88171 -8188 88212 -8154
rect 90939 -8188 90980 -8154
rect 91035 -8188 91076 -8154
rect 91131 -8188 91172 -8154
rect 91227 -8188 91268 -8154
rect 91323 -8188 91364 -8154
rect 91419 -8188 91460 -8154
rect 91515 -8188 91556 -8154
rect 94283 -8188 94324 -8154
rect 94379 -8188 94420 -8154
rect 94475 -8188 94516 -8154
rect 94571 -8188 94612 -8154
rect 94667 -8188 94708 -8154
rect 94763 -8188 94804 -8154
rect 94859 -8188 94900 -8154
rect 97627 -8188 97668 -8154
rect 97723 -8188 97764 -8154
rect 97819 -8188 97860 -8154
rect 97915 -8188 97956 -8154
rect 98011 -8188 98052 -8154
rect 98107 -8188 98148 -8154
rect 98203 -8188 98244 -8154
rect 100971 -8188 101012 -8154
rect 101067 -8188 101108 -8154
rect 101163 -8188 101204 -8154
rect 101259 -8188 101300 -8154
rect 101355 -8188 101396 -8154
rect 101451 -8188 101492 -8154
rect 101547 -8188 101588 -8154
rect 104315 -8188 104356 -8154
rect 104411 -8188 104452 -8154
rect 104507 -8188 104548 -8154
rect 104603 -8188 104644 -8154
rect 104699 -8188 104740 -8154
rect 104795 -8188 104836 -8154
rect 104891 -8188 104932 -8154
rect 107665 -8188 107700 -8154
rect 107761 -8188 107796 -8154
rect 107857 -8188 107892 -8154
rect 107953 -8188 107988 -8154
rect 108049 -8188 108084 -8154
rect 108145 -8188 108180 -8154
rect 108241 -8188 108276 -8154
rect 111009 -8188 111044 -8154
rect 111105 -8188 111140 -8154
rect 111201 -8188 111236 -8154
rect 111297 -8188 111332 -8154
rect 111393 -8188 111428 -8154
rect 111489 -8188 111524 -8154
rect 111585 -8188 111620 -8154
rect 114353 -8188 114388 -8154
rect 114449 -8188 114484 -8154
rect 114545 -8188 114580 -8154
rect 114641 -8188 114676 -8154
rect 114737 -8188 114772 -8154
rect 114833 -8188 114868 -8154
rect 114929 -8188 114964 -8154
rect 117697 -8188 117732 -8154
rect 117793 -8188 117828 -8154
rect 117889 -8188 117924 -8154
rect 117985 -8188 118020 -8154
rect 118081 -8188 118116 -8154
rect 118177 -8188 118212 -8154
rect 118273 -8188 118308 -8154
rect 121041 -8188 121076 -8154
rect 121137 -8188 121172 -8154
rect 121233 -8188 121268 -8154
rect 121329 -8188 121364 -8154
rect 121425 -8188 121460 -8154
rect 121521 -8188 121556 -8154
rect 121617 -8188 121652 -8154
rect 124385 -8188 124420 -8154
rect 124481 -8188 124516 -8154
rect 124577 -8188 124612 -8154
rect 124673 -8188 124708 -8154
rect 124769 -8188 124804 -8154
rect 124865 -8188 124900 -8154
rect 124961 -8188 124996 -8154
rect 127729 -8188 127764 -8154
rect 127825 -8188 127860 -8154
rect 127921 -8188 127956 -8154
rect 128017 -8188 128052 -8154
rect 128113 -8188 128148 -8154
rect 128209 -8188 128244 -8154
rect 128305 -8188 128340 -8154
rect 131073 -8188 131108 -8154
rect 131169 -8188 131204 -8154
rect 131265 -8188 131300 -8154
rect 131361 -8188 131396 -8154
rect 131457 -8188 131492 -8154
rect 131553 -8188 131588 -8154
rect 131649 -8188 131684 -8154
rect 134417 -8188 134452 -8154
rect 134513 -8188 134548 -8154
rect 134609 -8188 134644 -8154
rect 134705 -8188 134740 -8154
rect 134801 -8188 134836 -8154
rect 134897 -8188 134932 -8154
rect 134993 -8188 135028 -8154
rect 137761 -8188 137796 -8154
rect 137857 -8188 137892 -8154
rect 137953 -8188 137988 -8154
rect 138049 -8188 138084 -8154
rect 138145 -8188 138180 -8154
rect 138241 -8188 138276 -8154
rect 138337 -8188 138372 -8154
rect 141105 -8188 141140 -8154
rect 141201 -8188 141236 -8154
rect 141297 -8188 141332 -8154
rect 141393 -8188 141428 -8154
rect 141489 -8188 141524 -8154
rect 141585 -8188 141620 -8154
rect 141681 -8188 141716 -8154
rect 144449 -8188 144484 -8154
rect 144545 -8188 144580 -8154
rect 144641 -8188 144676 -8154
rect 144737 -8188 144772 -8154
rect 144833 -8188 144868 -8154
rect 144929 -8188 144964 -8154
rect 145025 -8188 145060 -8154
rect 147793 -8188 147828 -8154
rect 147889 -8188 147924 -8154
rect 147985 -8188 148020 -8154
rect 148081 -8188 148116 -8154
rect 148177 -8188 148212 -8154
rect 148273 -8188 148308 -8154
rect 148369 -8188 148404 -8154
rect 151137 -8188 151172 -8154
rect 151233 -8188 151268 -8154
rect 151329 -8188 151364 -8154
rect 151425 -8188 151460 -8154
rect 151521 -8188 151556 -8154
rect 151617 -8188 151652 -8154
rect 151713 -8188 151748 -8154
rect 154481 -8188 154516 -8154
rect 154577 -8188 154612 -8154
rect 154673 -8188 154708 -8154
rect 154769 -8188 154804 -8154
rect 154865 -8188 154900 -8154
rect 154961 -8188 154996 -8154
rect 155057 -8188 155092 -8154
rect 157825 -8188 157860 -8154
rect 157921 -8188 157956 -8154
rect 158017 -8188 158052 -8154
rect 158113 -8188 158148 -8154
rect 158209 -8188 158244 -8154
rect 158305 -8188 158340 -8154
rect 158401 -8188 158436 -8154
rect 161169 -8188 161204 -8154
rect 161265 -8188 161300 -8154
rect 161361 -8188 161396 -8154
rect 161457 -8188 161492 -8154
rect 161553 -8188 161588 -8154
rect 161649 -8188 161684 -8154
rect 161745 -8188 161780 -8154
rect 164513 -8188 164548 -8154
rect 164609 -8188 164644 -8154
rect 164705 -8188 164740 -8154
rect 164801 -8188 164836 -8154
rect 164897 -8188 164932 -8154
rect 164993 -8188 165028 -8154
rect 165089 -8188 165124 -8154
rect 167857 -8188 167892 -8154
rect 167953 -8188 167988 -8154
rect 168049 -8188 168084 -8154
rect 168145 -8188 168180 -8154
rect 168241 -8188 168276 -8154
rect 168337 -8188 168372 -8154
rect 168433 -8188 168468 -8154
rect 171201 -8188 171236 -8154
rect 171297 -8188 171332 -8154
rect 171393 -8188 171428 -8154
rect 171489 -8188 171524 -8154
rect 171585 -8188 171620 -8154
rect 171681 -8188 171716 -8154
rect 171777 -8188 171812 -8154
rect 174545 -8188 174580 -8154
rect 174641 -8188 174676 -8154
rect 174737 -8188 174772 -8154
rect 174833 -8188 174868 -8154
rect 174929 -8188 174964 -8154
rect 175025 -8188 175060 -8154
rect 175121 -8188 175156 -8154
rect 177889 -8188 177924 -8154
rect 177985 -8188 178020 -8154
rect 178081 -8188 178116 -8154
rect 178177 -8188 178212 -8154
rect 178273 -8188 178308 -8154
rect 178369 -8188 178404 -8154
rect 178465 -8188 178500 -8154
rect 181233 -8188 181268 -8154
rect 181329 -8188 181364 -8154
rect 181425 -8188 181460 -8154
rect 181521 -8188 181556 -8154
rect 181617 -8188 181652 -8154
rect 181713 -8188 181748 -8154
rect 181809 -8188 181844 -8154
rect 184577 -8188 184612 -8154
rect 184673 -8188 184708 -8154
rect 184769 -8188 184804 -8154
rect 184865 -8188 184900 -8154
rect 184961 -8188 184996 -8154
rect 185057 -8188 185092 -8154
rect 185153 -8188 185188 -8154
rect 187921 -8188 187956 -8154
rect 188017 -8188 188052 -8154
rect 188113 -8188 188148 -8154
rect 188209 -8188 188244 -8154
rect 188305 -8188 188340 -8154
rect 188401 -8188 188436 -8154
rect 188497 -8188 188532 -8154
rect 191265 -8188 191300 -8154
rect 191361 -8188 191396 -8154
rect 191457 -8188 191492 -8154
rect 191553 -8188 191588 -8154
rect 191649 -8188 191684 -8154
rect 191745 -8188 191780 -8154
rect 191841 -8188 191876 -8154
rect 194609 -8188 194644 -8154
rect 194705 -8188 194740 -8154
rect 194801 -8188 194836 -8154
rect 194897 -8188 194932 -8154
rect 194993 -8188 195028 -8154
rect 195089 -8188 195124 -8154
rect 195185 -8188 195220 -8154
rect 197953 -8188 197988 -8154
rect 198049 -8188 198084 -8154
rect 198145 -8188 198180 -8154
rect 198241 -8188 198276 -8154
rect 198337 -8188 198372 -8154
rect 198433 -8188 198468 -8154
rect 198529 -8188 198564 -8154
rect 201297 -8188 201332 -8154
rect 201393 -8188 201428 -8154
rect 201489 -8188 201524 -8154
rect 201585 -8188 201620 -8154
rect 201681 -8188 201716 -8154
rect 201777 -8188 201812 -8154
rect 201873 -8188 201908 -8154
rect 204641 -8188 204676 -8154
rect 204737 -8188 204772 -8154
rect 204833 -8188 204868 -8154
rect 204929 -8188 204964 -8154
rect 205025 -8188 205060 -8154
rect 205121 -8188 205156 -8154
rect 205217 -8188 205252 -8154
rect 207985 -8188 208020 -8154
rect 208081 -8188 208116 -8154
rect 208177 -8188 208212 -8154
rect 208273 -8188 208308 -8154
rect 208369 -8188 208404 -8154
rect 208465 -8188 208500 -8154
rect 208561 -8188 208596 -8154
rect 211329 -8188 211364 -8154
rect 211425 -8188 211460 -8154
rect 211521 -8188 211556 -8154
rect 211617 -8188 211652 -8154
rect 211713 -8188 211748 -8154
rect 211809 -8188 211844 -8154
rect 211905 -8188 211940 -8154
rect 153 -8199 203 -8191
rect 203 -8207 214 -8199
rect 280 -8207 289 -8191
rect 314 -8199 359 -8191
rect 368 -8199 375 -8191
rect 303 -8207 323 -8199
rect 359 -8207 375 -8199
rect 94 -8241 139 -8207
rect 158 -8241 214 -8207
rect 238 -8241 289 -8207
rect 203 -8290 214 -8279
rect 158 -8324 214 -8290
rect 124 -8369 164 -8340
rect 203 -8369 214 -8363
rect 280 -8369 289 -8241
rect 314 -8241 375 -8207
rect 314 -8279 323 -8241
rect 368 -8279 375 -8241
rect 303 -8290 323 -8279
rect 359 -8290 375 -8279
rect 314 -8324 375 -8290
rect 314 -8340 323 -8324
rect 314 -8363 356 -8340
rect 368 -8363 375 -8324
rect 303 -8369 356 -8363
rect 359 -8369 375 -8363
rect 402 -8207 409 -8191
rect 470 -8199 520 -8191
rect 459 -8207 470 -8199
rect 402 -8241 453 -8207
rect 470 -8241 525 -8207
rect 1385 -8231 1430 -8197
rect 1481 -8231 1526 -8197
rect 1577 -8231 1622 -8197
rect 3497 -8199 3547 -8191
rect 3547 -8207 3558 -8199
rect 3624 -8207 3633 -8191
rect 3658 -8199 3703 -8191
rect 3712 -8199 3719 -8191
rect 3647 -8207 3667 -8199
rect 3703 -8207 3719 -8199
rect 402 -8369 409 -8241
rect 1178 -8250 1187 -8234
rect 1212 -8242 1262 -8234
rect 1201 -8250 1221 -8242
rect 459 -8290 470 -8279
rect 638 -8284 683 -8250
rect 710 -8284 755 -8250
rect 782 -8284 827 -8250
rect 926 -8284 971 -8250
rect 998 -8284 1115 -8250
rect 1142 -8284 1187 -8250
rect 470 -8324 515 -8290
rect 459 -8369 470 -8363
rect 124 -8374 483 -8369
rect 495 -8374 527 -8358
rect 1035 -8367 1080 -8333
rect 130 -8378 527 -8374
rect 130 -8403 531 -8378
rect 158 -8408 214 -8403
rect 146 -8431 161 -8416
rect 146 -8446 203 -8431
rect 146 -8457 214 -8446
rect 280 -8449 289 -8403
rect 314 -8408 375 -8403
rect 314 -8415 323 -8408
rect 314 -8431 331 -8415
rect 314 -8446 359 -8431
rect 368 -8446 375 -8408
rect 303 -8449 375 -8446
rect 402 -8449 409 -8403
rect 470 -8408 531 -8403
rect 280 -8454 297 -8449
rect 158 -8491 214 -8457
rect 236 -8465 297 -8454
rect 303 -8457 370 -8449
rect 247 -8499 297 -8465
rect 236 -8524 297 -8499
rect 176 -8571 297 -8524
rect 223 -8582 297 -8571
rect 314 -8491 370 -8457
rect 392 -8465 448 -8454
rect 459 -8457 470 -8446
rect 495 -8457 531 -8408
rect 1060 -8412 1114 -8383
rect 1178 -8412 1187 -8284
rect 1212 -8284 1257 -8250
rect 1739 -8274 1784 -8240
rect 1835 -8274 1880 -8240
rect 1931 -8274 1976 -8240
rect 3438 -8241 3483 -8207
rect 3502 -8241 3558 -8207
rect 3582 -8241 3633 -8207
rect 1212 -8322 1221 -8284
rect 1401 -8285 1451 -8277
rect 1562 -8285 1612 -8277
rect 1451 -8293 1462 -8285
rect 1551 -8293 1562 -8285
rect 1201 -8333 1221 -8322
rect 1378 -8327 1495 -8293
rect 1562 -8327 1607 -8293
rect 2093 -8317 2138 -8283
rect 2189 -8317 2234 -8283
rect 2285 -8317 2330 -8283
rect 2381 -8317 2426 -8283
rect 2477 -8317 2522 -8283
rect 3547 -8290 3558 -8279
rect 1755 -8328 1805 -8320
rect 1916 -8328 1966 -8320
rect 3502 -8324 3558 -8290
rect 1212 -8367 1257 -8333
rect 1805 -8336 1816 -8328
rect 1905 -8336 1916 -8328
rect 1212 -8406 1221 -8367
rect 1451 -8376 1462 -8365
rect 1551 -8376 1562 -8365
rect 1732 -8370 1849 -8336
rect 1916 -8370 1961 -8336
rect 2641 -8360 2686 -8326
rect 2737 -8360 2782 -8326
rect 2833 -8360 2878 -8326
rect 2929 -8360 2974 -8326
rect 3025 -8360 3070 -8326
rect 3121 -8360 3166 -8326
rect 3217 -8360 3262 -8326
rect 2145 -8371 2195 -8363
rect 1201 -8412 1221 -8406
rect 549 -8446 581 -8412
rect 634 -8417 1221 -8412
rect 1233 -8417 1269 -8401
rect 1406 -8410 1462 -8376
rect 1562 -8410 1607 -8376
rect 2195 -8379 2206 -8371
rect 2272 -8379 2281 -8363
rect 2306 -8371 2351 -8363
rect 2360 -8371 2367 -8363
rect 2295 -8379 2315 -8371
rect 2351 -8379 2367 -8371
rect 634 -8421 1269 -8417
rect 1805 -8419 1816 -8408
rect 1905 -8419 1916 -8408
rect 2086 -8413 2131 -8379
rect 2150 -8413 2206 -8379
rect 2230 -8413 2281 -8379
rect 634 -8446 1278 -8421
rect 314 -8582 331 -8491
rect 403 -8499 448 -8465
rect 470 -8480 531 -8457
rect 688 -8472 745 -8458
rect 470 -8491 527 -8480
rect 495 -8499 527 -8491
rect 223 -8605 331 -8582
rect 236 -8655 297 -8605
rect 314 -8637 331 -8605
rect 392 -8537 449 -8499
rect 470 -8507 520 -8499
rect 688 -8500 756 -8472
rect 700 -8517 756 -8500
rect 822 -8534 831 -8446
rect 856 -8472 901 -8450
rect 845 -8483 912 -8472
rect 856 -8517 912 -8483
rect 926 -8492 935 -8446
rect 1023 -8458 1027 -8446
rect 1035 -8451 1080 -8446
rect 1012 -8497 1023 -8458
rect 957 -8500 1023 -8497
rect 1034 -8500 1101 -8474
rect 1178 -8492 1187 -8446
rect 1212 -8451 1278 -8446
rect 1212 -8458 1221 -8451
rect 1233 -8458 1278 -8451
rect 1414 -8455 1448 -8426
rect 1451 -8455 1462 -8449
rect 1551 -8455 1562 -8449
rect 1212 -8489 1278 -8458
rect 1287 -8489 1323 -8455
rect 1394 -8460 1575 -8455
rect 1587 -8460 1619 -8444
rect 1760 -8453 1816 -8419
rect 1916 -8453 1961 -8419
rect 1394 -8464 1619 -8460
rect 2195 -8462 2206 -8451
rect 1394 -8489 1634 -8464
rect 1178 -8497 1200 -8492
rect 957 -8508 1012 -8500
rect 392 -8613 453 -8537
rect 465 -8587 487 -8571
rect 465 -8613 520 -8587
rect 533 -8613 536 -8571
rect 567 -8613 570 -8542
rect 392 -8655 581 -8613
rect 120 -8823 581 -8655
rect 676 -8666 721 -8632
rect 676 -8716 721 -8700
rect 725 -8716 753 -8536
rect 856 -8568 865 -8517
rect 968 -8542 1012 -8508
rect 1034 -8534 1091 -8500
rect 1134 -8508 1200 -8497
rect 1201 -8500 1278 -8489
rect 1406 -8494 1462 -8489
rect 1562 -8494 1634 -8489
rect 1034 -8542 1054 -8534
rect 1145 -8542 1200 -8508
rect 759 -8716 787 -8570
rect 799 -8606 810 -8595
rect 795 -8637 810 -8606
rect 795 -8648 804 -8637
rect 792 -8690 810 -8648
rect 829 -8674 838 -8640
rect 841 -8674 852 -8637
rect 857 -8674 902 -8654
rect 829 -8688 902 -8674
rect 795 -8708 804 -8690
rect 795 -8716 823 -8708
rect 829 -8716 857 -8688
rect 956 -8716 1012 -8542
rect 1134 -8543 1200 -8542
rect 1074 -8590 1200 -8543
rect 1121 -8624 1200 -8590
rect 1134 -8660 1200 -8624
rect 1212 -8523 1278 -8500
rect 1212 -8542 1269 -8523
rect 1212 -8550 1262 -8542
rect 1212 -8660 1234 -8550
rect 1271 -8660 1278 -8523
rect 1394 -8517 1409 -8502
rect 1394 -8532 1451 -8517
rect 1305 -8660 1312 -8535
rect 1394 -8543 1462 -8532
rect 1406 -8577 1462 -8543
rect 1484 -8551 1540 -8540
rect 1551 -8543 1562 -8532
rect 1587 -8543 1634 -8494
rect 1768 -8498 1802 -8469
rect 1805 -8498 1816 -8492
rect 1905 -8498 1916 -8492
rect 1641 -8532 1673 -8498
rect 1748 -8503 1929 -8498
rect 1941 -8503 1973 -8487
rect 2150 -8496 2206 -8462
rect 1748 -8507 1973 -8503
rect 1748 -8532 1988 -8507
rect 1760 -8537 1816 -8532
rect 1916 -8537 1988 -8532
rect 1495 -8585 1540 -8551
rect 1562 -8566 1634 -8543
rect 1562 -8577 1619 -8566
rect 1587 -8585 1619 -8577
rect 1484 -8593 1541 -8585
rect 1562 -8593 1612 -8585
rect 1484 -8610 1556 -8593
rect 1424 -8657 1556 -8610
rect 1134 -8702 1337 -8660
rect 1471 -8691 1556 -8657
rect 641 -8722 1012 -8716
rect 641 -8731 825 -8722
rect 656 -8734 823 -8731
rect 656 -8768 678 -8734
rect 725 -8768 753 -8734
rect 759 -8768 823 -8734
rect 829 -8756 1012 -8722
rect 829 -8768 857 -8756
rect 934 -8768 1012 -8756
rect 1022 -8768 1337 -8702
rect 1484 -8703 1556 -8691
rect 1557 -8703 1590 -8593
rect 1625 -8703 1634 -8566
rect 1748 -8560 1763 -8545
rect 1748 -8575 1805 -8560
rect 1659 -8703 1668 -8578
rect 1748 -8586 1816 -8575
rect 1760 -8620 1816 -8586
rect 1838 -8594 1894 -8583
rect 1905 -8586 1916 -8575
rect 1941 -8586 1988 -8537
rect 2116 -8541 2156 -8512
rect 2195 -8541 2206 -8535
rect 2272 -8541 2281 -8413
rect 2306 -8413 2367 -8379
rect 2306 -8451 2315 -8413
rect 2360 -8451 2367 -8413
rect 2295 -8462 2315 -8451
rect 2351 -8462 2367 -8451
rect 2306 -8496 2367 -8462
rect 2306 -8512 2315 -8496
rect 2306 -8535 2348 -8512
rect 2360 -8535 2367 -8496
rect 2295 -8541 2348 -8535
rect 2351 -8541 2367 -8535
rect 2394 -8379 2401 -8363
rect 2462 -8371 2512 -8363
rect 2451 -8379 2462 -8371
rect 3547 -8374 3558 -8363
rect 2394 -8413 2445 -8379
rect 2462 -8413 2517 -8379
rect 2394 -8541 2401 -8413
rect 3172 -8422 3181 -8406
rect 3206 -8414 3256 -8406
rect 3502 -8408 3558 -8374
rect 3195 -8422 3215 -8414
rect 2451 -8462 2462 -8451
rect 2632 -8456 2677 -8422
rect 2704 -8456 2749 -8422
rect 2776 -8456 2821 -8422
rect 2920 -8456 2965 -8422
rect 2992 -8456 3109 -8422
rect 3136 -8456 3181 -8422
rect 2462 -8496 2507 -8462
rect 2451 -8541 2462 -8535
rect 1995 -8575 2027 -8541
rect 2116 -8546 2475 -8541
rect 2489 -8546 2519 -8530
rect 3029 -8539 3074 -8505
rect 2122 -8550 2519 -8546
rect 2122 -8575 2523 -8550
rect 2150 -8580 2206 -8575
rect 1849 -8628 1894 -8594
rect 1916 -8609 1988 -8586
rect 1916 -8620 1973 -8609
rect 1941 -8628 1973 -8620
rect 1838 -8636 1895 -8628
rect 1916 -8636 1966 -8628
rect 1838 -8653 1910 -8636
rect 1778 -8700 1910 -8653
rect 1484 -8745 1691 -8703
rect 1825 -8734 1910 -8700
rect 94 -8863 139 -8829
rect 146 -8831 228 -8823
rect 314 -8829 345 -8823
rect 166 -8863 211 -8831
rect 238 -8863 283 -8829
rect 310 -8863 355 -8829
rect 370 -8831 480 -8823
rect 483 -8831 581 -8823
rect 620 -8816 1337 -8768
rect 1372 -8816 1691 -8745
rect 1838 -8746 1910 -8734
rect 1911 -8746 1944 -8636
rect 1979 -8746 1988 -8609
rect 2138 -8603 2153 -8588
rect 2138 -8618 2195 -8603
rect 2013 -8746 2022 -8621
rect 2138 -8629 2206 -8618
rect 2272 -8621 2281 -8575
rect 2306 -8580 2367 -8575
rect 2306 -8587 2315 -8580
rect 2306 -8603 2323 -8587
rect 2306 -8618 2351 -8603
rect 2360 -8618 2367 -8580
rect 2295 -8621 2367 -8618
rect 2394 -8621 2401 -8575
rect 2462 -8580 2523 -8575
rect 2272 -8626 2289 -8621
rect 2150 -8663 2206 -8629
rect 2228 -8637 2289 -8626
rect 2295 -8629 2362 -8621
rect 2239 -8671 2289 -8637
rect 2228 -8696 2289 -8671
rect 2168 -8743 2289 -8696
rect 1838 -8788 2045 -8746
rect 2215 -8754 2289 -8743
rect 2306 -8663 2362 -8629
rect 2384 -8637 2440 -8626
rect 2451 -8629 2462 -8618
rect 2489 -8629 2523 -8580
rect 3054 -8584 3108 -8555
rect 3172 -8584 3181 -8456
rect 3206 -8456 3251 -8422
rect 3206 -8494 3215 -8456
rect 3547 -8457 3558 -8446
rect 3502 -8491 3558 -8457
rect 3195 -8505 3215 -8494
rect 3206 -8539 3251 -8505
rect 3206 -8578 3215 -8539
rect 3359 -8565 3464 -8499
rect 3497 -8507 3547 -8499
rect 3624 -8507 3633 -8241
rect 3658 -8241 3719 -8207
rect 3658 -8279 3667 -8241
rect 3712 -8279 3719 -8241
rect 3647 -8290 3667 -8279
rect 3703 -8290 3719 -8279
rect 3658 -8324 3719 -8290
rect 3658 -8363 3667 -8324
rect 3712 -8363 3719 -8324
rect 3647 -8374 3667 -8363
rect 3703 -8374 3719 -8363
rect 3658 -8408 3719 -8374
rect 3658 -8446 3667 -8408
rect 3712 -8446 3719 -8408
rect 3647 -8457 3667 -8446
rect 3703 -8457 3719 -8446
rect 3658 -8483 3719 -8457
rect 3647 -8491 3719 -8483
rect 3647 -8499 3667 -8491
rect 3647 -8507 3703 -8499
rect 3647 -8525 3667 -8507
rect 3658 -8541 3667 -8525
rect 3195 -8584 3215 -8578
rect 2543 -8618 2573 -8584
rect 2628 -8589 3215 -8584
rect 2628 -8618 3251 -8589
rect 3567 -8605 3612 -8571
rect 2306 -8754 2323 -8663
rect 2395 -8671 2440 -8637
rect 2462 -8652 2523 -8629
rect 2682 -8644 2739 -8630
rect 2462 -8663 2519 -8652
rect 2489 -8671 2519 -8663
rect 2215 -8777 2323 -8754
rect 456 -8833 539 -8831
rect 483 -8866 539 -8833
rect 620 -8843 1691 -8816
rect 620 -8866 1337 -8843
rect 622 -8874 642 -8866
rect 646 -8878 699 -8866
rect 819 -8874 852 -8866
rect 1019 -8870 1116 -8866
rect 1019 -8872 1126 -8870
rect 752 -8878 852 -8874
rect 408 -8879 442 -8878
rect 247 -8895 319 -8891
rect 398 -8895 458 -8891
rect 70 -8929 530 -8925
rect 70 -8939 242 -8929
rect 278 -8939 378 -8929
rect 389 -8939 434 -8929
rect 70 -8959 435 -8939
rect 485 -8959 530 -8929
rect 540 -8959 561 -8925
rect 574 -8992 595 -8891
rect 834 -8895 852 -8878
rect 953 -8906 998 -8872
rect 1019 -8878 1142 -8872
rect 1025 -8906 1070 -8878
rect 1097 -8906 1142 -8878
rect 1178 -8920 1200 -8866
rect 1212 -8878 1337 -8866
rect 1372 -8859 1691 -8843
rect 1726 -8859 2045 -8788
rect 2228 -8827 2289 -8777
rect 2306 -8809 2323 -8777
rect 2384 -8709 2441 -8671
rect 2462 -8679 2512 -8671
rect 2682 -8672 2750 -8644
rect 2694 -8689 2750 -8672
rect 2816 -8706 2825 -8618
rect 2850 -8644 2895 -8622
rect 2839 -8655 2906 -8644
rect 2850 -8689 2906 -8655
rect 2920 -8664 2929 -8618
rect 3017 -8630 3021 -8618
rect 3029 -8623 3074 -8618
rect 3006 -8669 3017 -8630
rect 2951 -8672 3017 -8669
rect 3028 -8672 3095 -8646
rect 3172 -8664 3181 -8618
rect 3206 -8623 3251 -8618
rect 3206 -8630 3215 -8623
rect 3206 -8661 3228 -8630
rect 3624 -8632 3628 -8555
rect 3658 -8637 3662 -8541
rect 3172 -8669 3194 -8664
rect 2951 -8680 3006 -8672
rect 2384 -8785 2445 -8709
rect 2457 -8759 2479 -8743
rect 2457 -8785 2512 -8759
rect 2527 -8785 2528 -8743
rect 2561 -8785 2562 -8714
rect 2384 -8827 2573 -8785
rect 1212 -8886 1295 -8878
rect 1221 -8909 1295 -8886
rect 1372 -8886 2045 -8859
rect 1372 -8909 1691 -8886
rect 1398 -8915 1476 -8909
rect 1378 -8921 1495 -8915
rect 1034 -8960 1038 -8957
rect 616 -8978 732 -8968
rect 743 -8978 934 -8968
rect 935 -8978 980 -8968
rect 616 -8986 981 -8978
rect 1031 -8986 1172 -8968
rect 616 -9002 1191 -8986
rect 1223 -9002 1299 -8968
rect 1312 -8976 1333 -8934
rect 1378 -8949 1423 -8921
rect 1450 -8949 1495 -8921
rect 1523 -8963 1556 -8909
rect 1557 -8921 1691 -8909
rect 1557 -8929 1649 -8921
rect 1575 -8952 1649 -8929
rect 1726 -8952 2045 -8886
rect 2071 -8921 2083 -8902
rect 2112 -8921 2573 -8827
rect 2670 -8838 2715 -8804
rect 2670 -8888 2715 -8872
rect 2719 -8888 2747 -8708
rect 2850 -8740 2859 -8689
rect 2962 -8714 3006 -8680
rect 3028 -8706 3085 -8672
rect 3128 -8680 3194 -8669
rect 3195 -8672 3228 -8661
rect 3028 -8714 3048 -8706
rect 3139 -8714 3194 -8680
rect 2753 -8888 2781 -8742
rect 2793 -8778 2804 -8767
rect 2789 -8809 2804 -8778
rect 2789 -8820 2798 -8809
rect 2786 -8862 2804 -8820
rect 2823 -8846 2832 -8812
rect 2835 -8846 2846 -8809
rect 2851 -8846 2896 -8826
rect 2823 -8860 2896 -8846
rect 2789 -8880 2798 -8862
rect 2789 -8888 2817 -8880
rect 2823 -8888 2851 -8860
rect 2950 -8888 3006 -8714
rect 3128 -8715 3194 -8714
rect 3068 -8762 3194 -8715
rect 3115 -8796 3194 -8762
rect 3128 -8832 3194 -8796
rect 3206 -8706 3251 -8672
rect 3689 -8673 3700 -8525
rect 3712 -8541 3719 -8491
rect 3746 -8207 3753 -8191
rect 3814 -8199 3864 -8191
rect 3803 -8207 3814 -8199
rect 3746 -8241 3797 -8207
rect 3814 -8241 3869 -8207
rect 4729 -8231 4774 -8197
rect 4825 -8231 4870 -8197
rect 4921 -8231 4966 -8197
rect 6892 -8207 6902 -8199
rect 6969 -8207 6977 -8191
rect 6992 -8207 7002 -8199
rect 7003 -8207 7011 -8191
rect 7057 -8199 7063 -8191
rect 3746 -8507 3753 -8241
rect 4522 -8250 4531 -8234
rect 4556 -8242 4606 -8234
rect 4545 -8250 4565 -8242
rect 3803 -8290 3814 -8279
rect 3982 -8284 4027 -8250
rect 4054 -8284 4099 -8250
rect 4126 -8284 4171 -8250
rect 4270 -8284 4315 -8250
rect 4342 -8284 4459 -8250
rect 4486 -8284 4531 -8250
rect 3814 -8324 3859 -8290
rect 3803 -8374 3814 -8363
rect 4379 -8367 4424 -8333
rect 3814 -8408 3859 -8374
rect 3803 -8457 3814 -8446
rect 3814 -8491 3859 -8457
rect 4089 -8483 4100 -8472
rect 3814 -8507 3864 -8499
rect 4044 -8517 4100 -8483
rect 4166 -8534 4175 -8416
rect 4200 -8472 4209 -8450
rect 4189 -8483 4209 -8472
rect 4236 -8472 4245 -8450
rect 4236 -8483 4256 -8472
rect 4200 -8517 4256 -8483
rect 4200 -8568 4209 -8517
rect 4236 -8568 4245 -8517
rect 4270 -8534 4279 -8417
rect 4367 -8458 4371 -8417
rect 4379 -8451 4424 -8417
rect 4379 -8534 4424 -8500
rect 4522 -8534 4531 -8284
rect 4556 -8284 4601 -8250
rect 5083 -8274 5128 -8240
rect 5179 -8274 5224 -8240
rect 5275 -8274 5320 -8240
rect 6783 -8241 6827 -8207
rect 6847 -8241 6902 -8207
rect 6927 -8241 6977 -8207
rect 4556 -8322 4565 -8284
rect 4745 -8285 4795 -8277
rect 4906 -8285 4956 -8277
rect 4795 -8293 4806 -8285
rect 4895 -8293 4906 -8285
rect 4545 -8333 4565 -8322
rect 4722 -8327 4839 -8293
rect 4906 -8327 4951 -8293
rect 5437 -8317 5482 -8283
rect 5533 -8317 5578 -8283
rect 5629 -8317 5674 -8283
rect 5725 -8317 5770 -8283
rect 5821 -8317 5866 -8283
rect 5099 -8328 5149 -8320
rect 5260 -8328 5310 -8320
rect 6847 -8324 6891 -8290
rect 6892 -8324 6902 -8279
rect 4556 -8367 4601 -8333
rect 5149 -8336 5160 -8328
rect 5249 -8336 5260 -8328
rect 4556 -8406 4565 -8367
rect 4795 -8376 4806 -8365
rect 4895 -8376 4906 -8365
rect 5076 -8370 5193 -8336
rect 5260 -8370 5305 -8336
rect 5985 -8360 6030 -8326
rect 6081 -8360 6126 -8326
rect 6177 -8360 6222 -8326
rect 6273 -8360 6318 -8326
rect 6369 -8360 6414 -8326
rect 6465 -8360 6510 -8326
rect 6561 -8360 6606 -8326
rect 5489 -8371 5539 -8363
rect 4545 -8417 4565 -8406
rect 4750 -8410 4806 -8376
rect 4906 -8410 4951 -8376
rect 5539 -8379 5550 -8371
rect 5616 -8379 5625 -8363
rect 5650 -8371 5695 -8363
rect 5704 -8371 5711 -8363
rect 5639 -8379 5659 -8371
rect 5695 -8379 5711 -8371
rect 4556 -8451 4601 -8417
rect 5149 -8419 5160 -8408
rect 5249 -8419 5260 -8408
rect 5430 -8413 5475 -8379
rect 5494 -8413 5550 -8379
rect 5574 -8413 5625 -8379
rect 4556 -8489 4565 -8451
rect 4795 -8460 4806 -8449
rect 4895 -8460 4906 -8449
rect 5104 -8453 5160 -8419
rect 5260 -8453 5305 -8419
rect 4545 -8500 4565 -8489
rect 4750 -8494 4806 -8460
rect 4906 -8494 4951 -8460
rect 5539 -8462 5550 -8451
rect 4556 -8534 4601 -8500
rect 5149 -8503 5160 -8492
rect 5249 -8503 5260 -8492
rect 5494 -8496 5550 -8462
rect 4556 -8542 4565 -8534
rect 4556 -8550 4606 -8542
rect 4795 -8543 4806 -8532
rect 4895 -8543 4906 -8532
rect 5104 -8537 5160 -8503
rect 5260 -8537 5305 -8503
rect 4556 -8568 4565 -8550
rect 3497 -8681 3547 -8673
rect 3547 -8689 3558 -8681
rect 3206 -8714 3228 -8706
rect 3206 -8722 3256 -8714
rect 3206 -8819 3228 -8722
rect 3502 -8723 3558 -8689
rect 3689 -8741 3705 -8673
rect 3730 -8707 3739 -8639
rect 3775 -8671 3784 -8603
rect 3809 -8637 3818 -8571
rect 3819 -8621 3864 -8587
rect 4020 -8666 4065 -8632
rect 3800 -8681 3850 -8673
rect 3789 -8689 3800 -8681
rect 3800 -8723 3845 -8689
rect 4020 -8734 4065 -8700
rect 3689 -8753 3700 -8741
rect 4069 -8750 4078 -8616
rect 3464 -8819 3861 -8753
rect 4103 -8784 4112 -8590
rect 4143 -8606 4154 -8595
rect 4139 -8637 4154 -8606
rect 4465 -8624 4510 -8590
rect 4043 -8819 4054 -8808
rect 3200 -8832 3228 -8819
rect 3128 -8874 3228 -8832
rect 3262 -8874 3861 -8819
rect 3998 -8853 4054 -8819
rect 4139 -8820 4148 -8637
rect 4173 -8823 4182 -8640
rect 2635 -8894 3006 -8888
rect 2635 -8903 2819 -8894
rect 2071 -8929 2573 -8921
rect 1752 -8958 1830 -8952
rect 1732 -8964 1849 -8958
rect 1384 -9003 1388 -9000
rect 1305 -9029 1333 -9021
rect 1354 -9029 1526 -9011
rect 1305 -9036 1545 -9029
rect 1331 -9045 1545 -9036
rect 1577 -9045 1653 -9011
rect 1666 -9019 1687 -8977
rect 1732 -8992 1777 -8964
rect 1804 -8992 1849 -8964
rect 1877 -9006 1910 -8952
rect 1911 -8964 2045 -8952
rect 1911 -8972 2003 -8964
rect 1929 -8995 2003 -8972
rect 2112 -8995 2573 -8929
rect 2650 -8906 2817 -8903
rect 2650 -8940 2672 -8906
rect 2719 -8940 2747 -8906
rect 2753 -8940 2817 -8906
rect 2823 -8928 3006 -8894
rect 2823 -8940 2851 -8928
rect 2928 -8940 3006 -8928
rect 3016 -8877 3861 -8874
rect 3016 -8940 3289 -8877
rect 3464 -8899 3861 -8877
rect 732 -9076 774 -9052
rect 934 -9076 981 -9052
rect 1331 -9071 1373 -9045
rect 1738 -9046 1742 -9043
rect 1659 -9072 1687 -9064
rect 1708 -9072 1880 -9054
rect 1659 -9079 1899 -9072
rect 1685 -9088 1899 -9079
rect 1931 -9088 1976 -9054
rect 1986 -9069 2007 -9054
rect 2020 -9062 2041 -9020
rect 2086 -9035 2131 -9001
rect 2138 -9003 2220 -8995
rect 2306 -9001 2337 -8995
rect 2158 -9035 2203 -9003
rect 2230 -9035 2275 -9001
rect 2302 -9035 2347 -9001
rect 2362 -9003 2472 -8995
rect 2477 -9003 2573 -8995
rect 2448 -9005 2531 -9003
rect 2477 -9038 2531 -9005
rect 2614 -9038 3289 -8940
rect 3388 -8925 3861 -8899
rect 4185 -8904 4196 -8637
rect 4522 -8640 4526 -8570
rect 4201 -8688 4246 -8654
rect 4556 -8674 4560 -8568
rect 4750 -8577 4806 -8543
rect 4906 -8577 4951 -8543
rect 5539 -8546 5550 -8535
rect 4745 -8593 4795 -8585
rect 4906 -8593 4956 -8585
rect 5149 -8586 5160 -8575
rect 5249 -8586 5260 -8575
rect 5494 -8580 5550 -8546
rect 4201 -8756 4246 -8722
rect 4253 -8823 4262 -8688
rect 4815 -8691 4860 -8657
rect 4867 -8718 4876 -8641
rect 4287 -8808 4296 -8720
rect 4399 -8728 4449 -8720
rect 4560 -8728 4610 -8724
rect 4449 -8736 4460 -8728
rect 4404 -8770 4460 -8736
rect 4549 -8740 4560 -8729
rect 4560 -8774 4605 -8740
rect 4901 -8752 4910 -8607
rect 5104 -8620 5160 -8586
rect 5260 -8620 5305 -8586
rect 5099 -8636 5149 -8628
rect 5260 -8636 5310 -8628
rect 5539 -8629 5550 -8618
rect 5169 -8734 5214 -8700
rect 5221 -8761 5230 -8684
rect 4749 -8771 4799 -8763
rect 4910 -8771 4960 -8763
rect 4799 -8779 4810 -8771
rect 4899 -8779 4910 -8771
rect 4285 -8819 4296 -8808
rect 4754 -8813 4810 -8779
rect 4910 -8813 4955 -8779
rect 5255 -8795 5264 -8650
rect 5494 -8663 5550 -8629
rect 5489 -8679 5539 -8671
rect 5616 -8679 5625 -8413
rect 5650 -8413 5711 -8379
rect 5650 -8451 5659 -8413
rect 5704 -8451 5711 -8413
rect 5639 -8462 5659 -8451
rect 5695 -8462 5711 -8451
rect 5650 -8496 5711 -8462
rect 5650 -8535 5659 -8496
rect 5704 -8535 5711 -8496
rect 5639 -8546 5659 -8535
rect 5695 -8546 5711 -8535
rect 5650 -8580 5711 -8546
rect 5650 -8618 5659 -8580
rect 5704 -8618 5711 -8580
rect 5639 -8629 5659 -8618
rect 5695 -8629 5711 -8618
rect 5650 -8655 5711 -8629
rect 5639 -8663 5711 -8655
rect 5639 -8671 5659 -8663
rect 5639 -8679 5695 -8671
rect 5639 -8697 5659 -8679
rect 5650 -8713 5659 -8697
rect 5559 -8777 5604 -8743
rect 5616 -8804 5620 -8727
rect 5103 -8814 5153 -8806
rect 5264 -8814 5314 -8806
rect 5650 -8809 5654 -8713
rect 4287 -8853 4341 -8819
rect 4449 -8836 4460 -8825
rect 4549 -8832 4560 -8821
rect 5153 -8822 5164 -8814
rect 5253 -8822 5264 -8814
rect 4404 -8870 4460 -8836
rect 4560 -8866 4605 -8832
rect 5108 -8856 5164 -8822
rect 5264 -8856 5309 -8822
rect 5681 -8845 5692 -8697
rect 5704 -8713 5711 -8663
rect 5738 -8379 5745 -8363
rect 5806 -8371 5856 -8363
rect 5795 -8379 5806 -8371
rect 5738 -8413 5789 -8379
rect 5806 -8413 5861 -8379
rect 5738 -8679 5745 -8413
rect 6516 -8422 6525 -8406
rect 6550 -8414 6600 -8406
rect 6847 -8408 6891 -8374
rect 6892 -8408 6902 -8363
rect 6539 -8422 6559 -8414
rect 5795 -8462 5806 -8451
rect 5976 -8456 6021 -8422
rect 6048 -8456 6093 -8422
rect 6120 -8456 6165 -8422
rect 6264 -8456 6309 -8422
rect 6336 -8456 6453 -8422
rect 6480 -8456 6525 -8422
rect 5806 -8496 5851 -8462
rect 5795 -8546 5806 -8535
rect 6373 -8539 6418 -8505
rect 5806 -8580 5851 -8546
rect 5795 -8629 5806 -8618
rect 5806 -8663 5851 -8629
rect 6083 -8655 6094 -8644
rect 5806 -8679 5856 -8671
rect 6038 -8689 6094 -8655
rect 6160 -8706 6169 -8588
rect 6194 -8644 6203 -8622
rect 6183 -8655 6203 -8644
rect 6230 -8644 6239 -8622
rect 6230 -8655 6250 -8644
rect 6194 -8689 6250 -8655
rect 6194 -8740 6203 -8689
rect 6230 -8740 6239 -8689
rect 6264 -8706 6273 -8589
rect 6361 -8630 6365 -8589
rect 6373 -8623 6418 -8589
rect 6373 -8706 6418 -8672
rect 6516 -8706 6525 -8456
rect 6550 -8456 6595 -8422
rect 6550 -8494 6559 -8456
rect 6847 -8491 6891 -8457
rect 6892 -8491 6902 -8446
rect 6539 -8505 6559 -8494
rect 6550 -8539 6595 -8505
rect 6550 -8578 6559 -8539
rect 6703 -8565 6809 -8499
rect 6969 -8507 6977 -8241
rect 7003 -8241 7047 -8207
rect 7048 -8241 7063 -8199
rect 6992 -8290 7002 -8279
rect 7003 -8290 7011 -8241
rect 7057 -8279 7063 -8241
rect 7003 -8324 7047 -8290
rect 7048 -8324 7063 -8279
rect 6992 -8374 7002 -8363
rect 7003 -8374 7011 -8324
rect 7057 -8363 7063 -8324
rect 7003 -8408 7047 -8374
rect 7048 -8408 7063 -8363
rect 6992 -8457 7002 -8446
rect 7003 -8457 7011 -8408
rect 7057 -8446 7063 -8408
rect 6992 -8525 7002 -8483
rect 7003 -8491 7047 -8457
rect 7048 -8491 7063 -8446
rect 7003 -8541 7011 -8491
rect 6539 -8589 6559 -8578
rect 6550 -8623 6595 -8589
rect 6912 -8605 6956 -8571
rect 6550 -8661 6559 -8623
rect 6969 -8632 6972 -8555
rect 7003 -8637 7006 -8541
rect 6539 -8672 6559 -8661
rect 6550 -8706 6595 -8672
rect 7034 -8673 7044 -8525
rect 7057 -8541 7063 -8491
rect 7091 -8207 7097 -8191
rect 7148 -8207 7158 -8199
rect 7091 -8241 7141 -8207
rect 7159 -8241 7213 -8207
rect 8074 -8231 8118 -8197
rect 8170 -8231 8214 -8197
rect 8266 -8231 8310 -8197
rect 10236 -8207 10246 -8199
rect 10313 -8207 10321 -8191
rect 10336 -8207 10346 -8199
rect 10347 -8207 10355 -8191
rect 10401 -8199 10407 -8191
rect 7091 -8507 7097 -8241
rect 7867 -8250 7875 -8234
rect 7890 -8250 7900 -8242
rect 7901 -8250 7909 -8234
rect 7148 -8290 7158 -8279
rect 7327 -8284 7371 -8250
rect 7399 -8284 7443 -8250
rect 7471 -8284 7515 -8250
rect 7615 -8284 7659 -8250
rect 7687 -8284 7803 -8250
rect 7831 -8284 7875 -8250
rect 7159 -8324 7203 -8290
rect 7148 -8374 7158 -8363
rect 7724 -8367 7768 -8333
rect 7159 -8408 7203 -8374
rect 7148 -8457 7158 -8446
rect 7159 -8491 7203 -8457
rect 7389 -8517 7433 -8483
rect 7434 -8517 7444 -8472
rect 7511 -8534 7519 -8416
rect 7534 -8483 7544 -8472
rect 7545 -8483 7553 -8450
rect 7581 -8483 7589 -8450
rect 7545 -8517 7589 -8483
rect 7590 -8517 7600 -8472
rect 7545 -8568 7553 -8517
rect 7581 -8568 7589 -8517
rect 7615 -8534 7623 -8417
rect 7712 -8458 7715 -8417
rect 7724 -8451 7768 -8417
rect 7724 -8534 7768 -8500
rect 7867 -8534 7875 -8284
rect 7901 -8284 7945 -8250
rect 8428 -8274 8472 -8240
rect 8524 -8274 8568 -8240
rect 8620 -8274 8664 -8240
rect 10127 -8241 10171 -8207
rect 10191 -8241 10246 -8207
rect 10271 -8241 10321 -8207
rect 7890 -8333 7900 -8322
rect 7901 -8333 7909 -8284
rect 8140 -8293 8150 -8285
rect 8240 -8293 8250 -8285
rect 8067 -8327 8183 -8293
rect 8251 -8327 8295 -8293
rect 8782 -8317 8826 -8283
rect 8878 -8317 8922 -8283
rect 8974 -8317 9018 -8283
rect 9070 -8317 9114 -8283
rect 9166 -8317 9210 -8283
rect 10191 -8324 10235 -8290
rect 10236 -8324 10246 -8279
rect 7901 -8367 7945 -8333
rect 8494 -8336 8504 -8328
rect 8594 -8336 8604 -8328
rect 7890 -8417 7900 -8406
rect 7901 -8417 7909 -8367
rect 8095 -8410 8139 -8376
rect 8140 -8410 8150 -8365
rect 8240 -8376 8250 -8365
rect 8421 -8370 8537 -8336
rect 8605 -8370 8649 -8336
rect 9330 -8360 9374 -8326
rect 9426 -8360 9470 -8326
rect 9522 -8360 9566 -8326
rect 9618 -8360 9662 -8326
rect 9714 -8360 9758 -8326
rect 9810 -8360 9854 -8326
rect 9906 -8360 9950 -8326
rect 8251 -8410 8295 -8376
rect 8884 -8379 8894 -8371
rect 8961 -8379 8969 -8363
rect 8984 -8379 8994 -8371
rect 8995 -8379 9003 -8363
rect 9049 -8371 9055 -8363
rect 7901 -8451 7945 -8417
rect 7890 -8500 7900 -8489
rect 7901 -8500 7909 -8451
rect 8095 -8494 8139 -8460
rect 8140 -8494 8150 -8449
rect 8240 -8460 8250 -8449
rect 8449 -8453 8493 -8419
rect 8494 -8453 8504 -8408
rect 8594 -8419 8604 -8408
rect 8775 -8413 8819 -8379
rect 8839 -8413 8894 -8379
rect 8919 -8413 8969 -8379
rect 8605 -8453 8649 -8419
rect 8251 -8494 8295 -8460
rect 7901 -8534 7945 -8500
rect 7901 -8568 7909 -8534
rect 6550 -8714 6559 -8706
rect 6550 -8722 6600 -8714
rect 6550 -8740 6559 -8722
rect 6847 -8723 6891 -8689
rect 6892 -8723 6902 -8681
rect 5489 -8853 5539 -8845
rect 5539 -8861 5550 -8853
rect 4297 -8906 4342 -8872
rect 4369 -8878 4414 -8872
rect 4441 -8878 4486 -8872
rect 4369 -8886 4486 -8878
rect 4560 -8882 4610 -8878
rect 4799 -8879 4810 -8868
rect 4899 -8879 4910 -8868
rect 4369 -8906 4414 -8886
rect 4441 -8906 4486 -8886
rect 4754 -8913 4810 -8879
rect 4910 -8913 4955 -8879
rect 5494 -8895 5550 -8861
rect 4722 -8921 4767 -8915
rect 4794 -8921 4839 -8915
rect 3388 -8959 3874 -8925
rect 4722 -8929 4839 -8921
rect 4910 -8929 4960 -8921
rect 5153 -8922 5164 -8911
rect 5253 -8922 5264 -8911
rect 5681 -8913 5697 -8845
rect 5722 -8879 5731 -8811
rect 5767 -8843 5776 -8775
rect 5801 -8809 5810 -8743
rect 5811 -8793 5856 -8759
rect 6014 -8838 6059 -8804
rect 5792 -8853 5842 -8845
rect 5781 -8861 5792 -8853
rect 5792 -8895 5837 -8861
rect 6014 -8906 6059 -8872
rect 4722 -8949 4767 -8929
rect 4794 -8949 4839 -8929
rect 5108 -8956 5164 -8922
rect 5264 -8956 5309 -8922
rect 3388 -8985 3861 -8959
rect 5076 -8964 5121 -8958
rect 5148 -8964 5193 -8958
rect 5539 -8961 5550 -8950
rect 3392 -8993 3603 -8985
rect 3408 -9003 3587 -8993
rect 3738 -9023 3783 -8985
rect 3991 -9002 4036 -8968
rect 4087 -9002 4132 -8968
rect 4183 -9002 4228 -8968
rect 4279 -9002 4324 -8968
rect 4375 -9002 4420 -8968
rect 4471 -9002 4516 -8968
rect 4567 -9002 4612 -8968
rect 5076 -8972 5193 -8964
rect 5264 -8972 5314 -8964
rect 5076 -8992 5121 -8972
rect 5148 -8992 5193 -8972
rect 5494 -8995 5550 -8961
rect 5681 -9001 5692 -8913
rect 6063 -8922 6072 -8788
rect 5781 -8961 5792 -8950
rect 6097 -8956 6106 -8762
rect 6137 -8778 6148 -8767
rect 6133 -8809 6148 -8778
rect 6459 -8796 6504 -8762
rect 5792 -8995 5837 -8961
rect 6037 -8991 6048 -8980
rect 2616 -9046 2636 -9038
rect 2640 -9050 2693 -9038
rect 2813 -9046 2846 -9038
rect 2746 -9050 2846 -9046
rect 2400 -9051 2434 -9050
rect 2239 -9067 2311 -9063
rect 2390 -9067 2450 -9063
rect 1979 -9088 2007 -9069
rect 1685 -9114 1727 -9088
rect 2062 -9101 2522 -9097
rect 2013 -9122 2041 -9103
rect 2062 -9111 2234 -9101
rect 2270 -9111 2370 -9101
rect 2381 -9111 2426 -9101
rect 2062 -9131 2427 -9111
rect 2477 -9131 2522 -9101
rect 2534 -9131 2553 -9097
rect 2568 -9164 2587 -9063
rect 2828 -9067 2846 -9050
rect 2947 -9078 2992 -9044
rect 3013 -9050 3289 -9038
rect 3346 -9050 3391 -9046
rect 3019 -9078 3064 -9050
rect 3067 -9077 3289 -9050
rect 3334 -9077 3445 -9050
rect 3593 -9062 3603 -9051
rect 3604 -9077 3649 -9062
rect 3028 -9132 3032 -9129
rect 3067 -9135 3661 -9077
rect 3672 -9123 3717 -9077
rect 3067 -9140 3319 -9135
rect 2610 -9150 2726 -9140
rect 2737 -9150 2928 -9140
rect 2929 -9150 2974 -9140
rect 2610 -9158 2975 -9150
rect 3025 -9158 3319 -9140
rect 2610 -9174 3319 -9158
rect 3067 -9200 3319 -9174
rect 3334 -9174 3445 -9135
rect 2726 -9248 2768 -9224
rect 2928 -9248 2975 -9224
rect 3067 -9458 3257 -9200
rect 3334 -9211 3391 -9174
rect 3392 -9211 3402 -9174
rect 3334 -9227 3393 -9211
rect 3509 -9227 3556 -9180
rect 3334 -9261 3556 -9227
rect 2687 -9970 3066 -9936
rect 3145 -9971 3191 -9458
rect 3200 -9971 3257 -9458
rect 3267 -9971 3269 -9308
rect 3279 -9971 3291 -9304
rect 3312 -9308 3313 -9304
rect 3334 -9308 3392 -9261
rect 3604 -9280 3649 -9135
rect 3570 -9308 3571 -9304
rect 3312 -9320 3319 -9308
rect 3308 -9971 3319 -9320
rect 3340 -9971 3391 -9308
rect 3570 -9309 3577 -9308
rect 3526 -9320 3577 -9309
rect 3537 -9971 3577 -9320
rect 3598 -9971 3649 -9280
rect 3659 -9971 3661 -9135
rect 3671 -9971 3717 -9123
rect 3726 -9971 3783 -9023
rect 4729 -9045 4774 -9011
rect 4825 -9045 4870 -9011
rect 4921 -9045 4966 -9011
rect 5430 -9035 5475 -9001
rect 5502 -9003 5547 -9001
rect 5489 -9011 5547 -9003
rect 5502 -9035 5547 -9011
rect 5574 -9035 5619 -9001
rect 5646 -9029 5692 -9001
rect 5792 -9011 5842 -9003
rect 5992 -9025 6048 -8991
rect 6133 -8992 6142 -8809
rect 6167 -8995 6176 -8812
rect 5646 -9035 5691 -9029
rect 5083 -9088 5128 -9054
rect 5179 -9088 5224 -9054
rect 5275 -9088 5320 -9054
rect 6179 -9076 6190 -8809
rect 6516 -8812 6520 -8742
rect 6550 -8819 6554 -8740
rect 7034 -8741 7049 -8673
rect 7075 -8707 7083 -8639
rect 7120 -8671 7128 -8603
rect 7154 -8637 7162 -8571
rect 7164 -8621 7208 -8587
rect 7365 -8666 7409 -8632
rect 7134 -8689 7144 -8681
rect 7145 -8723 7189 -8689
rect 7365 -8734 7409 -8700
rect 7034 -8753 7044 -8741
rect 7414 -8750 7422 -8616
rect 6809 -8819 7205 -8753
rect 7448 -8784 7456 -8590
rect 7488 -8606 7498 -8595
rect 7484 -8637 7498 -8606
rect 7810 -8624 7854 -8590
rect 6195 -8860 6240 -8826
rect 6544 -8830 6565 -8819
rect 6544 -8832 6554 -8830
rect 6195 -8928 6240 -8894
rect 6247 -8995 6256 -8860
rect 6478 -8874 6554 -8832
rect 6607 -8874 7205 -8819
rect 7343 -8853 7387 -8819
rect 7388 -8853 7398 -8808
rect 7484 -8820 7492 -8637
rect 7518 -8823 7526 -8640
rect 6478 -8877 7205 -8874
rect 6281 -8980 6290 -8892
rect 6393 -8900 6443 -8892
rect 6443 -8908 6454 -8900
rect 6398 -8942 6454 -8908
rect 6279 -8991 6290 -8980
rect 6281 -9025 6335 -8991
rect 6443 -9008 6454 -8997
rect 6398 -9042 6454 -9008
rect 6478 -9044 6633 -8877
rect 6809 -8899 7205 -8877
rect 6733 -8925 7205 -8899
rect 7530 -8904 7540 -8637
rect 7867 -8640 7870 -8570
rect 7546 -8688 7590 -8654
rect 7901 -8674 7904 -8568
rect 8095 -8577 8139 -8543
rect 8140 -8577 8150 -8532
rect 8240 -8543 8250 -8532
rect 8449 -8537 8493 -8503
rect 8494 -8537 8504 -8492
rect 8594 -8503 8604 -8492
rect 8839 -8496 8883 -8462
rect 8884 -8496 8894 -8451
rect 8605 -8537 8649 -8503
rect 8251 -8577 8295 -8543
rect 7546 -8756 7590 -8722
rect 7598 -8823 7606 -8688
rect 8160 -8691 8204 -8657
rect 8212 -8718 8220 -8641
rect 7632 -8808 7640 -8720
rect 7749 -8770 7793 -8736
rect 7794 -8770 7804 -8728
rect 7894 -8740 7904 -8729
rect 7905 -8774 7949 -8740
rect 8246 -8752 8254 -8607
rect 8449 -8620 8493 -8586
rect 8494 -8620 8504 -8575
rect 8594 -8586 8604 -8575
rect 8839 -8580 8883 -8546
rect 8884 -8580 8894 -8535
rect 8605 -8620 8649 -8586
rect 8514 -8734 8558 -8700
rect 8566 -8761 8574 -8684
rect 7630 -8819 7640 -8808
rect 8099 -8813 8143 -8779
rect 8144 -8813 8154 -8771
rect 8244 -8779 8254 -8771
rect 8255 -8813 8299 -8779
rect 8600 -8795 8608 -8650
rect 8839 -8663 8883 -8629
rect 8884 -8663 8894 -8618
rect 8961 -8679 8969 -8413
rect 8995 -8413 9039 -8379
rect 9040 -8413 9055 -8371
rect 8984 -8462 8994 -8451
rect 8995 -8462 9003 -8413
rect 9049 -8451 9055 -8413
rect 8995 -8496 9039 -8462
rect 9040 -8496 9055 -8451
rect 8984 -8546 8994 -8535
rect 8995 -8546 9003 -8496
rect 9049 -8535 9055 -8496
rect 8995 -8580 9039 -8546
rect 9040 -8580 9055 -8535
rect 8984 -8629 8994 -8618
rect 8995 -8629 9003 -8580
rect 9049 -8618 9055 -8580
rect 8984 -8697 8994 -8655
rect 8995 -8663 9039 -8629
rect 9040 -8663 9055 -8618
rect 8995 -8713 9003 -8663
rect 8904 -8777 8948 -8743
rect 8961 -8804 8964 -8727
rect 8995 -8809 8998 -8713
rect 7632 -8853 7640 -8819
rect 7641 -8853 7685 -8819
rect 7749 -8870 7793 -8836
rect 7794 -8870 7804 -8825
rect 7894 -8832 7904 -8821
rect 7905 -8866 7949 -8832
rect 8453 -8856 8497 -8822
rect 8498 -8856 8508 -8814
rect 8598 -8822 8608 -8814
rect 8609 -8856 8653 -8822
rect 9026 -8845 9036 -8697
rect 9049 -8713 9055 -8663
rect 9083 -8379 9089 -8363
rect 9140 -8379 9150 -8371
rect 9083 -8413 9133 -8379
rect 9151 -8413 9205 -8379
rect 9083 -8679 9089 -8413
rect 9861 -8422 9869 -8406
rect 9884 -8422 9894 -8414
rect 9895 -8422 9903 -8406
rect 10191 -8408 10235 -8374
rect 10236 -8408 10246 -8363
rect 9140 -8462 9150 -8451
rect 9321 -8456 9365 -8422
rect 9393 -8456 9437 -8422
rect 9465 -8456 9509 -8422
rect 9609 -8456 9653 -8422
rect 9681 -8456 9797 -8422
rect 9825 -8456 9869 -8422
rect 9151 -8496 9195 -8462
rect 9140 -8546 9150 -8535
rect 9718 -8539 9762 -8505
rect 9151 -8580 9195 -8546
rect 9140 -8629 9150 -8618
rect 9151 -8663 9195 -8629
rect 9383 -8689 9427 -8655
rect 9428 -8689 9438 -8644
rect 9505 -8706 9513 -8588
rect 9528 -8655 9538 -8644
rect 9539 -8655 9547 -8622
rect 9575 -8655 9583 -8622
rect 9539 -8689 9583 -8655
rect 9584 -8689 9594 -8644
rect 9539 -8740 9547 -8689
rect 9575 -8740 9583 -8689
rect 9609 -8706 9617 -8589
rect 9706 -8630 9709 -8589
rect 9718 -8623 9762 -8589
rect 9718 -8706 9762 -8672
rect 9861 -8706 9869 -8456
rect 9895 -8456 9939 -8422
rect 9884 -8505 9894 -8494
rect 9895 -8505 9903 -8456
rect 10191 -8491 10235 -8457
rect 10236 -8491 10246 -8446
rect 9895 -8539 9939 -8505
rect 9884 -8589 9894 -8578
rect 9895 -8589 9903 -8539
rect 10047 -8565 10153 -8499
rect 10313 -8507 10321 -8241
rect 10347 -8241 10391 -8207
rect 10392 -8241 10407 -8199
rect 10336 -8290 10346 -8279
rect 10347 -8290 10355 -8241
rect 10401 -8279 10407 -8241
rect 10347 -8324 10391 -8290
rect 10392 -8324 10407 -8279
rect 10336 -8374 10346 -8363
rect 10347 -8374 10355 -8324
rect 10401 -8363 10407 -8324
rect 10347 -8408 10391 -8374
rect 10392 -8408 10407 -8363
rect 10336 -8457 10346 -8446
rect 10347 -8457 10355 -8408
rect 10401 -8446 10407 -8408
rect 10336 -8525 10346 -8483
rect 10347 -8491 10391 -8457
rect 10392 -8491 10407 -8446
rect 10347 -8541 10355 -8491
rect 9895 -8623 9939 -8589
rect 10256 -8605 10300 -8571
rect 9884 -8672 9894 -8661
rect 9895 -8672 9903 -8623
rect 10313 -8632 10316 -8555
rect 10347 -8637 10350 -8541
rect 9895 -8706 9939 -8672
rect 10378 -8673 10388 -8525
rect 10401 -8541 10407 -8491
rect 10435 -8207 10441 -8191
rect 10492 -8207 10502 -8199
rect 10435 -8241 10485 -8207
rect 10503 -8241 10557 -8207
rect 11418 -8231 11462 -8197
rect 11514 -8231 11558 -8197
rect 11610 -8231 11654 -8197
rect 13581 -8207 13590 -8199
rect 13658 -8207 13665 -8191
rect 13681 -8207 13690 -8199
rect 13692 -8207 13699 -8191
rect 13746 -8199 13751 -8191
rect 10435 -8507 10441 -8241
rect 11211 -8250 11219 -8234
rect 11234 -8250 11244 -8242
rect 11245 -8250 11253 -8234
rect 10492 -8290 10502 -8279
rect 10671 -8284 10715 -8250
rect 10743 -8284 10787 -8250
rect 10815 -8284 10859 -8250
rect 10959 -8284 11003 -8250
rect 11031 -8284 11147 -8250
rect 11175 -8284 11219 -8250
rect 10503 -8324 10547 -8290
rect 10492 -8374 10502 -8363
rect 11068 -8367 11112 -8333
rect 10503 -8408 10547 -8374
rect 10492 -8457 10502 -8446
rect 10503 -8491 10547 -8457
rect 10733 -8517 10777 -8483
rect 10778 -8517 10788 -8472
rect 10855 -8534 10863 -8416
rect 10878 -8483 10888 -8472
rect 10889 -8483 10897 -8450
rect 10925 -8483 10933 -8450
rect 10889 -8517 10933 -8483
rect 10934 -8517 10944 -8472
rect 10889 -8568 10897 -8517
rect 10925 -8568 10933 -8517
rect 10959 -8534 10967 -8417
rect 11056 -8458 11059 -8417
rect 11068 -8451 11112 -8417
rect 11068 -8534 11112 -8500
rect 11211 -8534 11219 -8284
rect 11245 -8284 11289 -8250
rect 11772 -8274 11816 -8240
rect 11868 -8274 11912 -8240
rect 11964 -8274 12008 -8240
rect 13472 -8241 13515 -8207
rect 13536 -8241 13590 -8207
rect 13616 -8241 13665 -8207
rect 11234 -8333 11244 -8322
rect 11245 -8333 11253 -8284
rect 11484 -8293 11494 -8285
rect 11584 -8293 11594 -8285
rect 11411 -8327 11527 -8293
rect 11595 -8327 11639 -8293
rect 12126 -8317 12170 -8283
rect 12222 -8317 12266 -8283
rect 12318 -8317 12362 -8283
rect 12414 -8317 12458 -8283
rect 12510 -8317 12554 -8283
rect 13536 -8324 13579 -8290
rect 13581 -8324 13590 -8279
rect 11245 -8367 11289 -8333
rect 11838 -8336 11848 -8328
rect 11938 -8336 11948 -8328
rect 11234 -8417 11244 -8406
rect 11245 -8417 11253 -8367
rect 11439 -8410 11483 -8376
rect 11484 -8410 11494 -8365
rect 11584 -8376 11594 -8365
rect 11765 -8370 11881 -8336
rect 11949 -8370 11993 -8336
rect 12674 -8360 12718 -8326
rect 12770 -8360 12814 -8326
rect 12866 -8360 12910 -8326
rect 12962 -8360 13006 -8326
rect 13058 -8360 13102 -8326
rect 13154 -8360 13198 -8326
rect 13250 -8360 13294 -8326
rect 11595 -8410 11639 -8376
rect 12228 -8379 12238 -8371
rect 12305 -8379 12313 -8363
rect 12328 -8379 12338 -8371
rect 12339 -8379 12347 -8363
rect 12393 -8371 12399 -8363
rect 11245 -8451 11289 -8417
rect 11234 -8500 11244 -8489
rect 11245 -8500 11253 -8451
rect 11439 -8494 11483 -8460
rect 11484 -8494 11494 -8449
rect 11584 -8460 11594 -8449
rect 11793 -8453 11837 -8419
rect 11838 -8453 11848 -8408
rect 11938 -8419 11948 -8408
rect 12119 -8413 12163 -8379
rect 12183 -8413 12238 -8379
rect 12263 -8413 12313 -8379
rect 11949 -8453 11993 -8419
rect 11595 -8494 11639 -8460
rect 11245 -8534 11289 -8500
rect 11245 -8568 11253 -8534
rect 9895 -8740 9903 -8706
rect 10191 -8723 10235 -8689
rect 10236 -8723 10246 -8681
rect 7642 -8906 7686 -8872
rect 7714 -8906 7758 -8872
rect 7786 -8906 7830 -8872
rect 8099 -8913 8143 -8879
rect 8144 -8913 8154 -8868
rect 8244 -8879 8254 -8868
rect 8255 -8913 8299 -8879
rect 8839 -8895 8883 -8861
rect 8884 -8895 8894 -8853
rect 6733 -8959 7218 -8925
rect 8067 -8949 8111 -8915
rect 8139 -8949 8183 -8915
rect 8453 -8956 8497 -8922
rect 8498 -8956 8508 -8911
rect 8598 -8922 8608 -8911
rect 9026 -8913 9041 -8845
rect 9067 -8879 9075 -8811
rect 9112 -8843 9120 -8775
rect 9146 -8809 9154 -8743
rect 9156 -8793 9200 -8759
rect 9359 -8838 9403 -8804
rect 9126 -8861 9136 -8853
rect 9137 -8895 9181 -8861
rect 9359 -8906 9403 -8872
rect 8609 -8956 8653 -8922
rect 6733 -8985 7205 -8959
rect 6736 -8993 6947 -8985
rect 6752 -9003 6931 -8993
rect 6291 -9078 6336 -9044
rect 6363 -9050 6408 -9044
rect 6435 -9050 6633 -9044
rect 6363 -9058 6633 -9050
rect 6363 -9078 6408 -9058
rect 6435 -9078 6633 -9058
rect 5437 -9131 5482 -9097
rect 5533 -9131 5578 -9097
rect 5629 -9131 5674 -9097
rect 5725 -9131 5770 -9097
rect 5821 -9131 5866 -9097
rect 6478 -9114 6633 -9078
rect 6478 -9140 6663 -9114
rect 5985 -9174 6030 -9140
rect 6081 -9174 6126 -9140
rect 6177 -9174 6222 -9140
rect 6273 -9174 6318 -9140
rect 6369 -9174 6414 -9140
rect 6465 -9174 6663 -9140
rect 6478 -9200 6663 -9174
rect 6678 -9174 6789 -9050
rect 6937 -9062 6947 -9051
rect 6556 -9870 6601 -9200
rect 6678 -9228 6735 -9174
rect 6031 -9970 6410 -9936
rect 6490 -9971 6518 -9924
rect 6544 -9971 6601 -9870
rect 6690 -9971 6735 -9228
rect 6736 -9971 6746 -9174
rect 6948 -9971 6993 -9062
rect 7082 -9971 7127 -8985
rect 7336 -9002 7380 -8968
rect 7432 -9002 7476 -8968
rect 7528 -9002 7572 -8968
rect 7624 -9002 7668 -8968
rect 7720 -9002 7764 -8968
rect 7816 -9002 7860 -8968
rect 7912 -9002 7956 -8968
rect 8421 -8992 8465 -8958
rect 8493 -8992 8537 -8958
rect 8839 -8995 8883 -8961
rect 8884 -8995 8894 -8950
rect 9026 -9001 9036 -8913
rect 9408 -8922 9416 -8788
rect 9126 -8961 9136 -8950
rect 9442 -8956 9450 -8762
rect 9482 -8778 9492 -8767
rect 9478 -8809 9492 -8778
rect 9804 -8796 9848 -8762
rect 9137 -8995 9181 -8961
rect 8074 -9045 8118 -9011
rect 8170 -9045 8214 -9011
rect 8266 -9045 8310 -9011
rect 8775 -9035 8819 -9001
rect 8847 -9035 8891 -9001
rect 8919 -9035 8963 -9001
rect 8991 -9029 9036 -9001
rect 9337 -9025 9381 -8991
rect 9382 -9025 9392 -8980
rect 9478 -8992 9486 -8809
rect 9512 -8995 9520 -8812
rect 8991 -9035 9035 -9029
rect 8428 -9088 8472 -9054
rect 8524 -9088 8568 -9054
rect 8620 -9088 8664 -9054
rect 9524 -9076 9534 -8809
rect 9861 -8812 9864 -8742
rect 9895 -8819 9898 -8740
rect 10378 -8741 10393 -8673
rect 10419 -8707 10427 -8639
rect 10464 -8671 10472 -8603
rect 10498 -8637 10506 -8571
rect 10508 -8621 10552 -8587
rect 10709 -8666 10753 -8632
rect 10478 -8689 10488 -8681
rect 10489 -8723 10533 -8689
rect 10709 -8734 10753 -8700
rect 10378 -8753 10388 -8741
rect 10758 -8750 10766 -8616
rect 10153 -8819 10549 -8753
rect 10792 -8784 10800 -8590
rect 10832 -8606 10842 -8595
rect 10828 -8637 10842 -8606
rect 11154 -8624 11198 -8590
rect 9540 -8860 9584 -8826
rect 9889 -8830 9909 -8819
rect 9889 -8832 9898 -8830
rect 9540 -8928 9584 -8894
rect 9592 -8995 9600 -8860
rect 9823 -8874 9898 -8832
rect 9951 -8874 10549 -8819
rect 10687 -8853 10731 -8819
rect 10732 -8853 10742 -8808
rect 10828 -8820 10836 -8637
rect 10862 -8823 10870 -8640
rect 9823 -8877 10549 -8874
rect 9626 -8980 9634 -8892
rect 9743 -8942 9787 -8908
rect 9788 -8942 9798 -8900
rect 9624 -8991 9634 -8980
rect 9626 -9025 9634 -8991
rect 9635 -9025 9679 -8991
rect 9743 -9042 9787 -9008
rect 9788 -9042 9798 -8997
rect 9823 -9044 9977 -8877
rect 10153 -8899 10549 -8877
rect 10077 -8925 10549 -8899
rect 10874 -8904 10884 -8637
rect 11211 -8640 11214 -8570
rect 10890 -8688 10934 -8654
rect 11245 -8674 11248 -8568
rect 11439 -8577 11483 -8543
rect 11484 -8577 11494 -8532
rect 11584 -8543 11594 -8532
rect 11793 -8537 11837 -8503
rect 11838 -8537 11848 -8492
rect 11938 -8503 11948 -8492
rect 12183 -8496 12227 -8462
rect 12228 -8496 12238 -8451
rect 11949 -8537 11993 -8503
rect 11595 -8577 11639 -8543
rect 10890 -8756 10934 -8722
rect 10942 -8823 10950 -8688
rect 11504 -8691 11548 -8657
rect 11556 -8718 11564 -8641
rect 10976 -8808 10984 -8720
rect 11093 -8770 11137 -8736
rect 11138 -8770 11148 -8728
rect 11238 -8740 11248 -8729
rect 11249 -8774 11293 -8740
rect 11590 -8752 11598 -8607
rect 11793 -8620 11837 -8586
rect 11838 -8620 11848 -8575
rect 11938 -8586 11948 -8575
rect 12183 -8580 12227 -8546
rect 12228 -8580 12238 -8535
rect 11949 -8620 11993 -8586
rect 11858 -8734 11902 -8700
rect 11910 -8761 11918 -8684
rect 10974 -8819 10984 -8808
rect 11443 -8813 11487 -8779
rect 11488 -8813 11498 -8771
rect 11588 -8779 11598 -8771
rect 11599 -8813 11643 -8779
rect 11944 -8795 11952 -8650
rect 12183 -8663 12227 -8629
rect 12228 -8663 12238 -8618
rect 12305 -8679 12313 -8413
rect 12339 -8413 12383 -8379
rect 12384 -8413 12399 -8371
rect 12328 -8462 12338 -8451
rect 12339 -8462 12347 -8413
rect 12393 -8451 12399 -8413
rect 12339 -8496 12383 -8462
rect 12384 -8496 12399 -8451
rect 12328 -8546 12338 -8535
rect 12339 -8546 12347 -8496
rect 12393 -8535 12399 -8496
rect 12339 -8580 12383 -8546
rect 12384 -8580 12399 -8535
rect 12328 -8629 12338 -8618
rect 12339 -8629 12347 -8580
rect 12393 -8618 12399 -8580
rect 12328 -8697 12338 -8655
rect 12339 -8663 12383 -8629
rect 12384 -8663 12399 -8618
rect 12339 -8713 12347 -8663
rect 12248 -8777 12292 -8743
rect 12305 -8804 12308 -8727
rect 12339 -8809 12342 -8713
rect 10976 -8853 10984 -8819
rect 10985 -8853 11029 -8819
rect 11093 -8870 11137 -8836
rect 11138 -8870 11148 -8825
rect 11238 -8832 11248 -8821
rect 11249 -8866 11293 -8832
rect 11797 -8856 11841 -8822
rect 11842 -8856 11852 -8814
rect 11942 -8822 11952 -8814
rect 11953 -8856 11997 -8822
rect 12370 -8845 12380 -8697
rect 12393 -8713 12399 -8663
rect 12427 -8379 12433 -8363
rect 12484 -8379 12494 -8371
rect 12427 -8413 12477 -8379
rect 12495 -8413 12549 -8379
rect 12427 -8679 12433 -8413
rect 13205 -8422 13213 -8406
rect 13228 -8422 13238 -8414
rect 13239 -8422 13247 -8406
rect 13536 -8408 13579 -8374
rect 13581 -8408 13590 -8363
rect 12484 -8462 12494 -8451
rect 12665 -8456 12709 -8422
rect 12737 -8456 12781 -8422
rect 12809 -8456 12853 -8422
rect 12953 -8456 12997 -8422
rect 13025 -8456 13141 -8422
rect 13169 -8456 13213 -8422
rect 12495 -8496 12539 -8462
rect 12484 -8546 12494 -8535
rect 13062 -8539 13106 -8505
rect 12495 -8580 12539 -8546
rect 12484 -8629 12494 -8618
rect 12495 -8663 12539 -8629
rect 12727 -8689 12771 -8655
rect 12772 -8689 12782 -8644
rect 12849 -8706 12857 -8588
rect 12872 -8655 12882 -8644
rect 12883 -8655 12891 -8622
rect 12919 -8655 12927 -8622
rect 12883 -8689 12927 -8655
rect 12928 -8689 12938 -8644
rect 12883 -8740 12891 -8689
rect 12919 -8740 12927 -8689
rect 12953 -8706 12961 -8589
rect 13050 -8630 13053 -8589
rect 13062 -8623 13106 -8589
rect 13062 -8706 13106 -8672
rect 13205 -8706 13213 -8456
rect 13239 -8456 13283 -8422
rect 13228 -8505 13238 -8494
rect 13239 -8505 13247 -8456
rect 13536 -8491 13579 -8457
rect 13581 -8491 13590 -8446
rect 13239 -8539 13283 -8505
rect 13228 -8589 13238 -8578
rect 13239 -8589 13247 -8539
rect 13391 -8565 13498 -8499
rect 13658 -8507 13665 -8241
rect 13692 -8241 13735 -8207
rect 13737 -8241 13751 -8199
rect 13681 -8290 13690 -8279
rect 13692 -8290 13699 -8241
rect 13746 -8279 13751 -8241
rect 13692 -8324 13735 -8290
rect 13737 -8324 13751 -8279
rect 13681 -8374 13690 -8363
rect 13692 -8374 13699 -8324
rect 13746 -8363 13751 -8324
rect 13692 -8408 13735 -8374
rect 13737 -8408 13751 -8363
rect 13681 -8457 13690 -8446
rect 13692 -8457 13699 -8408
rect 13746 -8446 13751 -8408
rect 13692 -8491 13735 -8457
rect 13737 -8491 13751 -8446
rect 13681 -8525 13690 -8499
rect 13692 -8541 13699 -8491
rect 13239 -8623 13283 -8589
rect 13601 -8605 13644 -8571
rect 13228 -8672 13238 -8661
rect 13239 -8672 13247 -8623
rect 13658 -8632 13660 -8555
rect 13692 -8637 13694 -8541
rect 13239 -8706 13283 -8672
rect 13723 -8673 13732 -8525
rect 13746 -8541 13751 -8491
rect 13780 -8507 13785 -8191
rect 13837 -8207 13846 -8199
rect 13786 -8241 13829 -8207
rect 13848 -8241 13901 -8207
rect 14763 -8231 14806 -8197
rect 14859 -8231 14902 -8197
rect 14955 -8231 14998 -8197
rect 16925 -8207 16934 -8199
rect 17002 -8207 17009 -8191
rect 17025 -8207 17034 -8199
rect 17036 -8207 17043 -8191
rect 17090 -8199 17095 -8191
rect 14556 -8250 14563 -8234
rect 14579 -8250 14588 -8242
rect 14590 -8250 14597 -8234
rect 13837 -8290 13846 -8279
rect 14016 -8284 14059 -8250
rect 14088 -8284 14131 -8250
rect 14160 -8284 14203 -8250
rect 14304 -8284 14347 -8250
rect 14376 -8284 14491 -8250
rect 14520 -8284 14563 -8250
rect 13848 -8324 13891 -8290
rect 13837 -8374 13846 -8363
rect 14413 -8367 14456 -8333
rect 13848 -8408 13891 -8374
rect 13837 -8457 13846 -8446
rect 13848 -8491 13891 -8457
rect 14078 -8517 14121 -8483
rect 14123 -8517 14132 -8472
rect 14200 -8534 14207 -8416
rect 14223 -8483 14232 -8472
rect 14234 -8483 14241 -8450
rect 14270 -8483 14277 -8450
rect 14234 -8517 14277 -8483
rect 14279 -8517 14288 -8472
rect 14234 -8568 14241 -8517
rect 14270 -8568 14277 -8517
rect 14304 -8534 14311 -8417
rect 14401 -8458 14403 -8417
rect 14413 -8451 14456 -8417
rect 14413 -8534 14456 -8500
rect 14556 -8534 14563 -8284
rect 14590 -8284 14633 -8250
rect 15117 -8274 15160 -8240
rect 15213 -8274 15256 -8240
rect 15309 -8274 15352 -8240
rect 16816 -8241 16859 -8207
rect 16880 -8241 16934 -8207
rect 16960 -8241 17009 -8207
rect 14579 -8333 14588 -8322
rect 14590 -8333 14597 -8284
rect 14829 -8293 14838 -8285
rect 14929 -8293 14938 -8285
rect 14756 -8327 14827 -8293
rect 14828 -8327 14871 -8293
rect 14940 -8327 14983 -8293
rect 15471 -8317 15514 -8283
rect 15567 -8317 15610 -8283
rect 15663 -8317 15706 -8283
rect 15759 -8317 15802 -8283
rect 15855 -8317 15898 -8283
rect 16880 -8324 16923 -8290
rect 16925 -8324 16934 -8279
rect 14590 -8367 14633 -8333
rect 15183 -8336 15192 -8328
rect 15283 -8336 15292 -8328
rect 14579 -8417 14588 -8406
rect 14590 -8417 14597 -8367
rect 14784 -8410 14827 -8376
rect 14829 -8410 14838 -8365
rect 14929 -8376 14938 -8365
rect 15110 -8370 15181 -8336
rect 15182 -8370 15225 -8336
rect 15294 -8370 15337 -8336
rect 16019 -8360 16062 -8326
rect 16115 -8360 16158 -8326
rect 16211 -8360 16254 -8326
rect 16307 -8360 16350 -8326
rect 16403 -8360 16446 -8326
rect 16499 -8360 16542 -8326
rect 16595 -8360 16638 -8326
rect 14940 -8410 14983 -8376
rect 15573 -8379 15582 -8371
rect 15650 -8379 15657 -8363
rect 15673 -8379 15682 -8371
rect 15684 -8379 15691 -8363
rect 15738 -8371 15743 -8363
rect 14590 -8451 14633 -8417
rect 14579 -8500 14588 -8489
rect 14590 -8500 14597 -8451
rect 14784 -8494 14827 -8460
rect 14829 -8494 14838 -8449
rect 14929 -8460 14938 -8449
rect 15138 -8453 15181 -8419
rect 15183 -8453 15192 -8408
rect 15283 -8419 15292 -8408
rect 15464 -8413 15507 -8379
rect 15528 -8413 15582 -8379
rect 15608 -8413 15657 -8379
rect 15294 -8453 15337 -8419
rect 14940 -8494 14983 -8460
rect 14590 -8534 14633 -8500
rect 14590 -8568 14597 -8534
rect 13239 -8740 13247 -8706
rect 13536 -8723 13579 -8689
rect 13581 -8723 13590 -8681
rect 10986 -8906 11030 -8872
rect 11058 -8906 11102 -8872
rect 11130 -8906 11174 -8872
rect 11443 -8913 11487 -8879
rect 11488 -8913 11498 -8868
rect 11588 -8879 11598 -8868
rect 11599 -8913 11643 -8879
rect 12183 -8895 12227 -8861
rect 12228 -8895 12238 -8853
rect 10077 -8959 10562 -8925
rect 11411 -8949 11455 -8915
rect 11483 -8949 11527 -8915
rect 11797 -8956 11841 -8922
rect 11842 -8956 11852 -8911
rect 11942 -8922 11952 -8911
rect 12370 -8913 12385 -8845
rect 12411 -8879 12419 -8811
rect 12456 -8843 12464 -8775
rect 12490 -8809 12498 -8743
rect 12500 -8793 12544 -8759
rect 12703 -8838 12747 -8804
rect 12470 -8861 12480 -8853
rect 12481 -8895 12525 -8861
rect 12703 -8906 12747 -8872
rect 11953 -8956 11997 -8922
rect 10077 -8985 10549 -8959
rect 10081 -8993 10291 -8985
rect 10097 -9003 10275 -8993
rect 9636 -9078 9680 -9044
rect 9708 -9078 9752 -9044
rect 9780 -9078 9977 -9044
rect 8782 -9131 8826 -9097
rect 8878 -9131 8922 -9097
rect 8974 -9131 9018 -9097
rect 9070 -9131 9114 -9097
rect 9166 -9131 9210 -9097
rect 9823 -9114 9977 -9078
rect 9823 -9140 10007 -9114
rect 9330 -9174 9374 -9140
rect 9426 -9174 9470 -9140
rect 9522 -9174 9566 -9140
rect 9618 -9174 9662 -9140
rect 9714 -9174 9758 -9140
rect 9810 -9174 10007 -9140
rect 9823 -9200 10007 -9174
rect 10023 -9174 10133 -9050
rect 10282 -9062 10291 -9051
rect 9901 -9870 9945 -9200
rect 10023 -9228 10079 -9174
rect 9376 -9970 9754 -9936
rect 9835 -9971 9862 -9924
rect 9889 -9971 9945 -9870
rect 10035 -9971 10079 -9228
rect 10081 -9971 10090 -9174
rect 10293 -9971 10337 -9062
rect 10427 -9971 10471 -8985
rect 10680 -9002 10724 -8968
rect 10776 -9002 10820 -8968
rect 10872 -9002 10916 -8968
rect 10968 -9002 11012 -8968
rect 11064 -9002 11108 -8968
rect 11160 -9002 11204 -8968
rect 11256 -9002 11300 -8968
rect 11765 -8992 11809 -8958
rect 11837 -8992 11881 -8958
rect 12183 -8995 12227 -8961
rect 12228 -8995 12238 -8950
rect 12370 -9001 12380 -8913
rect 12752 -8922 12760 -8788
rect 12470 -8961 12480 -8950
rect 12786 -8956 12794 -8762
rect 12826 -8778 12836 -8767
rect 12822 -8809 12836 -8778
rect 13148 -8796 13192 -8762
rect 12481 -8995 12525 -8961
rect 11418 -9045 11462 -9011
rect 11514 -9045 11558 -9011
rect 11610 -9045 11654 -9011
rect 12119 -9035 12163 -9001
rect 12191 -9035 12235 -9001
rect 12263 -9035 12307 -9001
rect 12335 -9029 12380 -9001
rect 12681 -9025 12725 -8991
rect 12726 -9025 12736 -8980
rect 12822 -8992 12830 -8809
rect 12856 -8995 12864 -8812
rect 12335 -9035 12379 -9029
rect 11772 -9088 11816 -9054
rect 11868 -9088 11912 -9054
rect 11964 -9088 12008 -9054
rect 12868 -9076 12878 -8809
rect 13205 -8812 13208 -8742
rect 13239 -8819 13242 -8740
rect 13723 -8741 13737 -8673
rect 13764 -8707 13771 -8639
rect 13809 -8671 13816 -8603
rect 13843 -8637 13850 -8571
rect 13853 -8621 13896 -8587
rect 14054 -8666 14097 -8632
rect 13823 -8689 13832 -8681
rect 13834 -8723 13877 -8689
rect 14054 -8734 14097 -8700
rect 13723 -8753 13732 -8741
rect 14103 -8750 14110 -8616
rect 13498 -8819 13893 -8753
rect 14137 -8784 14144 -8590
rect 14177 -8606 14186 -8595
rect 14173 -8637 14186 -8606
rect 14499 -8624 14542 -8590
rect 12884 -8860 12928 -8826
rect 13233 -8830 13253 -8819
rect 13233 -8832 13242 -8830
rect 12884 -8928 12928 -8894
rect 12936 -8995 12944 -8860
rect 13167 -8874 13242 -8832
rect 13296 -8874 13893 -8819
rect 14032 -8853 14075 -8819
rect 14077 -8853 14086 -8808
rect 14173 -8820 14180 -8637
rect 14207 -8823 14214 -8640
rect 13167 -8877 13893 -8874
rect 12970 -8980 12978 -8892
rect 13087 -8942 13131 -8908
rect 13132 -8942 13142 -8900
rect 12968 -8991 12978 -8980
rect 12970 -9025 12978 -8991
rect 12979 -9025 13023 -8991
rect 13087 -9042 13131 -9008
rect 13132 -9042 13142 -8997
rect 13167 -9044 13321 -8877
rect 13498 -8899 13893 -8877
rect 13422 -8925 13893 -8899
rect 14219 -8904 14228 -8637
rect 14556 -8640 14558 -8570
rect 14235 -8688 14278 -8654
rect 14590 -8674 14592 -8568
rect 14784 -8577 14827 -8543
rect 14829 -8577 14838 -8532
rect 14929 -8543 14938 -8532
rect 15138 -8537 15181 -8503
rect 15183 -8537 15192 -8492
rect 15283 -8503 15292 -8492
rect 15528 -8496 15571 -8462
rect 15573 -8496 15582 -8451
rect 15294 -8537 15337 -8503
rect 14940 -8577 14983 -8543
rect 14235 -8756 14278 -8722
rect 14287 -8823 14294 -8688
rect 14849 -8691 14892 -8657
rect 14901 -8718 14908 -8641
rect 14321 -8808 14328 -8720
rect 14438 -8770 14481 -8736
rect 14483 -8770 14492 -8728
rect 14583 -8740 14592 -8729
rect 14594 -8774 14637 -8740
rect 14935 -8752 14942 -8607
rect 15138 -8620 15181 -8586
rect 15183 -8620 15192 -8575
rect 15283 -8586 15292 -8575
rect 15528 -8580 15571 -8546
rect 15573 -8580 15582 -8535
rect 15294 -8620 15337 -8586
rect 15203 -8734 15246 -8700
rect 15255 -8761 15262 -8684
rect 14319 -8819 14328 -8808
rect 14788 -8813 14831 -8779
rect 14833 -8813 14842 -8771
rect 14933 -8779 14942 -8771
rect 14944 -8813 14987 -8779
rect 15289 -8795 15296 -8650
rect 15528 -8663 15571 -8629
rect 15573 -8663 15582 -8618
rect 15650 -8679 15657 -8413
rect 15684 -8413 15727 -8379
rect 15729 -8413 15743 -8371
rect 15673 -8462 15682 -8451
rect 15684 -8462 15691 -8413
rect 15738 -8451 15743 -8413
rect 15684 -8496 15727 -8462
rect 15729 -8496 15743 -8451
rect 15673 -8546 15682 -8535
rect 15684 -8546 15691 -8496
rect 15738 -8535 15743 -8496
rect 15684 -8580 15727 -8546
rect 15729 -8580 15743 -8535
rect 15673 -8629 15682 -8618
rect 15684 -8629 15691 -8580
rect 15738 -8618 15743 -8580
rect 15684 -8663 15727 -8629
rect 15729 -8663 15743 -8618
rect 15673 -8697 15682 -8671
rect 15684 -8713 15691 -8663
rect 15593 -8777 15636 -8743
rect 15650 -8804 15652 -8727
rect 15684 -8809 15686 -8713
rect 14321 -8853 14328 -8819
rect 14330 -8853 14373 -8819
rect 14438 -8870 14481 -8836
rect 14483 -8870 14492 -8825
rect 14583 -8832 14592 -8821
rect 14594 -8866 14637 -8832
rect 15142 -8856 15185 -8822
rect 15187 -8856 15196 -8814
rect 15287 -8822 15296 -8814
rect 15298 -8856 15341 -8822
rect 15715 -8845 15724 -8697
rect 15738 -8713 15743 -8663
rect 15772 -8679 15777 -8363
rect 15829 -8379 15838 -8371
rect 15778 -8413 15821 -8379
rect 15840 -8413 15893 -8379
rect 16550 -8422 16557 -8406
rect 16573 -8422 16582 -8414
rect 16584 -8422 16591 -8406
rect 16880 -8408 16923 -8374
rect 16925 -8408 16934 -8363
rect 15829 -8462 15838 -8451
rect 16010 -8456 16053 -8422
rect 16082 -8456 16125 -8422
rect 16154 -8456 16197 -8422
rect 16298 -8456 16341 -8422
rect 16370 -8456 16485 -8422
rect 16514 -8456 16557 -8422
rect 15840 -8496 15883 -8462
rect 15829 -8546 15838 -8535
rect 16407 -8539 16450 -8505
rect 15840 -8580 15883 -8546
rect 15829 -8629 15838 -8618
rect 15840 -8663 15883 -8629
rect 16072 -8689 16115 -8655
rect 16117 -8689 16126 -8644
rect 16194 -8706 16201 -8588
rect 16217 -8655 16226 -8644
rect 16228 -8655 16235 -8622
rect 16264 -8655 16271 -8622
rect 16228 -8689 16271 -8655
rect 16273 -8689 16282 -8644
rect 16228 -8740 16235 -8689
rect 16264 -8740 16271 -8689
rect 16298 -8706 16305 -8589
rect 16395 -8630 16397 -8589
rect 16407 -8623 16450 -8589
rect 16407 -8706 16450 -8672
rect 16550 -8706 16557 -8456
rect 16584 -8456 16627 -8422
rect 16573 -8505 16582 -8494
rect 16584 -8505 16591 -8456
rect 16880 -8491 16923 -8457
rect 16925 -8491 16934 -8446
rect 16584 -8539 16627 -8505
rect 16573 -8589 16582 -8578
rect 16584 -8589 16591 -8539
rect 16735 -8565 16842 -8499
rect 17002 -8507 17009 -8241
rect 17036 -8241 17079 -8207
rect 17081 -8241 17095 -8199
rect 17025 -8290 17034 -8279
rect 17036 -8290 17043 -8241
rect 17090 -8279 17095 -8241
rect 17036 -8324 17079 -8290
rect 17081 -8324 17095 -8279
rect 17025 -8374 17034 -8363
rect 17036 -8374 17043 -8324
rect 17090 -8363 17095 -8324
rect 17036 -8408 17079 -8374
rect 17081 -8408 17095 -8363
rect 17025 -8457 17034 -8446
rect 17036 -8457 17043 -8408
rect 17090 -8446 17095 -8408
rect 17036 -8491 17079 -8457
rect 17081 -8491 17095 -8446
rect 17025 -8525 17034 -8499
rect 17036 -8541 17043 -8491
rect 16584 -8623 16627 -8589
rect 16945 -8605 16988 -8571
rect 16573 -8672 16582 -8661
rect 16584 -8672 16591 -8623
rect 17002 -8632 17004 -8555
rect 17036 -8637 17038 -8541
rect 16584 -8706 16627 -8672
rect 17067 -8673 17076 -8525
rect 17090 -8541 17095 -8491
rect 17124 -8507 17129 -8191
rect 17181 -8207 17190 -8199
rect 17130 -8241 17173 -8207
rect 17192 -8241 17245 -8207
rect 18107 -8231 18150 -8197
rect 18203 -8231 18246 -8197
rect 18299 -8231 18342 -8197
rect 20269 -8207 20278 -8199
rect 20346 -8207 20353 -8191
rect 20369 -8207 20378 -8199
rect 20380 -8207 20387 -8191
rect 20434 -8199 20439 -8191
rect 17900 -8250 17907 -8234
rect 17923 -8250 17932 -8242
rect 17934 -8250 17941 -8234
rect 17181 -8290 17190 -8279
rect 17360 -8284 17403 -8250
rect 17432 -8284 17475 -8250
rect 17504 -8284 17547 -8250
rect 17648 -8284 17691 -8250
rect 17720 -8284 17835 -8250
rect 17864 -8284 17907 -8250
rect 17192 -8324 17235 -8290
rect 17181 -8374 17190 -8363
rect 17757 -8367 17800 -8333
rect 17192 -8408 17235 -8374
rect 17181 -8457 17190 -8446
rect 17192 -8491 17235 -8457
rect 17422 -8517 17465 -8483
rect 17467 -8517 17476 -8472
rect 17544 -8534 17551 -8416
rect 17567 -8483 17576 -8472
rect 17578 -8483 17585 -8450
rect 17614 -8483 17621 -8450
rect 17578 -8517 17621 -8483
rect 17623 -8517 17632 -8472
rect 17578 -8568 17585 -8517
rect 17614 -8568 17621 -8517
rect 17648 -8534 17655 -8417
rect 17745 -8458 17747 -8417
rect 17757 -8451 17800 -8417
rect 17757 -8534 17800 -8500
rect 17900 -8534 17907 -8284
rect 17934 -8284 17977 -8250
rect 18461 -8274 18504 -8240
rect 18557 -8274 18600 -8240
rect 18653 -8274 18696 -8240
rect 20160 -8241 20203 -8207
rect 20224 -8241 20278 -8207
rect 20304 -8241 20353 -8207
rect 17923 -8333 17932 -8322
rect 17934 -8333 17941 -8284
rect 18173 -8293 18182 -8285
rect 18273 -8293 18282 -8285
rect 18100 -8327 18171 -8293
rect 18172 -8327 18215 -8293
rect 18284 -8327 18327 -8293
rect 18815 -8317 18858 -8283
rect 18911 -8317 18954 -8283
rect 19007 -8317 19050 -8283
rect 19103 -8317 19146 -8283
rect 19199 -8317 19242 -8283
rect 20224 -8324 20267 -8290
rect 20269 -8324 20278 -8279
rect 17934 -8367 17977 -8333
rect 18527 -8336 18536 -8328
rect 18627 -8336 18636 -8328
rect 17923 -8417 17932 -8406
rect 17934 -8417 17941 -8367
rect 18128 -8410 18171 -8376
rect 18173 -8410 18182 -8365
rect 18273 -8376 18282 -8365
rect 18454 -8370 18525 -8336
rect 18526 -8370 18569 -8336
rect 18638 -8370 18681 -8336
rect 19363 -8360 19406 -8326
rect 19459 -8360 19502 -8326
rect 19555 -8360 19598 -8326
rect 19651 -8360 19694 -8326
rect 19747 -8360 19790 -8326
rect 19843 -8360 19886 -8326
rect 19939 -8360 19982 -8326
rect 18284 -8410 18327 -8376
rect 18917 -8379 18926 -8371
rect 18994 -8379 19001 -8363
rect 19017 -8379 19026 -8371
rect 19028 -8379 19035 -8363
rect 19082 -8371 19087 -8363
rect 17934 -8451 17977 -8417
rect 17923 -8500 17932 -8489
rect 17934 -8500 17941 -8451
rect 18128 -8494 18171 -8460
rect 18173 -8494 18182 -8449
rect 18273 -8460 18282 -8449
rect 18482 -8453 18525 -8419
rect 18527 -8453 18536 -8408
rect 18627 -8419 18636 -8408
rect 18808 -8413 18851 -8379
rect 18872 -8413 18926 -8379
rect 18952 -8413 19001 -8379
rect 18638 -8453 18681 -8419
rect 18284 -8494 18327 -8460
rect 17934 -8534 17977 -8500
rect 17934 -8568 17941 -8534
rect 16584 -8740 16591 -8706
rect 16880 -8723 16923 -8689
rect 16925 -8723 16934 -8681
rect 14331 -8906 14374 -8872
rect 14403 -8906 14446 -8872
rect 14475 -8906 14518 -8872
rect 14788 -8913 14831 -8879
rect 14833 -8913 14842 -8868
rect 14933 -8879 14942 -8868
rect 14944 -8913 14987 -8879
rect 15528 -8895 15571 -8861
rect 15573 -8895 15582 -8853
rect 13422 -8959 13906 -8925
rect 14756 -8949 14799 -8915
rect 14828 -8949 14871 -8915
rect 15142 -8956 15185 -8922
rect 15187 -8956 15196 -8911
rect 15287 -8922 15296 -8911
rect 15715 -8913 15729 -8845
rect 15756 -8879 15763 -8811
rect 15801 -8843 15808 -8775
rect 15835 -8809 15842 -8743
rect 15845 -8793 15888 -8759
rect 16048 -8838 16091 -8804
rect 15815 -8861 15824 -8853
rect 15826 -8895 15869 -8861
rect 16048 -8906 16091 -8872
rect 15298 -8956 15341 -8922
rect 13422 -8985 13893 -8959
rect 13425 -8993 13635 -8985
rect 13441 -9003 13619 -8993
rect 12980 -9078 13024 -9044
rect 13052 -9078 13096 -9044
rect 13124 -9078 13321 -9044
rect 12126 -9131 12170 -9097
rect 12222 -9131 12266 -9097
rect 12318 -9131 12362 -9097
rect 12414 -9131 12458 -9097
rect 12510 -9131 12554 -9097
rect 13167 -9114 13321 -9078
rect 13167 -9140 13351 -9114
rect 12674 -9174 12718 -9140
rect 12770 -9174 12814 -9140
rect 12866 -9174 12910 -9140
rect 12962 -9174 13006 -9140
rect 13058 -9174 13102 -9140
rect 13154 -9174 13351 -9140
rect 13167 -9200 13351 -9174
rect 13367 -9174 13477 -9050
rect 13626 -9062 13635 -9051
rect 13245 -9870 13289 -9200
rect 13367 -9228 13423 -9174
rect 12720 -9970 13098 -9936
rect 13179 -9971 13206 -9924
rect 13233 -9971 13289 -9870
rect 13379 -9971 13423 -9228
rect 13425 -9971 13434 -9174
rect 13637 -9971 13681 -9062
rect 13771 -9971 13815 -8985
rect 14025 -9002 14068 -8968
rect 14121 -9002 14164 -8968
rect 14217 -9002 14260 -8968
rect 14313 -9002 14356 -8968
rect 14409 -9002 14452 -8968
rect 14505 -9002 14548 -8968
rect 14601 -9002 14644 -8968
rect 15110 -8992 15153 -8958
rect 15182 -8992 15225 -8958
rect 15528 -8995 15571 -8961
rect 15573 -8995 15582 -8950
rect 15715 -9001 15724 -8913
rect 16097 -8922 16104 -8788
rect 15815 -8961 15824 -8950
rect 16131 -8956 16138 -8762
rect 16171 -8778 16180 -8767
rect 16167 -8809 16180 -8778
rect 16493 -8796 16536 -8762
rect 15826 -8995 15869 -8961
rect 14763 -9045 14806 -9011
rect 14859 -9045 14902 -9011
rect 14955 -9045 14998 -9011
rect 15464 -9035 15507 -9001
rect 15536 -9035 15579 -9001
rect 15608 -9035 15651 -9001
rect 15680 -9029 15724 -9001
rect 16026 -9025 16069 -8991
rect 16071 -9025 16080 -8980
rect 16167 -8992 16174 -8809
rect 16201 -8995 16208 -8812
rect 15680 -9035 15723 -9029
rect 15117 -9088 15160 -9054
rect 15213 -9088 15256 -9054
rect 15309 -9088 15352 -9054
rect 16213 -9076 16222 -8809
rect 16550 -8812 16552 -8742
rect 16584 -8819 16586 -8740
rect 17067 -8741 17081 -8673
rect 17108 -8707 17115 -8639
rect 17153 -8671 17160 -8603
rect 17187 -8637 17194 -8571
rect 17197 -8621 17240 -8587
rect 17398 -8666 17441 -8632
rect 17167 -8689 17176 -8681
rect 17178 -8723 17221 -8689
rect 17398 -8734 17441 -8700
rect 17067 -8753 17076 -8741
rect 17447 -8750 17454 -8616
rect 16842 -8819 17237 -8753
rect 17481 -8784 17488 -8590
rect 17521 -8606 17530 -8595
rect 17517 -8637 17530 -8606
rect 17843 -8624 17886 -8590
rect 16229 -8860 16272 -8826
rect 16578 -8830 16597 -8819
rect 16578 -8832 16586 -8830
rect 16229 -8928 16272 -8894
rect 16281 -8995 16288 -8860
rect 16512 -8874 16586 -8832
rect 16640 -8874 17237 -8819
rect 17376 -8853 17419 -8819
rect 17421 -8853 17430 -8808
rect 17517 -8820 17524 -8637
rect 17551 -8823 17558 -8640
rect 16512 -8877 17237 -8874
rect 16315 -8980 16322 -8892
rect 16432 -8942 16475 -8908
rect 16477 -8942 16486 -8900
rect 16313 -8991 16322 -8980
rect 16315 -9025 16322 -8991
rect 16324 -9025 16367 -8991
rect 16432 -9042 16475 -9008
rect 16477 -9042 16486 -8997
rect 16512 -9044 16665 -8877
rect 16842 -8899 17237 -8877
rect 16766 -8925 17237 -8899
rect 17563 -8904 17572 -8637
rect 17900 -8640 17902 -8570
rect 17579 -8688 17622 -8654
rect 17934 -8674 17936 -8568
rect 18128 -8577 18171 -8543
rect 18173 -8577 18182 -8532
rect 18273 -8543 18282 -8532
rect 18482 -8537 18525 -8503
rect 18527 -8537 18536 -8492
rect 18627 -8503 18636 -8492
rect 18872 -8496 18915 -8462
rect 18917 -8496 18926 -8451
rect 18638 -8537 18681 -8503
rect 18284 -8577 18327 -8543
rect 17579 -8756 17622 -8722
rect 17631 -8823 17638 -8688
rect 18193 -8691 18236 -8657
rect 18245 -8718 18252 -8641
rect 17665 -8808 17672 -8720
rect 17782 -8770 17825 -8736
rect 17827 -8770 17836 -8728
rect 17927 -8740 17936 -8729
rect 17938 -8774 17981 -8740
rect 18279 -8752 18286 -8607
rect 18482 -8620 18525 -8586
rect 18527 -8620 18536 -8575
rect 18627 -8586 18636 -8575
rect 18872 -8580 18915 -8546
rect 18917 -8580 18926 -8535
rect 18638 -8620 18681 -8586
rect 18547 -8734 18590 -8700
rect 18599 -8761 18606 -8684
rect 17663 -8819 17672 -8808
rect 18132 -8813 18175 -8779
rect 18177 -8813 18186 -8771
rect 18277 -8779 18286 -8771
rect 18288 -8813 18331 -8779
rect 18633 -8795 18640 -8650
rect 18872 -8663 18915 -8629
rect 18917 -8663 18926 -8618
rect 18994 -8679 19001 -8413
rect 19028 -8413 19071 -8379
rect 19073 -8413 19087 -8371
rect 19017 -8462 19026 -8451
rect 19028 -8462 19035 -8413
rect 19082 -8451 19087 -8413
rect 19028 -8496 19071 -8462
rect 19073 -8496 19087 -8451
rect 19017 -8546 19026 -8535
rect 19028 -8546 19035 -8496
rect 19082 -8535 19087 -8496
rect 19028 -8580 19071 -8546
rect 19073 -8580 19087 -8535
rect 19017 -8629 19026 -8618
rect 19028 -8629 19035 -8580
rect 19082 -8618 19087 -8580
rect 19028 -8663 19071 -8629
rect 19073 -8663 19087 -8618
rect 19017 -8697 19026 -8671
rect 19028 -8713 19035 -8663
rect 18937 -8777 18980 -8743
rect 18994 -8804 18996 -8727
rect 19028 -8809 19030 -8713
rect 17665 -8853 17672 -8819
rect 17674 -8853 17717 -8819
rect 17782 -8870 17825 -8836
rect 17827 -8870 17836 -8825
rect 17927 -8832 17936 -8821
rect 17938 -8866 17981 -8832
rect 18486 -8856 18529 -8822
rect 18531 -8856 18540 -8814
rect 18631 -8822 18640 -8814
rect 18642 -8856 18685 -8822
rect 19059 -8845 19068 -8697
rect 19082 -8713 19087 -8663
rect 19116 -8679 19121 -8363
rect 19173 -8379 19182 -8371
rect 19122 -8413 19165 -8379
rect 19184 -8413 19237 -8379
rect 19894 -8422 19901 -8406
rect 19917 -8422 19926 -8414
rect 19928 -8422 19935 -8406
rect 20224 -8408 20267 -8374
rect 20269 -8408 20278 -8363
rect 19173 -8462 19182 -8451
rect 19354 -8456 19397 -8422
rect 19426 -8456 19469 -8422
rect 19498 -8456 19541 -8422
rect 19642 -8456 19685 -8422
rect 19714 -8456 19829 -8422
rect 19858 -8456 19901 -8422
rect 19184 -8496 19227 -8462
rect 19173 -8546 19182 -8535
rect 19751 -8539 19794 -8505
rect 19184 -8580 19227 -8546
rect 19173 -8629 19182 -8618
rect 19184 -8663 19227 -8629
rect 19416 -8689 19459 -8655
rect 19461 -8689 19470 -8644
rect 19538 -8706 19545 -8588
rect 19561 -8655 19570 -8644
rect 19572 -8655 19579 -8622
rect 19608 -8655 19615 -8622
rect 19572 -8689 19615 -8655
rect 19617 -8689 19626 -8644
rect 19572 -8740 19579 -8689
rect 19608 -8740 19615 -8689
rect 19642 -8706 19649 -8589
rect 19739 -8630 19741 -8589
rect 19751 -8623 19794 -8589
rect 19751 -8706 19794 -8672
rect 19894 -8706 19901 -8456
rect 19928 -8456 19971 -8422
rect 19917 -8505 19926 -8494
rect 19928 -8505 19935 -8456
rect 20224 -8491 20267 -8457
rect 20269 -8491 20278 -8446
rect 19928 -8539 19971 -8505
rect 19917 -8589 19926 -8578
rect 19928 -8589 19935 -8539
rect 20079 -8565 20186 -8499
rect 20346 -8507 20353 -8241
rect 20380 -8241 20423 -8207
rect 20425 -8241 20439 -8199
rect 20369 -8290 20378 -8279
rect 20380 -8290 20387 -8241
rect 20434 -8279 20439 -8241
rect 20380 -8324 20423 -8290
rect 20425 -8324 20439 -8279
rect 20369 -8374 20378 -8363
rect 20380 -8374 20387 -8324
rect 20434 -8363 20439 -8324
rect 20380 -8408 20423 -8374
rect 20425 -8408 20439 -8363
rect 20369 -8457 20378 -8446
rect 20380 -8457 20387 -8408
rect 20434 -8446 20439 -8408
rect 20380 -8491 20423 -8457
rect 20425 -8491 20439 -8446
rect 20369 -8525 20378 -8499
rect 20380 -8541 20387 -8491
rect 19928 -8623 19971 -8589
rect 20289 -8605 20332 -8571
rect 19917 -8672 19926 -8661
rect 19928 -8672 19935 -8623
rect 20346 -8632 20348 -8555
rect 20380 -8637 20382 -8541
rect 19928 -8706 19971 -8672
rect 20411 -8673 20420 -8525
rect 20434 -8541 20439 -8491
rect 20468 -8507 20473 -8191
rect 20525 -8207 20534 -8199
rect 20474 -8241 20517 -8207
rect 20536 -8241 20589 -8207
rect 21451 -8231 21494 -8197
rect 21547 -8231 21590 -8197
rect 21643 -8231 21686 -8197
rect 23613 -8207 23622 -8199
rect 23690 -8207 23697 -8191
rect 23713 -8207 23722 -8199
rect 23724 -8207 23731 -8191
rect 23778 -8199 23783 -8191
rect 21244 -8250 21251 -8234
rect 21267 -8250 21276 -8242
rect 21278 -8250 21285 -8234
rect 20525 -8290 20534 -8279
rect 20704 -8284 20747 -8250
rect 20776 -8284 20819 -8250
rect 20848 -8284 20891 -8250
rect 20992 -8284 21035 -8250
rect 21064 -8284 21179 -8250
rect 21208 -8284 21251 -8250
rect 20536 -8324 20579 -8290
rect 20525 -8374 20534 -8363
rect 21101 -8367 21144 -8333
rect 20536 -8408 20579 -8374
rect 20525 -8457 20534 -8446
rect 20536 -8491 20579 -8457
rect 20766 -8517 20809 -8483
rect 20811 -8517 20820 -8472
rect 20888 -8534 20895 -8416
rect 20911 -8483 20920 -8472
rect 20922 -8483 20929 -8450
rect 20958 -8483 20965 -8450
rect 20922 -8517 20965 -8483
rect 20967 -8517 20976 -8472
rect 20922 -8568 20929 -8517
rect 20958 -8568 20965 -8517
rect 20992 -8534 20999 -8417
rect 21089 -8458 21091 -8417
rect 21101 -8451 21144 -8417
rect 21101 -8534 21144 -8500
rect 21244 -8534 21251 -8284
rect 21278 -8284 21321 -8250
rect 21805 -8274 21848 -8240
rect 21901 -8274 21944 -8240
rect 21997 -8274 22040 -8240
rect 23504 -8241 23547 -8207
rect 23568 -8241 23622 -8207
rect 23648 -8241 23697 -8207
rect 21267 -8333 21276 -8322
rect 21278 -8333 21285 -8284
rect 21517 -8293 21526 -8285
rect 21617 -8293 21626 -8285
rect 21444 -8327 21515 -8293
rect 21516 -8327 21559 -8293
rect 21628 -8327 21671 -8293
rect 22159 -8317 22202 -8283
rect 22255 -8317 22298 -8283
rect 22351 -8317 22394 -8283
rect 22447 -8317 22490 -8283
rect 22543 -8317 22586 -8283
rect 23568 -8324 23611 -8290
rect 23613 -8324 23622 -8279
rect 21278 -8367 21321 -8333
rect 21871 -8336 21880 -8328
rect 21971 -8336 21980 -8328
rect 21267 -8417 21276 -8406
rect 21278 -8417 21285 -8367
rect 21472 -8410 21515 -8376
rect 21517 -8410 21526 -8365
rect 21617 -8376 21626 -8365
rect 21798 -8370 21869 -8336
rect 21870 -8370 21913 -8336
rect 21982 -8370 22025 -8336
rect 22707 -8360 22750 -8326
rect 22803 -8360 22846 -8326
rect 22899 -8360 22942 -8326
rect 22995 -8360 23038 -8326
rect 23091 -8360 23134 -8326
rect 23187 -8360 23230 -8326
rect 23283 -8360 23326 -8326
rect 21628 -8410 21671 -8376
rect 22261 -8379 22270 -8371
rect 22338 -8379 22345 -8363
rect 22361 -8379 22370 -8371
rect 22372 -8379 22379 -8363
rect 22426 -8371 22431 -8363
rect 21278 -8451 21321 -8417
rect 21267 -8500 21276 -8489
rect 21278 -8500 21285 -8451
rect 21472 -8494 21515 -8460
rect 21517 -8494 21526 -8449
rect 21617 -8460 21626 -8449
rect 21826 -8453 21869 -8419
rect 21871 -8453 21880 -8408
rect 21971 -8419 21980 -8408
rect 22152 -8413 22195 -8379
rect 22216 -8413 22270 -8379
rect 22296 -8413 22345 -8379
rect 21982 -8453 22025 -8419
rect 21628 -8494 21671 -8460
rect 21278 -8534 21321 -8500
rect 21278 -8568 21285 -8534
rect 19928 -8740 19935 -8706
rect 20224 -8723 20267 -8689
rect 20269 -8723 20278 -8681
rect 17675 -8906 17718 -8872
rect 17747 -8906 17790 -8872
rect 17819 -8906 17862 -8872
rect 18132 -8913 18175 -8879
rect 18177 -8913 18186 -8868
rect 18277 -8879 18286 -8868
rect 18288 -8913 18331 -8879
rect 18872 -8895 18915 -8861
rect 18917 -8895 18926 -8853
rect 16766 -8959 17250 -8925
rect 18100 -8949 18143 -8915
rect 18172 -8949 18215 -8915
rect 18486 -8956 18529 -8922
rect 18531 -8956 18540 -8911
rect 18631 -8922 18640 -8911
rect 19059 -8913 19073 -8845
rect 19100 -8879 19107 -8811
rect 19145 -8843 19152 -8775
rect 19179 -8809 19186 -8743
rect 19189 -8793 19232 -8759
rect 19392 -8838 19435 -8804
rect 19159 -8861 19168 -8853
rect 19170 -8895 19213 -8861
rect 19392 -8906 19435 -8872
rect 18642 -8956 18685 -8922
rect 16766 -8985 17237 -8959
rect 16770 -8993 16979 -8985
rect 16786 -9003 16963 -8993
rect 16325 -9078 16368 -9044
rect 16397 -9078 16440 -9044
rect 16469 -9078 16665 -9044
rect 15471 -9131 15514 -9097
rect 15567 -9131 15610 -9097
rect 15663 -9131 15706 -9097
rect 15759 -9131 15802 -9097
rect 15855 -9131 15898 -9097
rect 16512 -9114 16665 -9078
rect 16512 -9140 16695 -9114
rect 16019 -9174 16062 -9140
rect 16115 -9174 16158 -9140
rect 16211 -9174 16254 -9140
rect 16307 -9174 16350 -9140
rect 16403 -9174 16446 -9140
rect 16499 -9174 16695 -9140
rect 16512 -9200 16695 -9174
rect 16712 -9174 16821 -9050
rect 16971 -9062 16979 -9051
rect 16590 -9870 16633 -9200
rect 16712 -9228 16723 -9174
rect 16065 -9970 16442 -9936
rect 16524 -9971 16550 -9924
rect 16578 -9971 16633 -9870
rect 16724 -9971 16767 -9174
rect 16770 -9971 16778 -9174
rect 16982 -9971 17025 -9062
rect 17116 -9971 17159 -8985
rect 17369 -9002 17412 -8968
rect 17465 -9002 17508 -8968
rect 17561 -9002 17604 -8968
rect 17657 -9002 17700 -8968
rect 17753 -9002 17796 -8968
rect 17849 -9002 17892 -8968
rect 17945 -9002 17988 -8968
rect 18454 -8992 18497 -8958
rect 18526 -8992 18569 -8958
rect 18872 -8995 18915 -8961
rect 18917 -8995 18926 -8950
rect 19059 -9001 19068 -8913
rect 19441 -8922 19448 -8788
rect 19159 -8961 19168 -8950
rect 19475 -8956 19482 -8762
rect 19515 -8778 19524 -8767
rect 19511 -8809 19524 -8778
rect 19837 -8796 19880 -8762
rect 19170 -8995 19213 -8961
rect 18107 -9045 18150 -9011
rect 18203 -9045 18246 -9011
rect 18299 -9045 18342 -9011
rect 18808 -9035 18851 -9001
rect 18880 -9035 18923 -9001
rect 18952 -9035 18995 -9001
rect 19024 -9029 19068 -9001
rect 19370 -9025 19413 -8991
rect 19415 -9025 19424 -8980
rect 19511 -8992 19518 -8809
rect 19545 -8995 19552 -8812
rect 19024 -9035 19067 -9029
rect 18461 -9088 18504 -9054
rect 18557 -9088 18600 -9054
rect 18653 -9088 18696 -9054
rect 19557 -9076 19566 -8809
rect 19894 -8812 19896 -8742
rect 19928 -8819 19930 -8740
rect 20411 -8741 20425 -8673
rect 20452 -8707 20459 -8639
rect 20497 -8671 20504 -8603
rect 20531 -8637 20538 -8571
rect 20541 -8621 20584 -8587
rect 20742 -8666 20785 -8632
rect 20511 -8689 20520 -8681
rect 20522 -8723 20565 -8689
rect 20742 -8734 20785 -8700
rect 20411 -8753 20420 -8741
rect 20791 -8750 20798 -8616
rect 20186 -8819 20581 -8753
rect 20825 -8784 20832 -8590
rect 20865 -8606 20874 -8595
rect 20861 -8637 20874 -8606
rect 21187 -8624 21230 -8590
rect 19573 -8860 19616 -8826
rect 19922 -8830 19941 -8819
rect 19922 -8832 19930 -8830
rect 19573 -8928 19616 -8894
rect 19625 -8995 19632 -8860
rect 19856 -8874 19930 -8832
rect 19984 -8874 20581 -8819
rect 20720 -8853 20763 -8819
rect 20765 -8853 20774 -8808
rect 20861 -8820 20868 -8637
rect 20895 -8823 20902 -8640
rect 19856 -8877 20581 -8874
rect 19659 -8980 19666 -8892
rect 19776 -8942 19819 -8908
rect 19821 -8942 19830 -8900
rect 19657 -8991 19666 -8980
rect 19659 -9025 19666 -8991
rect 19668 -9025 19711 -8991
rect 19776 -9042 19819 -9008
rect 19821 -9042 19830 -8997
rect 19856 -9044 20009 -8877
rect 20186 -8899 20581 -8877
rect 20110 -8925 20581 -8899
rect 20907 -8904 20916 -8637
rect 21244 -8640 21246 -8570
rect 20923 -8688 20966 -8654
rect 21278 -8674 21280 -8568
rect 21472 -8577 21515 -8543
rect 21517 -8577 21526 -8532
rect 21617 -8543 21626 -8532
rect 21826 -8537 21869 -8503
rect 21871 -8537 21880 -8492
rect 21971 -8503 21980 -8492
rect 22216 -8496 22259 -8462
rect 22261 -8496 22270 -8451
rect 21982 -8537 22025 -8503
rect 21628 -8577 21671 -8543
rect 20923 -8756 20966 -8722
rect 20975 -8823 20982 -8688
rect 21537 -8691 21580 -8657
rect 21589 -8718 21596 -8641
rect 21009 -8808 21016 -8720
rect 21126 -8770 21169 -8736
rect 21171 -8770 21180 -8728
rect 21271 -8740 21280 -8729
rect 21282 -8774 21325 -8740
rect 21623 -8752 21630 -8607
rect 21826 -8620 21869 -8586
rect 21871 -8620 21880 -8575
rect 21971 -8586 21980 -8575
rect 22216 -8580 22259 -8546
rect 22261 -8580 22270 -8535
rect 21982 -8620 22025 -8586
rect 21891 -8734 21934 -8700
rect 21943 -8761 21950 -8684
rect 21007 -8819 21016 -8808
rect 21476 -8813 21519 -8779
rect 21521 -8813 21530 -8771
rect 21621 -8779 21630 -8771
rect 21632 -8813 21675 -8779
rect 21977 -8795 21984 -8650
rect 22216 -8663 22259 -8629
rect 22261 -8663 22270 -8618
rect 22338 -8679 22345 -8413
rect 22372 -8413 22415 -8379
rect 22417 -8413 22431 -8371
rect 22361 -8462 22370 -8451
rect 22372 -8462 22379 -8413
rect 22426 -8451 22431 -8413
rect 22372 -8496 22415 -8462
rect 22417 -8496 22431 -8451
rect 22361 -8546 22370 -8535
rect 22372 -8546 22379 -8496
rect 22426 -8535 22431 -8496
rect 22372 -8580 22415 -8546
rect 22417 -8580 22431 -8535
rect 22361 -8629 22370 -8618
rect 22372 -8629 22379 -8580
rect 22426 -8618 22431 -8580
rect 22372 -8663 22415 -8629
rect 22417 -8663 22431 -8618
rect 22361 -8697 22370 -8671
rect 22372 -8713 22379 -8663
rect 22281 -8777 22324 -8743
rect 22338 -8804 22340 -8727
rect 22372 -8809 22374 -8713
rect 21009 -8853 21016 -8819
rect 21018 -8853 21061 -8819
rect 21126 -8870 21169 -8836
rect 21171 -8870 21180 -8825
rect 21271 -8832 21280 -8821
rect 21282 -8866 21325 -8832
rect 21830 -8856 21873 -8822
rect 21875 -8856 21884 -8814
rect 21975 -8822 21984 -8814
rect 21986 -8856 22029 -8822
rect 22403 -8845 22412 -8697
rect 22426 -8713 22431 -8663
rect 22460 -8679 22465 -8363
rect 22517 -8379 22526 -8371
rect 22466 -8413 22509 -8379
rect 22528 -8413 22581 -8379
rect 23238 -8422 23245 -8406
rect 23261 -8422 23270 -8414
rect 23272 -8422 23279 -8406
rect 23568 -8408 23611 -8374
rect 23613 -8408 23622 -8363
rect 22517 -8462 22526 -8451
rect 22698 -8456 22741 -8422
rect 22770 -8456 22813 -8422
rect 22842 -8456 22885 -8422
rect 22986 -8456 23029 -8422
rect 23058 -8456 23173 -8422
rect 23202 -8456 23245 -8422
rect 22528 -8496 22571 -8462
rect 22517 -8546 22526 -8535
rect 23095 -8539 23138 -8505
rect 22528 -8580 22571 -8546
rect 22517 -8629 22526 -8618
rect 22528 -8663 22571 -8629
rect 22760 -8689 22803 -8655
rect 22805 -8689 22814 -8644
rect 22882 -8706 22889 -8588
rect 22905 -8655 22914 -8644
rect 22916 -8655 22923 -8622
rect 22952 -8655 22959 -8622
rect 22916 -8689 22959 -8655
rect 22961 -8689 22970 -8644
rect 22916 -8740 22923 -8689
rect 22952 -8740 22959 -8689
rect 22986 -8706 22993 -8589
rect 23083 -8630 23085 -8589
rect 23095 -8623 23138 -8589
rect 23095 -8706 23138 -8672
rect 23238 -8706 23245 -8456
rect 23272 -8456 23315 -8422
rect 23261 -8505 23270 -8494
rect 23272 -8505 23279 -8456
rect 23568 -8491 23611 -8457
rect 23613 -8491 23622 -8446
rect 23272 -8539 23315 -8505
rect 23261 -8589 23270 -8578
rect 23272 -8589 23279 -8539
rect 23423 -8565 23530 -8499
rect 23690 -8507 23697 -8241
rect 23724 -8241 23767 -8207
rect 23769 -8241 23783 -8199
rect 23713 -8290 23722 -8279
rect 23724 -8290 23731 -8241
rect 23778 -8279 23783 -8241
rect 23724 -8324 23767 -8290
rect 23769 -8324 23783 -8279
rect 23713 -8374 23722 -8363
rect 23724 -8374 23731 -8324
rect 23778 -8363 23783 -8324
rect 23724 -8408 23767 -8374
rect 23769 -8408 23783 -8363
rect 23713 -8457 23722 -8446
rect 23724 -8457 23731 -8408
rect 23778 -8446 23783 -8408
rect 23724 -8491 23767 -8457
rect 23769 -8491 23783 -8446
rect 23713 -8525 23722 -8499
rect 23724 -8541 23731 -8491
rect 23272 -8623 23315 -8589
rect 23633 -8605 23676 -8571
rect 23261 -8672 23270 -8661
rect 23272 -8672 23279 -8623
rect 23690 -8632 23692 -8555
rect 23724 -8637 23726 -8541
rect 23272 -8706 23315 -8672
rect 23755 -8673 23764 -8525
rect 23778 -8541 23783 -8491
rect 23812 -8507 23817 -8191
rect 23869 -8207 23878 -8199
rect 23818 -8241 23861 -8207
rect 23880 -8241 23933 -8207
rect 24795 -8231 24838 -8197
rect 24891 -8231 24934 -8197
rect 24987 -8231 25030 -8197
rect 26958 -8207 26966 -8199
rect 27035 -8207 27041 -8191
rect 27058 -8207 27066 -8199
rect 27069 -8207 27075 -8191
rect 24588 -8250 24595 -8234
rect 24611 -8250 24620 -8242
rect 24622 -8250 24629 -8234
rect 23869 -8290 23878 -8279
rect 24048 -8284 24091 -8250
rect 24120 -8284 24163 -8250
rect 24192 -8284 24235 -8250
rect 24336 -8284 24379 -8250
rect 24408 -8284 24523 -8250
rect 24552 -8284 24595 -8250
rect 23880 -8324 23923 -8290
rect 23869 -8374 23878 -8363
rect 24445 -8367 24488 -8333
rect 23880 -8408 23923 -8374
rect 23869 -8457 23878 -8446
rect 23880 -8491 23923 -8457
rect 24110 -8517 24153 -8483
rect 24155 -8517 24164 -8472
rect 24232 -8534 24239 -8416
rect 24255 -8483 24264 -8472
rect 24266 -8483 24273 -8450
rect 24302 -8483 24309 -8450
rect 24266 -8517 24309 -8483
rect 24311 -8517 24320 -8472
rect 24266 -8568 24273 -8517
rect 24302 -8568 24309 -8517
rect 24336 -8534 24343 -8417
rect 24433 -8458 24435 -8417
rect 24445 -8451 24488 -8417
rect 24445 -8534 24488 -8500
rect 24588 -8534 24595 -8284
rect 24622 -8284 24665 -8250
rect 25149 -8274 25192 -8240
rect 25245 -8274 25288 -8240
rect 25341 -8274 25384 -8240
rect 26849 -8241 26891 -8207
rect 26913 -8241 26966 -8207
rect 26993 -8241 27041 -8207
rect 24611 -8333 24620 -8322
rect 24622 -8333 24629 -8284
rect 24861 -8293 24870 -8285
rect 24961 -8293 24970 -8285
rect 24788 -8327 24859 -8293
rect 24860 -8327 24903 -8293
rect 24972 -8327 25015 -8293
rect 25503 -8317 25546 -8283
rect 25599 -8317 25642 -8283
rect 25695 -8317 25738 -8283
rect 25791 -8317 25834 -8283
rect 25887 -8317 25930 -8283
rect 26913 -8324 26955 -8290
rect 26958 -8324 26966 -8279
rect 24622 -8367 24665 -8333
rect 25215 -8336 25224 -8328
rect 25315 -8336 25324 -8328
rect 24611 -8417 24620 -8406
rect 24622 -8417 24629 -8367
rect 24816 -8410 24859 -8376
rect 24861 -8410 24870 -8365
rect 24961 -8376 24970 -8365
rect 25142 -8370 25213 -8336
rect 25214 -8370 25257 -8336
rect 25326 -8370 25369 -8336
rect 26051 -8360 26094 -8326
rect 26147 -8360 26190 -8326
rect 26243 -8360 26286 -8326
rect 26339 -8360 26382 -8326
rect 26435 -8360 26478 -8326
rect 26531 -8360 26574 -8326
rect 26627 -8360 26670 -8326
rect 24972 -8410 25015 -8376
rect 25605 -8379 25614 -8371
rect 25682 -8379 25689 -8363
rect 25705 -8379 25714 -8371
rect 25716 -8379 25723 -8363
rect 25770 -8371 25775 -8363
rect 24622 -8451 24665 -8417
rect 24611 -8500 24620 -8489
rect 24622 -8500 24629 -8451
rect 24816 -8494 24859 -8460
rect 24861 -8494 24870 -8449
rect 24961 -8460 24970 -8449
rect 25170 -8453 25213 -8419
rect 25215 -8453 25224 -8408
rect 25315 -8419 25324 -8408
rect 25496 -8413 25539 -8379
rect 25560 -8413 25614 -8379
rect 25640 -8413 25689 -8379
rect 25326 -8453 25369 -8419
rect 24972 -8494 25015 -8460
rect 24622 -8534 24665 -8500
rect 24622 -8568 24629 -8534
rect 23272 -8740 23279 -8706
rect 23568 -8723 23611 -8689
rect 23613 -8723 23622 -8681
rect 21019 -8906 21062 -8872
rect 21091 -8906 21134 -8872
rect 21163 -8906 21206 -8872
rect 21476 -8913 21519 -8879
rect 21521 -8913 21530 -8868
rect 21621 -8879 21630 -8868
rect 21632 -8913 21675 -8879
rect 22216 -8895 22259 -8861
rect 22261 -8895 22270 -8853
rect 20110 -8959 20594 -8925
rect 21444 -8949 21487 -8915
rect 21516 -8949 21559 -8915
rect 21830 -8956 21873 -8922
rect 21875 -8956 21884 -8911
rect 21975 -8922 21984 -8911
rect 22403 -8913 22417 -8845
rect 22444 -8879 22451 -8811
rect 22489 -8843 22496 -8775
rect 22523 -8809 22530 -8743
rect 22533 -8793 22576 -8759
rect 22736 -8838 22779 -8804
rect 22503 -8861 22512 -8853
rect 22514 -8895 22557 -8861
rect 22736 -8906 22779 -8872
rect 21986 -8956 22029 -8922
rect 20110 -8985 20581 -8959
rect 20114 -8993 20323 -8985
rect 20130 -9003 20307 -8993
rect 19669 -9078 19712 -9044
rect 19741 -9078 19784 -9044
rect 19813 -9078 20009 -9044
rect 18815 -9131 18858 -9097
rect 18911 -9131 18954 -9097
rect 19007 -9131 19050 -9097
rect 19103 -9131 19146 -9097
rect 19199 -9131 19242 -9097
rect 19856 -9114 20009 -9078
rect 19856 -9140 20039 -9114
rect 19363 -9174 19406 -9140
rect 19459 -9174 19502 -9140
rect 19555 -9174 19598 -9140
rect 19651 -9174 19694 -9140
rect 19747 -9174 19790 -9140
rect 19843 -9174 20039 -9140
rect 19856 -9200 20039 -9174
rect 20056 -9174 20165 -9050
rect 20315 -9062 20323 -9051
rect 19934 -9870 19977 -9200
rect 20056 -9228 20067 -9174
rect 19409 -9970 19786 -9936
rect 19868 -9971 19894 -9924
rect 19922 -9971 19977 -9870
rect 20068 -9971 20111 -9174
rect 20114 -9971 20122 -9174
rect 20326 -9971 20369 -9062
rect 20460 -9971 20503 -8985
rect 20713 -9002 20756 -8968
rect 20809 -9002 20852 -8968
rect 20905 -9002 20948 -8968
rect 21001 -9002 21044 -8968
rect 21097 -9002 21140 -8968
rect 21193 -9002 21236 -8968
rect 21289 -9002 21332 -8968
rect 21798 -8992 21841 -8958
rect 21870 -8992 21913 -8958
rect 22216 -8995 22259 -8961
rect 22261 -8995 22270 -8950
rect 22403 -9001 22412 -8913
rect 22785 -8922 22792 -8788
rect 22503 -8961 22512 -8950
rect 22819 -8956 22826 -8762
rect 22859 -8778 22868 -8767
rect 22855 -8809 22868 -8778
rect 23181 -8796 23224 -8762
rect 22514 -8995 22557 -8961
rect 21451 -9045 21494 -9011
rect 21547 -9045 21590 -9011
rect 21643 -9045 21686 -9011
rect 22152 -9035 22195 -9001
rect 22224 -9035 22267 -9001
rect 22296 -9035 22339 -9001
rect 22368 -9029 22412 -9001
rect 22714 -9025 22757 -8991
rect 22759 -9025 22768 -8980
rect 22855 -8992 22862 -8809
rect 22889 -8995 22896 -8812
rect 22368 -9035 22411 -9029
rect 21805 -9088 21848 -9054
rect 21901 -9088 21944 -9054
rect 21997 -9088 22040 -9054
rect 22901 -9076 22910 -8809
rect 23238 -8812 23240 -8742
rect 23272 -8819 23274 -8740
rect 23755 -8741 23769 -8673
rect 23796 -8707 23803 -8639
rect 23841 -8671 23848 -8603
rect 23875 -8637 23882 -8571
rect 23885 -8621 23928 -8587
rect 24086 -8666 24129 -8632
rect 23855 -8689 23864 -8681
rect 23866 -8723 23909 -8689
rect 24086 -8734 24129 -8700
rect 23755 -8753 23764 -8741
rect 24135 -8750 24142 -8616
rect 23530 -8819 23925 -8753
rect 24169 -8784 24176 -8590
rect 24209 -8606 24218 -8595
rect 24205 -8637 24218 -8606
rect 24531 -8624 24574 -8590
rect 22917 -8860 22960 -8826
rect 23266 -8830 23285 -8819
rect 23266 -8832 23274 -8830
rect 22917 -8928 22960 -8894
rect 22969 -8995 22976 -8860
rect 23200 -8874 23274 -8832
rect 23328 -8874 23925 -8819
rect 24064 -8853 24107 -8819
rect 24109 -8853 24118 -8808
rect 24205 -8820 24212 -8637
rect 24239 -8823 24246 -8640
rect 23200 -8877 23925 -8874
rect 23003 -8980 23010 -8892
rect 23120 -8942 23163 -8908
rect 23165 -8942 23174 -8900
rect 23001 -8991 23010 -8980
rect 23003 -9025 23010 -8991
rect 23012 -9025 23055 -8991
rect 23120 -9042 23163 -9008
rect 23165 -9042 23174 -8997
rect 23200 -9044 23353 -8877
rect 23530 -8899 23925 -8877
rect 23454 -8925 23925 -8899
rect 24251 -8904 24260 -8637
rect 24588 -8640 24590 -8570
rect 24267 -8688 24310 -8654
rect 24622 -8674 24624 -8568
rect 24816 -8577 24859 -8543
rect 24861 -8577 24870 -8532
rect 24961 -8543 24970 -8532
rect 25170 -8537 25213 -8503
rect 25215 -8537 25224 -8492
rect 25315 -8503 25324 -8492
rect 25560 -8496 25603 -8462
rect 25605 -8496 25614 -8451
rect 25326 -8537 25369 -8503
rect 24972 -8577 25015 -8543
rect 24267 -8756 24310 -8722
rect 24319 -8823 24326 -8688
rect 24881 -8691 24924 -8657
rect 24933 -8718 24940 -8641
rect 24353 -8808 24360 -8720
rect 24470 -8770 24513 -8736
rect 24515 -8770 24524 -8728
rect 24615 -8740 24624 -8729
rect 24626 -8774 24669 -8740
rect 24967 -8752 24974 -8607
rect 25170 -8620 25213 -8586
rect 25215 -8620 25224 -8575
rect 25315 -8586 25324 -8575
rect 25560 -8580 25603 -8546
rect 25605 -8580 25614 -8535
rect 25326 -8620 25369 -8586
rect 25235 -8734 25278 -8700
rect 25287 -8761 25294 -8684
rect 24351 -8819 24360 -8808
rect 24820 -8813 24863 -8779
rect 24865 -8813 24874 -8771
rect 24965 -8779 24974 -8771
rect 24976 -8813 25019 -8779
rect 25321 -8795 25328 -8650
rect 25560 -8663 25603 -8629
rect 25605 -8663 25614 -8618
rect 25682 -8679 25689 -8413
rect 25716 -8413 25759 -8379
rect 25761 -8413 25775 -8371
rect 25705 -8462 25714 -8451
rect 25716 -8462 25723 -8413
rect 25770 -8451 25775 -8413
rect 25716 -8496 25759 -8462
rect 25761 -8496 25775 -8451
rect 25705 -8546 25714 -8535
rect 25716 -8546 25723 -8496
rect 25770 -8535 25775 -8496
rect 25716 -8580 25759 -8546
rect 25761 -8580 25775 -8535
rect 25705 -8629 25714 -8618
rect 25716 -8629 25723 -8580
rect 25770 -8618 25775 -8580
rect 25716 -8663 25759 -8629
rect 25761 -8663 25775 -8618
rect 25705 -8697 25714 -8671
rect 25716 -8713 25723 -8663
rect 25625 -8777 25668 -8743
rect 25682 -8804 25684 -8727
rect 25716 -8809 25718 -8713
rect 24353 -8853 24360 -8819
rect 24362 -8853 24405 -8819
rect 24470 -8870 24513 -8836
rect 24515 -8870 24524 -8825
rect 24615 -8832 24624 -8821
rect 24626 -8866 24669 -8832
rect 25174 -8856 25217 -8822
rect 25219 -8856 25228 -8814
rect 25319 -8822 25328 -8814
rect 25330 -8856 25373 -8822
rect 25747 -8845 25756 -8697
rect 25770 -8713 25775 -8663
rect 25804 -8679 25809 -8363
rect 25861 -8379 25870 -8371
rect 25810 -8413 25853 -8379
rect 25872 -8413 25925 -8379
rect 26582 -8422 26589 -8406
rect 26605 -8422 26614 -8414
rect 26616 -8422 26623 -8406
rect 26913 -8408 26955 -8374
rect 26958 -8408 26966 -8363
rect 25861 -8462 25870 -8451
rect 26042 -8456 26085 -8422
rect 26114 -8456 26157 -8422
rect 26186 -8456 26229 -8422
rect 26330 -8456 26373 -8422
rect 26402 -8456 26517 -8422
rect 26546 -8456 26589 -8422
rect 25872 -8496 25915 -8462
rect 25861 -8546 25870 -8535
rect 26439 -8539 26482 -8505
rect 25872 -8580 25915 -8546
rect 25861 -8629 25870 -8618
rect 25872 -8663 25915 -8629
rect 26104 -8689 26147 -8655
rect 26149 -8689 26158 -8644
rect 26226 -8706 26233 -8588
rect 26249 -8655 26258 -8644
rect 26260 -8655 26267 -8622
rect 26296 -8655 26303 -8622
rect 26260 -8689 26303 -8655
rect 26305 -8689 26314 -8644
rect 26260 -8740 26267 -8689
rect 26296 -8740 26303 -8689
rect 26330 -8706 26337 -8589
rect 26427 -8630 26429 -8589
rect 26439 -8623 26482 -8589
rect 26439 -8706 26482 -8672
rect 26582 -8706 26589 -8456
rect 26616 -8456 26659 -8422
rect 26605 -8505 26614 -8494
rect 26616 -8505 26623 -8456
rect 26913 -8491 26955 -8457
rect 26958 -8491 26966 -8446
rect 26616 -8539 26659 -8505
rect 26605 -8589 26614 -8578
rect 26616 -8589 26623 -8539
rect 26767 -8565 26875 -8499
rect 27035 -8507 27041 -8241
rect 27069 -8241 27111 -8207
rect 27114 -8241 27122 -8199
rect 27058 -8290 27066 -8279
rect 27069 -8290 27075 -8241
rect 27069 -8324 27111 -8290
rect 27114 -8324 27122 -8279
rect 27058 -8374 27066 -8363
rect 27069 -8374 27075 -8324
rect 27069 -8408 27111 -8374
rect 27114 -8408 27122 -8363
rect 27058 -8457 27066 -8446
rect 27069 -8457 27075 -8408
rect 27069 -8491 27111 -8457
rect 27114 -8491 27122 -8446
rect 27058 -8525 27066 -8499
rect 27069 -8541 27075 -8491
rect 26616 -8623 26659 -8589
rect 26978 -8605 27020 -8571
rect 26605 -8672 26614 -8661
rect 26616 -8672 26623 -8623
rect 27035 -8632 27036 -8555
rect 27069 -8637 27070 -8541
rect 26616 -8706 26659 -8672
rect 27100 -8673 27108 -8525
rect 27123 -8541 27127 -8191
rect 27157 -8507 27161 -8191
rect 27214 -8207 27222 -8199
rect 27163 -8241 27205 -8207
rect 27225 -8241 27277 -8207
rect 28140 -8231 28182 -8197
rect 28236 -8231 28278 -8197
rect 28332 -8231 28374 -8197
rect 30302 -8207 30310 -8199
rect 30379 -8207 30385 -8191
rect 30402 -8207 30410 -8199
rect 30413 -8207 30419 -8191
rect 27933 -8250 27939 -8234
rect 27956 -8250 27964 -8242
rect 27967 -8250 27973 -8234
rect 27214 -8290 27222 -8279
rect 27393 -8284 27435 -8250
rect 27465 -8284 27507 -8250
rect 27537 -8284 27579 -8250
rect 27681 -8284 27723 -8250
rect 27753 -8284 27867 -8250
rect 27897 -8284 27939 -8250
rect 27225 -8324 27267 -8290
rect 27214 -8374 27222 -8363
rect 27790 -8367 27832 -8333
rect 27225 -8408 27267 -8374
rect 27214 -8457 27222 -8446
rect 27225 -8491 27267 -8457
rect 27455 -8517 27497 -8483
rect 27500 -8517 27508 -8472
rect 27577 -8534 27583 -8416
rect 27600 -8483 27608 -8472
rect 27611 -8483 27617 -8450
rect 27647 -8483 27653 -8450
rect 27611 -8517 27653 -8483
rect 27656 -8517 27664 -8472
rect 27611 -8568 27617 -8517
rect 27647 -8568 27653 -8517
rect 27681 -8534 27687 -8417
rect 27778 -8458 27779 -8417
rect 27790 -8451 27832 -8417
rect 27790 -8534 27832 -8500
rect 27933 -8534 27939 -8284
rect 27967 -8284 28009 -8250
rect 28494 -8274 28536 -8240
rect 28590 -8274 28632 -8240
rect 28686 -8274 28728 -8240
rect 30193 -8241 30235 -8207
rect 30257 -8241 30310 -8207
rect 30337 -8241 30385 -8207
rect 27956 -8333 27964 -8322
rect 27967 -8333 27973 -8284
rect 28206 -8293 28214 -8285
rect 28306 -8293 28314 -8285
rect 28133 -8327 28203 -8293
rect 28205 -8327 28247 -8293
rect 28317 -8327 28359 -8293
rect 28848 -8317 28890 -8283
rect 28944 -8317 28986 -8283
rect 29040 -8317 29082 -8283
rect 29136 -8317 29178 -8283
rect 29232 -8317 29274 -8283
rect 30257 -8324 30299 -8290
rect 30302 -8324 30310 -8279
rect 27967 -8367 28009 -8333
rect 28560 -8336 28568 -8328
rect 28660 -8336 28668 -8328
rect 27956 -8417 27964 -8406
rect 27967 -8417 27973 -8367
rect 28161 -8410 28203 -8376
rect 28206 -8410 28214 -8365
rect 28306 -8376 28314 -8365
rect 28487 -8370 28557 -8336
rect 28559 -8370 28601 -8336
rect 28671 -8370 28713 -8336
rect 29396 -8360 29438 -8326
rect 29492 -8360 29534 -8326
rect 29588 -8360 29630 -8326
rect 29684 -8360 29726 -8326
rect 29780 -8360 29822 -8326
rect 29876 -8360 29918 -8326
rect 29972 -8360 30014 -8326
rect 28317 -8410 28359 -8376
rect 28950 -8379 28958 -8371
rect 29027 -8379 29033 -8363
rect 29050 -8379 29058 -8371
rect 29061 -8379 29067 -8363
rect 27967 -8451 28009 -8417
rect 27956 -8500 27964 -8489
rect 27967 -8500 27973 -8451
rect 28161 -8494 28203 -8460
rect 28206 -8494 28214 -8449
rect 28306 -8460 28314 -8449
rect 28515 -8453 28557 -8419
rect 28560 -8453 28568 -8408
rect 28660 -8419 28668 -8408
rect 28841 -8413 28883 -8379
rect 28905 -8413 28958 -8379
rect 28985 -8413 29033 -8379
rect 28671 -8453 28713 -8419
rect 28317 -8494 28359 -8460
rect 27967 -8534 28009 -8500
rect 27967 -8568 27973 -8534
rect 26616 -8740 26623 -8706
rect 26913 -8723 26955 -8689
rect 26958 -8723 26966 -8681
rect 24363 -8906 24406 -8872
rect 24435 -8906 24478 -8872
rect 24507 -8906 24550 -8872
rect 24820 -8913 24863 -8879
rect 24865 -8913 24874 -8868
rect 24965 -8879 24974 -8868
rect 24976 -8913 25019 -8879
rect 25560 -8895 25603 -8861
rect 25605 -8895 25614 -8853
rect 23454 -8959 23938 -8925
rect 24788 -8949 24831 -8915
rect 24860 -8949 24903 -8915
rect 25174 -8956 25217 -8922
rect 25219 -8956 25228 -8911
rect 25319 -8922 25328 -8911
rect 25747 -8913 25761 -8845
rect 25788 -8879 25795 -8811
rect 25833 -8843 25840 -8775
rect 25867 -8809 25874 -8743
rect 25877 -8793 25920 -8759
rect 26080 -8838 26123 -8804
rect 25847 -8861 25856 -8853
rect 25858 -8895 25901 -8861
rect 26080 -8906 26123 -8872
rect 25330 -8956 25373 -8922
rect 23454 -8985 23925 -8959
rect 23458 -8993 23667 -8985
rect 23474 -9003 23651 -8993
rect 23013 -9078 23056 -9044
rect 23085 -9078 23128 -9044
rect 23157 -9078 23353 -9044
rect 22159 -9131 22202 -9097
rect 22255 -9131 22298 -9097
rect 22351 -9131 22394 -9097
rect 22447 -9131 22490 -9097
rect 22543 -9131 22586 -9097
rect 23200 -9114 23353 -9078
rect 23200 -9140 23383 -9114
rect 22707 -9174 22750 -9140
rect 22803 -9174 22846 -9140
rect 22899 -9174 22942 -9140
rect 22995 -9174 23038 -9140
rect 23091 -9174 23134 -9140
rect 23187 -9174 23383 -9140
rect 23200 -9200 23383 -9174
rect 23400 -9174 23509 -9050
rect 23659 -9062 23667 -9051
rect 23278 -9870 23321 -9200
rect 23400 -9228 23411 -9174
rect 22753 -9970 23130 -9936
rect 23212 -9971 23238 -9924
rect 23266 -9971 23321 -9870
rect 23412 -9971 23455 -9174
rect 23458 -9971 23466 -9174
rect 23670 -9971 23713 -9062
rect 23804 -9971 23847 -8985
rect 24057 -9002 24100 -8968
rect 24153 -9002 24196 -8968
rect 24249 -9002 24292 -8968
rect 24345 -9002 24388 -8968
rect 24441 -9002 24484 -8968
rect 24537 -9002 24580 -8968
rect 24633 -9002 24676 -8968
rect 25142 -8992 25185 -8958
rect 25214 -8992 25257 -8958
rect 25560 -8995 25603 -8961
rect 25605 -8995 25614 -8950
rect 25747 -9001 25756 -8913
rect 26129 -8922 26136 -8788
rect 25847 -8961 25856 -8950
rect 26163 -8956 26170 -8762
rect 26203 -8778 26212 -8767
rect 26199 -8809 26212 -8778
rect 26525 -8796 26568 -8762
rect 25858 -8995 25901 -8961
rect 24795 -9045 24838 -9011
rect 24891 -9045 24934 -9011
rect 24987 -9045 25030 -9011
rect 25496 -9035 25539 -9001
rect 25568 -9035 25611 -9001
rect 25640 -9035 25683 -9001
rect 25712 -9029 25756 -9001
rect 26058 -9025 26101 -8991
rect 26103 -9025 26112 -8980
rect 26199 -8992 26206 -8809
rect 26233 -8995 26240 -8812
rect 25712 -9035 25755 -9029
rect 25149 -9088 25192 -9054
rect 25245 -9088 25288 -9054
rect 25341 -9088 25384 -9054
rect 26245 -9076 26254 -8809
rect 26582 -8812 26584 -8742
rect 26616 -8819 26618 -8740
rect 27100 -8741 27113 -8673
rect 27141 -8707 27147 -8639
rect 27186 -8671 27192 -8603
rect 27220 -8637 27226 -8571
rect 27230 -8621 27272 -8587
rect 27431 -8666 27473 -8632
rect 27200 -8689 27208 -8681
rect 27211 -8723 27253 -8689
rect 27431 -8734 27473 -8700
rect 27100 -8753 27108 -8741
rect 27480 -8750 27486 -8616
rect 26875 -8819 27269 -8753
rect 27514 -8784 27520 -8590
rect 27554 -8606 27562 -8595
rect 27550 -8637 27562 -8606
rect 27876 -8624 27918 -8590
rect 26261 -8860 26304 -8826
rect 26610 -8830 26629 -8819
rect 26610 -8832 26618 -8830
rect 26261 -8928 26304 -8894
rect 26313 -8995 26320 -8860
rect 26544 -8874 26618 -8832
rect 26673 -8874 27269 -8819
rect 27409 -8853 27451 -8819
rect 27454 -8853 27462 -8808
rect 27550 -8820 27556 -8637
rect 27584 -8823 27590 -8640
rect 26544 -8877 27269 -8874
rect 26347 -8980 26354 -8892
rect 26464 -8942 26507 -8908
rect 26509 -8942 26518 -8900
rect 26345 -8991 26354 -8980
rect 26347 -9025 26354 -8991
rect 26356 -9025 26399 -8991
rect 26464 -9042 26507 -9008
rect 26509 -9042 26518 -8997
rect 26544 -9044 26697 -8877
rect 26875 -8899 27269 -8877
rect 26799 -8925 27269 -8899
rect 27596 -8904 27604 -8637
rect 27933 -8640 27934 -8570
rect 27612 -8688 27654 -8654
rect 27967 -8674 27968 -8568
rect 28161 -8577 28203 -8543
rect 28206 -8577 28214 -8532
rect 28306 -8543 28314 -8532
rect 28515 -8537 28557 -8503
rect 28560 -8537 28568 -8492
rect 28660 -8503 28668 -8492
rect 28905 -8496 28947 -8462
rect 28950 -8496 28958 -8451
rect 28671 -8537 28713 -8503
rect 28317 -8577 28359 -8543
rect 27612 -8756 27654 -8722
rect 27664 -8823 27670 -8688
rect 28226 -8691 28268 -8657
rect 28278 -8718 28284 -8641
rect 27698 -8808 27704 -8720
rect 27815 -8770 27857 -8736
rect 27860 -8770 27868 -8728
rect 27960 -8740 27968 -8729
rect 27971 -8774 28013 -8740
rect 28312 -8752 28318 -8607
rect 28515 -8620 28557 -8586
rect 28560 -8620 28568 -8575
rect 28660 -8586 28668 -8575
rect 28905 -8580 28947 -8546
rect 28950 -8580 28958 -8535
rect 28671 -8620 28713 -8586
rect 28580 -8734 28622 -8700
rect 28632 -8761 28638 -8684
rect 27696 -8819 27704 -8808
rect 28165 -8813 28207 -8779
rect 28210 -8813 28218 -8771
rect 28310 -8779 28318 -8771
rect 28321 -8813 28363 -8779
rect 28666 -8795 28672 -8650
rect 28905 -8663 28947 -8629
rect 28950 -8663 28958 -8618
rect 29027 -8679 29033 -8413
rect 29061 -8413 29103 -8379
rect 29106 -8413 29114 -8371
rect 29050 -8462 29058 -8451
rect 29061 -8462 29067 -8413
rect 29061 -8496 29103 -8462
rect 29106 -8496 29114 -8451
rect 29050 -8546 29058 -8535
rect 29061 -8546 29067 -8496
rect 29061 -8580 29103 -8546
rect 29106 -8580 29114 -8535
rect 29050 -8629 29058 -8618
rect 29061 -8629 29067 -8580
rect 29061 -8663 29103 -8629
rect 29106 -8663 29114 -8618
rect 29050 -8697 29058 -8671
rect 29061 -8713 29067 -8663
rect 28970 -8777 29012 -8743
rect 29027 -8804 29028 -8727
rect 29061 -8809 29062 -8713
rect 27698 -8853 27704 -8819
rect 27707 -8853 27749 -8819
rect 27815 -8870 27857 -8836
rect 27860 -8870 27868 -8825
rect 27960 -8832 27968 -8821
rect 27971 -8866 28013 -8832
rect 28519 -8856 28561 -8822
rect 28564 -8856 28572 -8814
rect 28664 -8822 28672 -8814
rect 28675 -8856 28717 -8822
rect 29092 -8845 29100 -8697
rect 29115 -8713 29119 -8363
rect 29149 -8679 29153 -8363
rect 29206 -8379 29214 -8371
rect 29155 -8413 29197 -8379
rect 29217 -8413 29269 -8379
rect 29927 -8422 29933 -8406
rect 29950 -8422 29958 -8414
rect 29961 -8422 29967 -8406
rect 30257 -8408 30299 -8374
rect 30302 -8408 30310 -8363
rect 29206 -8462 29214 -8451
rect 29387 -8456 29429 -8422
rect 29459 -8456 29501 -8422
rect 29531 -8456 29573 -8422
rect 29675 -8456 29717 -8422
rect 29747 -8456 29861 -8422
rect 29891 -8456 29933 -8422
rect 29217 -8496 29259 -8462
rect 29206 -8546 29214 -8535
rect 29784 -8539 29826 -8505
rect 29217 -8580 29259 -8546
rect 29206 -8629 29214 -8618
rect 29217 -8663 29259 -8629
rect 29449 -8689 29491 -8655
rect 29494 -8689 29502 -8644
rect 29571 -8706 29577 -8588
rect 29594 -8655 29602 -8644
rect 29605 -8655 29611 -8622
rect 29641 -8655 29647 -8622
rect 29605 -8689 29647 -8655
rect 29650 -8689 29658 -8644
rect 29605 -8740 29611 -8689
rect 29641 -8740 29647 -8689
rect 29675 -8706 29681 -8589
rect 29772 -8630 29773 -8589
rect 29784 -8623 29826 -8589
rect 29784 -8706 29826 -8672
rect 29927 -8706 29933 -8456
rect 29961 -8456 30003 -8422
rect 29950 -8505 29958 -8494
rect 29961 -8505 29967 -8456
rect 30257 -8491 30299 -8457
rect 30302 -8491 30310 -8446
rect 29961 -8539 30003 -8505
rect 29950 -8589 29958 -8578
rect 29961 -8589 29967 -8539
rect 30111 -8565 30219 -8499
rect 30379 -8507 30385 -8241
rect 30413 -8241 30455 -8207
rect 30458 -8241 30466 -8199
rect 30402 -8290 30410 -8279
rect 30413 -8290 30419 -8241
rect 30413 -8324 30455 -8290
rect 30458 -8324 30466 -8279
rect 30402 -8374 30410 -8363
rect 30413 -8374 30419 -8324
rect 30413 -8408 30455 -8374
rect 30458 -8408 30466 -8363
rect 30402 -8457 30410 -8446
rect 30413 -8457 30419 -8408
rect 30413 -8491 30455 -8457
rect 30458 -8491 30466 -8446
rect 30402 -8525 30410 -8499
rect 30413 -8541 30419 -8491
rect 29961 -8623 30003 -8589
rect 30322 -8605 30364 -8571
rect 29950 -8672 29958 -8661
rect 29961 -8672 29967 -8623
rect 30379 -8632 30380 -8555
rect 30413 -8637 30414 -8541
rect 29961 -8706 30003 -8672
rect 30444 -8673 30452 -8525
rect 30467 -8541 30471 -8191
rect 30501 -8507 30505 -8191
rect 30558 -8207 30566 -8199
rect 30507 -8241 30549 -8207
rect 30569 -8241 30621 -8207
rect 31484 -8231 31526 -8197
rect 31580 -8231 31622 -8197
rect 31676 -8231 31718 -8197
rect 33646 -8207 33654 -8199
rect 33723 -8207 33729 -8191
rect 33746 -8207 33754 -8199
rect 33757 -8207 33763 -8191
rect 31277 -8250 31283 -8234
rect 31300 -8250 31308 -8242
rect 31311 -8250 31317 -8234
rect 30558 -8290 30566 -8279
rect 30737 -8284 30779 -8250
rect 30809 -8284 30851 -8250
rect 30881 -8284 30923 -8250
rect 31025 -8284 31067 -8250
rect 31097 -8284 31211 -8250
rect 31241 -8284 31283 -8250
rect 30569 -8324 30611 -8290
rect 30558 -8374 30566 -8363
rect 31134 -8367 31176 -8333
rect 30569 -8408 30611 -8374
rect 30558 -8457 30566 -8446
rect 30569 -8491 30611 -8457
rect 30799 -8517 30841 -8483
rect 30844 -8517 30852 -8472
rect 30921 -8534 30927 -8416
rect 30944 -8483 30952 -8472
rect 30955 -8483 30961 -8450
rect 30991 -8483 30997 -8450
rect 30955 -8517 30997 -8483
rect 31000 -8517 31008 -8472
rect 30955 -8568 30961 -8517
rect 30991 -8568 30997 -8517
rect 31025 -8534 31031 -8417
rect 31122 -8458 31123 -8417
rect 31134 -8451 31176 -8417
rect 31134 -8534 31176 -8500
rect 31277 -8534 31283 -8284
rect 31311 -8284 31353 -8250
rect 31838 -8274 31880 -8240
rect 31934 -8274 31976 -8240
rect 32030 -8274 32072 -8240
rect 33537 -8241 33579 -8207
rect 33601 -8241 33654 -8207
rect 33681 -8241 33729 -8207
rect 31300 -8333 31308 -8322
rect 31311 -8333 31317 -8284
rect 31550 -8293 31558 -8285
rect 31650 -8293 31658 -8285
rect 31477 -8327 31547 -8293
rect 31549 -8327 31591 -8293
rect 31661 -8327 31703 -8293
rect 32192 -8317 32234 -8283
rect 32288 -8317 32330 -8283
rect 32384 -8317 32426 -8283
rect 32480 -8317 32522 -8283
rect 32576 -8317 32618 -8283
rect 33601 -8324 33643 -8290
rect 33646 -8324 33654 -8279
rect 31311 -8367 31353 -8333
rect 31904 -8336 31912 -8328
rect 32004 -8336 32012 -8328
rect 31300 -8417 31308 -8406
rect 31311 -8417 31317 -8367
rect 31505 -8410 31547 -8376
rect 31550 -8410 31558 -8365
rect 31650 -8376 31658 -8365
rect 31831 -8370 31901 -8336
rect 31903 -8370 31945 -8336
rect 32015 -8370 32057 -8336
rect 32740 -8360 32782 -8326
rect 32836 -8360 32878 -8326
rect 32932 -8360 32974 -8326
rect 33028 -8360 33070 -8326
rect 33124 -8360 33166 -8326
rect 33220 -8360 33262 -8326
rect 33316 -8360 33358 -8326
rect 31661 -8410 31703 -8376
rect 32294 -8379 32302 -8371
rect 32371 -8379 32377 -8363
rect 32394 -8379 32402 -8371
rect 32405 -8379 32411 -8363
rect 31311 -8451 31353 -8417
rect 31300 -8500 31308 -8489
rect 31311 -8500 31317 -8451
rect 31505 -8494 31547 -8460
rect 31550 -8494 31558 -8449
rect 31650 -8460 31658 -8449
rect 31859 -8453 31901 -8419
rect 31904 -8453 31912 -8408
rect 32004 -8419 32012 -8408
rect 32185 -8413 32227 -8379
rect 32249 -8413 32302 -8379
rect 32329 -8413 32377 -8379
rect 32015 -8453 32057 -8419
rect 31661 -8494 31703 -8460
rect 31311 -8534 31353 -8500
rect 31311 -8568 31317 -8534
rect 29961 -8740 29967 -8706
rect 30257 -8723 30299 -8689
rect 30302 -8723 30310 -8681
rect 27708 -8906 27750 -8872
rect 27780 -8906 27822 -8872
rect 27852 -8906 27894 -8872
rect 28165 -8913 28207 -8879
rect 28210 -8913 28218 -8868
rect 28310 -8879 28318 -8868
rect 28321 -8913 28363 -8879
rect 28905 -8895 28947 -8861
rect 28950 -8895 28958 -8853
rect 26799 -8959 27282 -8925
rect 28133 -8949 28175 -8915
rect 28205 -8949 28247 -8915
rect 28519 -8956 28561 -8922
rect 28564 -8956 28572 -8911
rect 28664 -8922 28672 -8911
rect 29092 -8913 29105 -8845
rect 29133 -8879 29139 -8811
rect 29178 -8843 29184 -8775
rect 29212 -8809 29218 -8743
rect 29222 -8793 29264 -8759
rect 29425 -8838 29467 -8804
rect 29192 -8861 29200 -8853
rect 29203 -8895 29245 -8861
rect 29425 -8906 29467 -8872
rect 28675 -8956 28717 -8922
rect 26799 -8985 27269 -8959
rect 26802 -8993 27011 -8985
rect 26818 -9003 26995 -8993
rect 26357 -9078 26400 -9044
rect 26429 -9078 26472 -9044
rect 26501 -9078 26697 -9044
rect 25503 -9131 25546 -9097
rect 25599 -9131 25642 -9097
rect 25695 -9131 25738 -9097
rect 25791 -9131 25834 -9097
rect 25887 -9131 25930 -9097
rect 26544 -9114 26697 -9078
rect 26544 -9140 26727 -9114
rect 26051 -9174 26094 -9140
rect 26147 -9174 26190 -9140
rect 26243 -9174 26286 -9140
rect 26339 -9174 26382 -9140
rect 26435 -9174 26478 -9140
rect 26531 -9174 26727 -9140
rect 26544 -9200 26727 -9174
rect 26744 -9174 26853 -9050
rect 27003 -9062 27011 -9051
rect 26622 -9870 26665 -9200
rect 26744 -9228 26755 -9174
rect 26097 -9970 26474 -9936
rect 26556 -9971 26582 -9924
rect 26610 -9971 26665 -9870
rect 26756 -9971 26799 -9174
rect 26802 -9971 26810 -9174
rect 27014 -9971 27057 -9062
rect 27148 -9971 27191 -8985
rect 27402 -9002 27444 -8968
rect 27498 -9002 27540 -8968
rect 27594 -9002 27636 -8968
rect 27690 -9002 27732 -8968
rect 27786 -9002 27828 -8968
rect 27882 -9002 27924 -8968
rect 27978 -9002 28020 -8968
rect 28487 -8992 28529 -8958
rect 28559 -8992 28601 -8958
rect 28905 -8995 28947 -8961
rect 28950 -8995 28958 -8950
rect 29092 -9001 29100 -8913
rect 29474 -8922 29480 -8788
rect 29192 -8961 29200 -8950
rect 29508 -8956 29514 -8762
rect 29548 -8778 29556 -8767
rect 29544 -8809 29556 -8778
rect 29870 -8796 29912 -8762
rect 29203 -8995 29245 -8961
rect 28140 -9045 28182 -9011
rect 28236 -9045 28278 -9011
rect 28332 -9045 28374 -9011
rect 28841 -9035 28883 -9001
rect 28913 -9035 28955 -9001
rect 28985 -9035 29027 -9001
rect 29057 -9029 29100 -9001
rect 29403 -9025 29445 -8991
rect 29448 -9025 29456 -8980
rect 29544 -8992 29550 -8809
rect 29578 -8995 29584 -8812
rect 29057 -9035 29099 -9029
rect 28494 -9088 28536 -9054
rect 28590 -9088 28632 -9054
rect 28686 -9088 28728 -9054
rect 29590 -9076 29598 -8809
rect 29927 -8812 29928 -8742
rect 29961 -8819 29962 -8740
rect 30444 -8741 30457 -8673
rect 30485 -8707 30491 -8639
rect 30530 -8671 30536 -8603
rect 30564 -8637 30570 -8571
rect 30574 -8621 30616 -8587
rect 30775 -8666 30817 -8632
rect 30544 -8689 30552 -8681
rect 30555 -8723 30597 -8689
rect 30775 -8734 30817 -8700
rect 30444 -8753 30452 -8741
rect 30824 -8750 30830 -8616
rect 30219 -8819 30613 -8753
rect 30858 -8784 30864 -8590
rect 30898 -8606 30906 -8595
rect 30894 -8637 30906 -8606
rect 31220 -8624 31262 -8590
rect 29606 -8860 29648 -8826
rect 29955 -8830 29973 -8819
rect 29955 -8832 29962 -8830
rect 29606 -8928 29648 -8894
rect 29658 -8995 29664 -8860
rect 29889 -8874 29962 -8832
rect 30017 -8874 30613 -8819
rect 30753 -8853 30795 -8819
rect 30798 -8853 30806 -8808
rect 30894 -8820 30900 -8637
rect 30928 -8823 30934 -8640
rect 29889 -8877 30613 -8874
rect 29692 -8980 29698 -8892
rect 29809 -8942 29851 -8908
rect 29854 -8942 29862 -8900
rect 29690 -8991 29698 -8980
rect 29692 -9025 29698 -8991
rect 29701 -9025 29743 -8991
rect 29809 -9042 29851 -9008
rect 29854 -9042 29862 -8997
rect 29702 -9078 29744 -9044
rect 29774 -9078 29816 -9044
rect 29846 -9078 29888 -9044
rect 28848 -9131 28890 -9097
rect 28944 -9131 28986 -9097
rect 29040 -9131 29082 -9097
rect 29136 -9131 29178 -9097
rect 29232 -9131 29274 -9097
rect 29889 -9114 30041 -8877
rect 30219 -8899 30613 -8877
rect 30143 -8925 30613 -8899
rect 30940 -8904 30948 -8637
rect 31277 -8640 31278 -8570
rect 30956 -8688 30998 -8654
rect 31311 -8674 31312 -8568
rect 31505 -8577 31547 -8543
rect 31550 -8577 31558 -8532
rect 31650 -8543 31658 -8532
rect 31859 -8537 31901 -8503
rect 31904 -8537 31912 -8492
rect 32004 -8503 32012 -8492
rect 32249 -8496 32291 -8462
rect 32294 -8496 32302 -8451
rect 32015 -8537 32057 -8503
rect 31661 -8577 31703 -8543
rect 30956 -8756 30998 -8722
rect 31008 -8823 31014 -8688
rect 31570 -8691 31612 -8657
rect 31622 -8718 31628 -8641
rect 31042 -8808 31048 -8720
rect 31159 -8770 31201 -8736
rect 31204 -8770 31212 -8728
rect 31304 -8740 31312 -8729
rect 31315 -8774 31357 -8740
rect 31656 -8752 31662 -8607
rect 31859 -8620 31901 -8586
rect 31904 -8620 31912 -8575
rect 32004 -8586 32012 -8575
rect 32249 -8580 32291 -8546
rect 32294 -8580 32302 -8535
rect 32015 -8620 32057 -8586
rect 31924 -8734 31966 -8700
rect 31976 -8761 31982 -8684
rect 31040 -8819 31048 -8808
rect 31509 -8813 31551 -8779
rect 31554 -8813 31562 -8771
rect 31654 -8779 31662 -8771
rect 31665 -8813 31707 -8779
rect 32010 -8795 32016 -8650
rect 32249 -8663 32291 -8629
rect 32294 -8663 32302 -8618
rect 32371 -8679 32377 -8413
rect 32405 -8413 32447 -8379
rect 32450 -8413 32458 -8371
rect 32394 -8462 32402 -8451
rect 32405 -8462 32411 -8413
rect 32405 -8496 32447 -8462
rect 32450 -8496 32458 -8451
rect 32394 -8546 32402 -8535
rect 32405 -8546 32411 -8496
rect 32405 -8580 32447 -8546
rect 32450 -8580 32458 -8535
rect 32394 -8629 32402 -8618
rect 32405 -8629 32411 -8580
rect 32405 -8663 32447 -8629
rect 32450 -8663 32458 -8618
rect 32394 -8697 32402 -8671
rect 32405 -8713 32411 -8663
rect 32314 -8777 32356 -8743
rect 32371 -8804 32372 -8727
rect 32405 -8809 32406 -8713
rect 31042 -8853 31048 -8819
rect 31051 -8853 31093 -8819
rect 31159 -8870 31201 -8836
rect 31204 -8870 31212 -8825
rect 31304 -8832 31312 -8821
rect 31315 -8866 31357 -8832
rect 31863 -8856 31905 -8822
rect 31908 -8856 31916 -8814
rect 32008 -8822 32016 -8814
rect 32019 -8856 32061 -8822
rect 32436 -8845 32444 -8697
rect 32459 -8713 32463 -8363
rect 32493 -8679 32497 -8363
rect 32550 -8379 32558 -8371
rect 32499 -8413 32541 -8379
rect 32561 -8413 32613 -8379
rect 33271 -8422 33277 -8406
rect 33294 -8422 33302 -8414
rect 33305 -8422 33311 -8406
rect 33601 -8408 33643 -8374
rect 33646 -8408 33654 -8363
rect 32550 -8462 32558 -8451
rect 32731 -8456 32773 -8422
rect 32803 -8456 32845 -8422
rect 32875 -8456 32917 -8422
rect 33019 -8456 33061 -8422
rect 33091 -8456 33205 -8422
rect 33235 -8456 33277 -8422
rect 32561 -8496 32603 -8462
rect 32550 -8546 32558 -8535
rect 33128 -8539 33170 -8505
rect 32561 -8580 32603 -8546
rect 32550 -8629 32558 -8618
rect 32561 -8663 32603 -8629
rect 32793 -8689 32835 -8655
rect 32838 -8689 32846 -8644
rect 32915 -8706 32921 -8588
rect 32938 -8655 32946 -8644
rect 32949 -8655 32955 -8622
rect 32985 -8655 32991 -8622
rect 32949 -8689 32991 -8655
rect 32994 -8689 33002 -8644
rect 32949 -8740 32955 -8689
rect 32985 -8740 32991 -8689
rect 33019 -8706 33025 -8589
rect 33116 -8630 33117 -8589
rect 33128 -8623 33170 -8589
rect 33128 -8706 33170 -8672
rect 33271 -8706 33277 -8456
rect 33305 -8456 33347 -8422
rect 33294 -8505 33302 -8494
rect 33305 -8505 33311 -8456
rect 33601 -8491 33643 -8457
rect 33646 -8491 33654 -8446
rect 33305 -8539 33347 -8505
rect 33294 -8589 33302 -8578
rect 33305 -8589 33311 -8539
rect 33455 -8565 33563 -8499
rect 33723 -8507 33729 -8241
rect 33757 -8241 33799 -8207
rect 33802 -8241 33810 -8199
rect 33746 -8290 33754 -8279
rect 33757 -8290 33763 -8241
rect 33757 -8324 33799 -8290
rect 33802 -8324 33810 -8279
rect 33746 -8374 33754 -8363
rect 33757 -8374 33763 -8324
rect 33757 -8408 33799 -8374
rect 33802 -8408 33810 -8363
rect 33746 -8457 33754 -8446
rect 33757 -8457 33763 -8408
rect 33757 -8491 33799 -8457
rect 33802 -8491 33810 -8446
rect 33746 -8525 33754 -8499
rect 33757 -8541 33763 -8491
rect 33305 -8623 33347 -8589
rect 33666 -8605 33708 -8571
rect 33294 -8672 33302 -8661
rect 33305 -8672 33311 -8623
rect 33723 -8632 33724 -8555
rect 33757 -8637 33758 -8541
rect 33305 -8706 33347 -8672
rect 33788 -8673 33796 -8525
rect 33811 -8541 33815 -8191
rect 33845 -8507 33849 -8191
rect 33902 -8207 33910 -8199
rect 33851 -8241 33893 -8207
rect 33913 -8241 33965 -8207
rect 34828 -8231 34870 -8197
rect 34924 -8231 34966 -8197
rect 35020 -8231 35062 -8197
rect 36990 -8207 36998 -8199
rect 37067 -8207 37073 -8191
rect 37090 -8207 37098 -8199
rect 37101 -8207 37107 -8191
rect 34621 -8250 34627 -8234
rect 34644 -8250 34652 -8242
rect 34655 -8250 34661 -8234
rect 33902 -8290 33910 -8279
rect 34081 -8284 34123 -8250
rect 34153 -8284 34195 -8250
rect 34225 -8284 34267 -8250
rect 34369 -8284 34411 -8250
rect 34441 -8284 34555 -8250
rect 34585 -8284 34627 -8250
rect 33913 -8324 33955 -8290
rect 33902 -8374 33910 -8363
rect 34478 -8367 34520 -8333
rect 33913 -8408 33955 -8374
rect 33902 -8457 33910 -8446
rect 33913 -8491 33955 -8457
rect 34143 -8517 34185 -8483
rect 34188 -8517 34196 -8472
rect 34265 -8534 34271 -8416
rect 34288 -8483 34296 -8472
rect 34299 -8483 34305 -8450
rect 34335 -8483 34341 -8450
rect 34299 -8517 34341 -8483
rect 34344 -8517 34352 -8472
rect 34299 -8568 34305 -8517
rect 34335 -8568 34341 -8517
rect 34369 -8534 34375 -8417
rect 34466 -8458 34467 -8417
rect 34478 -8451 34520 -8417
rect 34478 -8534 34520 -8500
rect 34621 -8534 34627 -8284
rect 34655 -8284 34697 -8250
rect 35182 -8274 35224 -8240
rect 35278 -8274 35320 -8240
rect 35374 -8274 35416 -8240
rect 36881 -8241 36923 -8207
rect 36945 -8241 36998 -8207
rect 37025 -8241 37073 -8207
rect 34644 -8333 34652 -8322
rect 34655 -8333 34661 -8284
rect 34894 -8293 34902 -8285
rect 34994 -8293 35002 -8285
rect 34821 -8327 34891 -8293
rect 34893 -8327 34935 -8293
rect 35005 -8327 35047 -8293
rect 35536 -8317 35578 -8283
rect 35632 -8317 35674 -8283
rect 35728 -8317 35770 -8283
rect 35824 -8317 35866 -8283
rect 35920 -8317 35962 -8283
rect 36945 -8324 36987 -8290
rect 36990 -8324 36998 -8279
rect 34655 -8367 34697 -8333
rect 35248 -8336 35256 -8328
rect 35348 -8336 35356 -8328
rect 34644 -8417 34652 -8406
rect 34655 -8417 34661 -8367
rect 34849 -8410 34891 -8376
rect 34894 -8410 34902 -8365
rect 34994 -8376 35002 -8365
rect 35175 -8370 35245 -8336
rect 35247 -8370 35289 -8336
rect 35359 -8370 35401 -8336
rect 36084 -8360 36126 -8326
rect 36180 -8360 36222 -8326
rect 36276 -8360 36318 -8326
rect 36372 -8360 36414 -8326
rect 36468 -8360 36510 -8326
rect 36564 -8360 36606 -8326
rect 36660 -8360 36702 -8326
rect 35005 -8410 35047 -8376
rect 35638 -8379 35646 -8371
rect 35715 -8379 35721 -8363
rect 35738 -8379 35746 -8371
rect 35749 -8379 35755 -8363
rect 34655 -8451 34697 -8417
rect 34644 -8500 34652 -8489
rect 34655 -8500 34661 -8451
rect 34849 -8494 34891 -8460
rect 34894 -8494 34902 -8449
rect 34994 -8460 35002 -8449
rect 35203 -8453 35245 -8419
rect 35248 -8453 35256 -8408
rect 35348 -8419 35356 -8408
rect 35529 -8413 35571 -8379
rect 35593 -8413 35646 -8379
rect 35673 -8413 35721 -8379
rect 35359 -8453 35401 -8419
rect 35005 -8494 35047 -8460
rect 34655 -8534 34697 -8500
rect 34655 -8568 34661 -8534
rect 33305 -8740 33311 -8706
rect 33601 -8723 33643 -8689
rect 33646 -8723 33654 -8681
rect 31052 -8906 31094 -8872
rect 31124 -8906 31166 -8872
rect 31196 -8906 31238 -8872
rect 31509 -8913 31551 -8879
rect 31554 -8913 31562 -8868
rect 31654 -8879 31662 -8868
rect 31665 -8913 31707 -8879
rect 32249 -8895 32291 -8861
rect 32294 -8895 32302 -8853
rect 30143 -8959 30626 -8925
rect 31477 -8949 31519 -8915
rect 31549 -8949 31591 -8915
rect 31863 -8956 31905 -8922
rect 31908 -8956 31916 -8911
rect 32008 -8922 32016 -8911
rect 32436 -8913 32449 -8845
rect 32477 -8879 32483 -8811
rect 32522 -8843 32528 -8775
rect 32556 -8809 32562 -8743
rect 32566 -8793 32608 -8759
rect 32769 -8838 32811 -8804
rect 32536 -8861 32544 -8853
rect 32547 -8895 32589 -8861
rect 32769 -8906 32811 -8872
rect 32019 -8956 32061 -8922
rect 30143 -8985 30613 -8959
rect 30147 -8993 30355 -8985
rect 30163 -9003 30339 -8993
rect 29889 -9140 30071 -9114
rect 29396 -9174 29438 -9140
rect 29492 -9174 29534 -9140
rect 29588 -9174 29630 -9140
rect 29684 -9174 29726 -9140
rect 29780 -9174 29822 -9140
rect 29876 -9174 30071 -9140
rect 29889 -9200 30071 -9174
rect 30089 -9174 30197 -9050
rect 30348 -9062 30355 -9051
rect 29967 -9870 30009 -9200
rect 30089 -9228 30099 -9174
rect 29774 -9936 29926 -9924
rect 29442 -9970 29926 -9936
rect 29774 -9971 29926 -9970
rect 29955 -9971 30009 -9870
rect 30101 -9971 30143 -9174
rect 30147 -9971 30154 -9174
rect 30359 -9971 30401 -9062
rect 30493 -9971 30535 -8985
rect 30746 -9002 30788 -8968
rect 30842 -9002 30884 -8968
rect 30938 -9002 30980 -8968
rect 31034 -9002 31076 -8968
rect 31130 -9002 31172 -8968
rect 31226 -9002 31268 -8968
rect 31322 -9002 31364 -8968
rect 31831 -8992 31873 -8958
rect 31903 -8992 31945 -8958
rect 32249 -8995 32291 -8961
rect 32294 -8995 32302 -8950
rect 32436 -9001 32444 -8913
rect 32818 -8922 32824 -8788
rect 32536 -8961 32544 -8950
rect 32852 -8956 32858 -8762
rect 32892 -8778 32900 -8767
rect 32888 -8809 32900 -8778
rect 33214 -8796 33256 -8762
rect 32547 -8995 32589 -8961
rect 31484 -9045 31526 -9011
rect 31580 -9045 31622 -9011
rect 31676 -9045 31718 -9011
rect 32185 -9035 32227 -9001
rect 32257 -9035 32299 -9001
rect 32329 -9035 32371 -9001
rect 32401 -9029 32444 -9001
rect 32747 -9025 32789 -8991
rect 32792 -9025 32800 -8980
rect 32888 -8992 32894 -8809
rect 32922 -8995 32928 -8812
rect 32401 -9035 32443 -9029
rect 31838 -9088 31880 -9054
rect 31934 -9088 31976 -9054
rect 32030 -9088 32072 -9054
rect 32934 -9076 32942 -8809
rect 33271 -8812 33272 -8742
rect 33305 -8819 33306 -8740
rect 33788 -8741 33801 -8673
rect 33829 -8707 33835 -8639
rect 33874 -8671 33880 -8603
rect 33908 -8637 33914 -8571
rect 33918 -8621 33960 -8587
rect 34119 -8666 34161 -8632
rect 33888 -8689 33896 -8681
rect 33899 -8723 33941 -8689
rect 34119 -8734 34161 -8700
rect 33788 -8753 33796 -8741
rect 34168 -8750 34174 -8616
rect 33563 -8819 33957 -8753
rect 34202 -8784 34208 -8590
rect 34242 -8606 34250 -8595
rect 34238 -8637 34250 -8606
rect 34564 -8624 34606 -8590
rect 32950 -8860 32992 -8826
rect 33299 -8830 33317 -8819
rect 33299 -8832 33306 -8830
rect 32950 -8928 32992 -8894
rect 33002 -8995 33008 -8860
rect 33233 -8874 33306 -8832
rect 33361 -8874 33957 -8819
rect 34097 -8853 34139 -8819
rect 34142 -8853 34150 -8808
rect 34238 -8820 34244 -8637
rect 34272 -8823 34278 -8640
rect 33233 -8877 33957 -8874
rect 33036 -8980 33042 -8892
rect 33153 -8942 33195 -8908
rect 33198 -8942 33206 -8900
rect 33034 -8991 33042 -8980
rect 33036 -9025 33042 -8991
rect 33045 -9025 33087 -8991
rect 33153 -9042 33195 -9008
rect 33198 -9042 33206 -8997
rect 33046 -9078 33088 -9044
rect 33118 -9078 33160 -9044
rect 33190 -9078 33232 -9044
rect 32192 -9131 32234 -9097
rect 32288 -9131 32330 -9097
rect 32384 -9131 32426 -9097
rect 32480 -9131 32522 -9097
rect 32576 -9131 32618 -9097
rect 33233 -9114 33385 -8877
rect 33563 -8899 33957 -8877
rect 33487 -8925 33957 -8899
rect 34284 -8904 34292 -8637
rect 34621 -8640 34622 -8570
rect 34300 -8688 34342 -8654
rect 34655 -8674 34656 -8568
rect 34849 -8577 34891 -8543
rect 34894 -8577 34902 -8532
rect 34994 -8543 35002 -8532
rect 35203 -8537 35245 -8503
rect 35248 -8537 35256 -8492
rect 35348 -8503 35356 -8492
rect 35593 -8496 35635 -8462
rect 35638 -8496 35646 -8451
rect 35359 -8537 35401 -8503
rect 35005 -8577 35047 -8543
rect 34300 -8756 34342 -8722
rect 34352 -8823 34358 -8688
rect 34914 -8691 34956 -8657
rect 34966 -8718 34972 -8641
rect 34386 -8808 34392 -8720
rect 34503 -8770 34545 -8736
rect 34548 -8770 34556 -8728
rect 34648 -8740 34656 -8729
rect 34659 -8774 34701 -8740
rect 35000 -8752 35006 -8607
rect 35203 -8620 35245 -8586
rect 35248 -8620 35256 -8575
rect 35348 -8586 35356 -8575
rect 35593 -8580 35635 -8546
rect 35638 -8580 35646 -8535
rect 35359 -8620 35401 -8586
rect 35268 -8734 35310 -8700
rect 35320 -8761 35326 -8684
rect 34384 -8819 34392 -8808
rect 34853 -8813 34895 -8779
rect 34898 -8813 34906 -8771
rect 34998 -8779 35006 -8771
rect 35009 -8813 35051 -8779
rect 35354 -8795 35360 -8650
rect 35593 -8663 35635 -8629
rect 35638 -8663 35646 -8618
rect 35715 -8679 35721 -8413
rect 35749 -8413 35791 -8379
rect 35794 -8413 35802 -8371
rect 35738 -8462 35746 -8451
rect 35749 -8462 35755 -8413
rect 35749 -8496 35791 -8462
rect 35794 -8496 35802 -8451
rect 35738 -8546 35746 -8535
rect 35749 -8546 35755 -8496
rect 35749 -8580 35791 -8546
rect 35794 -8580 35802 -8535
rect 35738 -8629 35746 -8618
rect 35749 -8629 35755 -8580
rect 35749 -8663 35791 -8629
rect 35794 -8663 35802 -8618
rect 35738 -8697 35746 -8671
rect 35749 -8713 35755 -8663
rect 35658 -8777 35700 -8743
rect 35715 -8804 35716 -8727
rect 35749 -8809 35750 -8713
rect 34386 -8853 34392 -8819
rect 34395 -8853 34437 -8819
rect 34503 -8870 34545 -8836
rect 34548 -8870 34556 -8825
rect 34648 -8832 34656 -8821
rect 34659 -8866 34701 -8832
rect 35207 -8856 35249 -8822
rect 35252 -8856 35260 -8814
rect 35352 -8822 35360 -8814
rect 35363 -8856 35405 -8822
rect 35780 -8845 35788 -8697
rect 35803 -8713 35807 -8363
rect 35837 -8679 35841 -8363
rect 35894 -8379 35902 -8371
rect 35843 -8413 35885 -8379
rect 35905 -8413 35957 -8379
rect 36615 -8422 36621 -8406
rect 36638 -8422 36646 -8414
rect 36649 -8422 36655 -8406
rect 36945 -8408 36987 -8374
rect 36990 -8408 36998 -8363
rect 35894 -8462 35902 -8451
rect 36075 -8456 36117 -8422
rect 36147 -8456 36189 -8422
rect 36219 -8456 36261 -8422
rect 36363 -8456 36405 -8422
rect 36435 -8456 36549 -8422
rect 36579 -8456 36621 -8422
rect 35905 -8496 35947 -8462
rect 35894 -8546 35902 -8535
rect 36472 -8539 36514 -8505
rect 35905 -8580 35947 -8546
rect 35894 -8629 35902 -8618
rect 35905 -8663 35947 -8629
rect 36137 -8689 36179 -8655
rect 36182 -8689 36190 -8644
rect 36259 -8706 36265 -8588
rect 36282 -8655 36290 -8644
rect 36293 -8655 36299 -8622
rect 36329 -8655 36335 -8622
rect 36293 -8689 36335 -8655
rect 36338 -8689 36346 -8644
rect 36293 -8740 36299 -8689
rect 36329 -8740 36335 -8689
rect 36363 -8706 36369 -8589
rect 36460 -8630 36461 -8589
rect 36472 -8623 36514 -8589
rect 36472 -8706 36514 -8672
rect 36615 -8706 36621 -8456
rect 36649 -8456 36691 -8422
rect 36638 -8505 36646 -8494
rect 36649 -8505 36655 -8456
rect 36945 -8491 36987 -8457
rect 36990 -8491 36998 -8446
rect 36649 -8539 36691 -8505
rect 36638 -8589 36646 -8578
rect 36649 -8589 36655 -8539
rect 36799 -8565 36907 -8499
rect 37067 -8507 37073 -8241
rect 37101 -8241 37143 -8207
rect 37146 -8241 37154 -8199
rect 37090 -8290 37098 -8279
rect 37101 -8290 37107 -8241
rect 37101 -8324 37143 -8290
rect 37146 -8324 37154 -8279
rect 37090 -8374 37098 -8363
rect 37101 -8374 37107 -8324
rect 37101 -8408 37143 -8374
rect 37146 -8408 37154 -8363
rect 37090 -8457 37098 -8446
rect 37101 -8457 37107 -8408
rect 37101 -8491 37143 -8457
rect 37146 -8491 37154 -8446
rect 37090 -8525 37098 -8499
rect 37101 -8541 37107 -8491
rect 36649 -8623 36691 -8589
rect 37010 -8605 37052 -8571
rect 36638 -8672 36646 -8661
rect 36649 -8672 36655 -8623
rect 37067 -8632 37068 -8555
rect 37101 -8637 37102 -8541
rect 36649 -8706 36691 -8672
rect 37132 -8673 37140 -8525
rect 37155 -8541 37159 -8191
rect 37189 -8507 37193 -8191
rect 37246 -8207 37254 -8199
rect 37195 -8241 37237 -8207
rect 37257 -8241 37309 -8207
rect 38172 -8231 38214 -8197
rect 38268 -8231 38310 -8197
rect 38364 -8231 38406 -8197
rect 40334 -8207 40342 -8199
rect 40411 -8207 40417 -8191
rect 40434 -8207 40442 -8199
rect 40445 -8207 40451 -8191
rect 37965 -8250 37971 -8234
rect 37988 -8250 37996 -8242
rect 37999 -8250 38005 -8234
rect 37246 -8290 37254 -8279
rect 37425 -8284 37467 -8250
rect 37497 -8284 37539 -8250
rect 37569 -8284 37611 -8250
rect 37713 -8284 37755 -8250
rect 37785 -8284 37899 -8250
rect 37929 -8284 37971 -8250
rect 37257 -8324 37299 -8290
rect 37246 -8374 37254 -8363
rect 37822 -8367 37864 -8333
rect 37257 -8408 37299 -8374
rect 37246 -8457 37254 -8446
rect 37257 -8491 37299 -8457
rect 37487 -8517 37529 -8483
rect 37532 -8517 37540 -8472
rect 37609 -8534 37615 -8416
rect 37632 -8483 37640 -8472
rect 37643 -8483 37649 -8450
rect 37679 -8483 37685 -8450
rect 37643 -8517 37685 -8483
rect 37688 -8517 37696 -8472
rect 37643 -8568 37649 -8517
rect 37679 -8568 37685 -8517
rect 37713 -8534 37719 -8417
rect 37810 -8458 37811 -8417
rect 37822 -8451 37864 -8417
rect 37822 -8534 37864 -8500
rect 37965 -8534 37971 -8284
rect 37999 -8284 38041 -8250
rect 38526 -8274 38568 -8240
rect 38622 -8274 38664 -8240
rect 38718 -8274 38760 -8240
rect 40225 -8241 40267 -8207
rect 40289 -8241 40342 -8207
rect 40369 -8241 40417 -8207
rect 37988 -8333 37996 -8322
rect 37999 -8333 38005 -8284
rect 38238 -8293 38246 -8285
rect 38338 -8293 38346 -8285
rect 38165 -8327 38235 -8293
rect 38237 -8327 38279 -8293
rect 38349 -8327 38391 -8293
rect 38880 -8317 38922 -8283
rect 38976 -8317 39018 -8283
rect 39072 -8317 39114 -8283
rect 39168 -8317 39210 -8283
rect 39264 -8317 39306 -8283
rect 40289 -8324 40331 -8290
rect 40334 -8324 40342 -8279
rect 37999 -8367 38041 -8333
rect 38592 -8336 38600 -8328
rect 38692 -8336 38700 -8328
rect 37988 -8417 37996 -8406
rect 37999 -8417 38005 -8367
rect 38193 -8410 38235 -8376
rect 38238 -8410 38246 -8365
rect 38338 -8376 38346 -8365
rect 38519 -8370 38589 -8336
rect 38591 -8370 38633 -8336
rect 38703 -8370 38745 -8336
rect 39428 -8360 39470 -8326
rect 39524 -8360 39566 -8326
rect 39620 -8360 39662 -8326
rect 39716 -8360 39758 -8326
rect 39812 -8360 39854 -8326
rect 39908 -8360 39950 -8326
rect 40004 -8360 40046 -8326
rect 38349 -8410 38391 -8376
rect 38982 -8379 38990 -8371
rect 39059 -8379 39065 -8363
rect 39082 -8379 39090 -8371
rect 39093 -8379 39099 -8363
rect 37999 -8451 38041 -8417
rect 37988 -8500 37996 -8489
rect 37999 -8500 38005 -8451
rect 38193 -8494 38235 -8460
rect 38238 -8494 38246 -8449
rect 38338 -8460 38346 -8449
rect 38547 -8453 38589 -8419
rect 38592 -8453 38600 -8408
rect 38692 -8419 38700 -8408
rect 38873 -8413 38915 -8379
rect 38937 -8413 38990 -8379
rect 39017 -8413 39065 -8379
rect 38703 -8453 38745 -8419
rect 38349 -8494 38391 -8460
rect 37999 -8534 38041 -8500
rect 37999 -8568 38005 -8534
rect 36649 -8740 36655 -8706
rect 36945 -8723 36987 -8689
rect 36990 -8723 36998 -8681
rect 34396 -8906 34438 -8872
rect 34468 -8906 34510 -8872
rect 34540 -8906 34582 -8872
rect 34853 -8913 34895 -8879
rect 34898 -8913 34906 -8868
rect 34998 -8879 35006 -8868
rect 35009 -8913 35051 -8879
rect 35593 -8895 35635 -8861
rect 35638 -8895 35646 -8853
rect 33487 -8959 33970 -8925
rect 34821 -8949 34863 -8915
rect 34893 -8949 34935 -8915
rect 35207 -8956 35249 -8922
rect 35252 -8956 35260 -8911
rect 35352 -8922 35360 -8911
rect 35780 -8913 35793 -8845
rect 35821 -8879 35827 -8811
rect 35866 -8843 35872 -8775
rect 35900 -8809 35906 -8743
rect 35910 -8793 35952 -8759
rect 36113 -8838 36155 -8804
rect 35880 -8861 35888 -8853
rect 35891 -8895 35933 -8861
rect 36113 -8906 36155 -8872
rect 35363 -8956 35405 -8922
rect 33487 -8985 33957 -8959
rect 33491 -8993 33699 -8985
rect 33507 -9003 33683 -8993
rect 33233 -9140 33415 -9114
rect 32740 -9174 32782 -9140
rect 32836 -9174 32878 -9140
rect 32932 -9174 32974 -9140
rect 33028 -9174 33070 -9140
rect 33124 -9174 33166 -9140
rect 33220 -9174 33415 -9140
rect 33233 -9200 33415 -9174
rect 33433 -9174 33541 -9050
rect 33692 -9062 33699 -9051
rect 33311 -9870 33353 -9200
rect 33433 -9228 33443 -9174
rect 33118 -9936 33270 -9924
rect 32786 -9970 33270 -9936
rect 33118 -9971 33270 -9970
rect 33299 -9971 33353 -9870
rect 33445 -9971 33487 -9174
rect 33491 -9971 33498 -9174
rect 33703 -9971 33745 -9062
rect 33837 -9971 33879 -8985
rect 34090 -9002 34132 -8968
rect 34186 -9002 34228 -8968
rect 34282 -9002 34324 -8968
rect 34378 -9002 34420 -8968
rect 34474 -9002 34516 -8968
rect 34570 -9002 34612 -8968
rect 34666 -9002 34708 -8968
rect 35175 -8992 35217 -8958
rect 35247 -8992 35289 -8958
rect 35593 -8995 35635 -8961
rect 35638 -8995 35646 -8950
rect 35780 -9001 35788 -8913
rect 36162 -8922 36168 -8788
rect 35880 -8961 35888 -8950
rect 36196 -8956 36202 -8762
rect 36236 -8778 36244 -8767
rect 36232 -8809 36244 -8778
rect 36558 -8796 36600 -8762
rect 35891 -8995 35933 -8961
rect 34828 -9045 34870 -9011
rect 34924 -9045 34966 -9011
rect 35020 -9045 35062 -9011
rect 35529 -9035 35571 -9001
rect 35601 -9035 35643 -9001
rect 35673 -9035 35715 -9001
rect 35745 -9029 35788 -9001
rect 36091 -9025 36133 -8991
rect 36136 -9025 36144 -8980
rect 36232 -8992 36238 -8809
rect 36266 -8995 36272 -8812
rect 35745 -9035 35787 -9029
rect 35182 -9088 35224 -9054
rect 35278 -9088 35320 -9054
rect 35374 -9088 35416 -9054
rect 36278 -9076 36286 -8809
rect 36615 -8812 36616 -8742
rect 36649 -8819 36650 -8740
rect 37132 -8741 37145 -8673
rect 37173 -8707 37179 -8639
rect 37218 -8671 37224 -8603
rect 37252 -8637 37258 -8571
rect 37262 -8621 37304 -8587
rect 37463 -8666 37505 -8632
rect 37232 -8689 37240 -8681
rect 37243 -8723 37285 -8689
rect 37463 -8734 37505 -8700
rect 37132 -8753 37140 -8741
rect 37512 -8750 37518 -8616
rect 36907 -8819 37301 -8753
rect 37546 -8784 37552 -8590
rect 37586 -8606 37594 -8595
rect 37582 -8637 37594 -8606
rect 37908 -8624 37950 -8590
rect 36294 -8860 36336 -8826
rect 36643 -8830 36661 -8819
rect 36643 -8832 36650 -8830
rect 36294 -8928 36336 -8894
rect 36346 -8995 36352 -8860
rect 36577 -8874 36650 -8832
rect 36705 -8874 37301 -8819
rect 37441 -8853 37483 -8819
rect 37486 -8853 37494 -8808
rect 37582 -8820 37588 -8637
rect 37616 -8823 37622 -8640
rect 36577 -8877 37301 -8874
rect 36380 -8980 36386 -8892
rect 36497 -8942 36539 -8908
rect 36542 -8942 36550 -8900
rect 36378 -8991 36386 -8980
rect 36380 -9025 36386 -8991
rect 36389 -9025 36431 -8991
rect 36497 -9042 36539 -9008
rect 36542 -9042 36550 -8997
rect 36390 -9078 36432 -9044
rect 36462 -9078 36504 -9044
rect 36534 -9078 36576 -9044
rect 35536 -9131 35578 -9097
rect 35632 -9131 35674 -9097
rect 35728 -9131 35770 -9097
rect 35824 -9131 35866 -9097
rect 35920 -9131 35962 -9097
rect 36577 -9114 36729 -8877
rect 36907 -8899 37301 -8877
rect 36831 -8925 37301 -8899
rect 37628 -8904 37636 -8637
rect 37965 -8640 37966 -8570
rect 37644 -8688 37686 -8654
rect 37999 -8674 38000 -8568
rect 38193 -8577 38235 -8543
rect 38238 -8577 38246 -8532
rect 38338 -8543 38346 -8532
rect 38547 -8537 38589 -8503
rect 38592 -8537 38600 -8492
rect 38692 -8503 38700 -8492
rect 38937 -8496 38979 -8462
rect 38982 -8496 38990 -8451
rect 38703 -8537 38745 -8503
rect 38349 -8577 38391 -8543
rect 37644 -8756 37686 -8722
rect 37696 -8823 37702 -8688
rect 38258 -8691 38300 -8657
rect 38310 -8718 38316 -8641
rect 37730 -8808 37736 -8720
rect 37847 -8770 37889 -8736
rect 37892 -8770 37900 -8728
rect 37992 -8740 38000 -8729
rect 38003 -8774 38045 -8740
rect 38344 -8752 38350 -8607
rect 38547 -8620 38589 -8586
rect 38592 -8620 38600 -8575
rect 38692 -8586 38700 -8575
rect 38937 -8580 38979 -8546
rect 38982 -8580 38990 -8535
rect 38703 -8620 38745 -8586
rect 38612 -8734 38654 -8700
rect 38664 -8761 38670 -8684
rect 37728 -8819 37736 -8808
rect 38197 -8813 38239 -8779
rect 38242 -8813 38250 -8771
rect 38342 -8779 38350 -8771
rect 38353 -8813 38395 -8779
rect 38698 -8795 38704 -8650
rect 38937 -8663 38979 -8629
rect 38982 -8663 38990 -8618
rect 39059 -8679 39065 -8413
rect 39093 -8413 39135 -8379
rect 39138 -8413 39146 -8371
rect 39082 -8462 39090 -8451
rect 39093 -8462 39099 -8413
rect 39093 -8496 39135 -8462
rect 39138 -8496 39146 -8451
rect 39082 -8546 39090 -8535
rect 39093 -8546 39099 -8496
rect 39093 -8580 39135 -8546
rect 39138 -8580 39146 -8535
rect 39082 -8629 39090 -8618
rect 39093 -8629 39099 -8580
rect 39093 -8663 39135 -8629
rect 39138 -8663 39146 -8618
rect 39082 -8697 39090 -8671
rect 39093 -8713 39099 -8663
rect 39002 -8777 39044 -8743
rect 39059 -8804 39060 -8727
rect 39093 -8809 39094 -8713
rect 37730 -8853 37736 -8819
rect 37739 -8853 37781 -8819
rect 37847 -8870 37889 -8836
rect 37892 -8870 37900 -8825
rect 37992 -8832 38000 -8821
rect 38003 -8866 38045 -8832
rect 38551 -8856 38593 -8822
rect 38596 -8856 38604 -8814
rect 38696 -8822 38704 -8814
rect 38707 -8856 38749 -8822
rect 39124 -8845 39132 -8697
rect 39147 -8713 39151 -8363
rect 39181 -8679 39185 -8363
rect 39238 -8379 39246 -8371
rect 39187 -8413 39229 -8379
rect 39249 -8413 39301 -8379
rect 39959 -8422 39965 -8406
rect 39982 -8422 39990 -8414
rect 39993 -8422 39999 -8406
rect 40289 -8408 40331 -8374
rect 40334 -8408 40342 -8363
rect 39238 -8462 39246 -8451
rect 39419 -8456 39461 -8422
rect 39491 -8456 39533 -8422
rect 39563 -8456 39605 -8422
rect 39707 -8456 39749 -8422
rect 39779 -8456 39893 -8422
rect 39923 -8456 39965 -8422
rect 39249 -8496 39291 -8462
rect 39238 -8546 39246 -8535
rect 39816 -8539 39858 -8505
rect 39249 -8580 39291 -8546
rect 39238 -8629 39246 -8618
rect 39249 -8663 39291 -8629
rect 39481 -8689 39523 -8655
rect 39526 -8689 39534 -8644
rect 39603 -8706 39609 -8588
rect 39626 -8655 39634 -8644
rect 39637 -8655 39643 -8622
rect 39673 -8655 39679 -8622
rect 39637 -8689 39679 -8655
rect 39682 -8689 39690 -8644
rect 39637 -8740 39643 -8689
rect 39673 -8740 39679 -8689
rect 39707 -8706 39713 -8589
rect 39804 -8630 39805 -8589
rect 39816 -8623 39858 -8589
rect 39816 -8706 39858 -8672
rect 39959 -8706 39965 -8456
rect 39993 -8456 40035 -8422
rect 39982 -8505 39990 -8494
rect 39993 -8505 39999 -8456
rect 40289 -8491 40331 -8457
rect 40334 -8491 40342 -8446
rect 39993 -8539 40035 -8505
rect 39982 -8589 39990 -8578
rect 39993 -8589 39999 -8539
rect 40143 -8565 40251 -8499
rect 40411 -8507 40417 -8241
rect 40445 -8241 40487 -8207
rect 40490 -8241 40498 -8199
rect 40434 -8290 40442 -8279
rect 40445 -8290 40451 -8241
rect 40445 -8324 40487 -8290
rect 40490 -8324 40498 -8279
rect 40434 -8374 40442 -8363
rect 40445 -8374 40451 -8324
rect 40445 -8408 40487 -8374
rect 40490 -8408 40498 -8363
rect 40434 -8457 40442 -8446
rect 40445 -8457 40451 -8408
rect 40445 -8491 40487 -8457
rect 40490 -8491 40498 -8446
rect 40434 -8525 40442 -8499
rect 40445 -8541 40451 -8491
rect 39993 -8623 40035 -8589
rect 40354 -8605 40396 -8571
rect 39982 -8672 39990 -8661
rect 39993 -8672 39999 -8623
rect 40411 -8632 40412 -8555
rect 40445 -8637 40446 -8541
rect 39993 -8706 40035 -8672
rect 40476 -8673 40484 -8525
rect 40499 -8541 40503 -8191
rect 40533 -8507 40537 -8191
rect 40590 -8207 40598 -8199
rect 40539 -8241 40581 -8207
rect 40601 -8241 40653 -8207
rect 41516 -8231 41558 -8197
rect 41612 -8231 41654 -8197
rect 41708 -8231 41750 -8197
rect 43678 -8207 43686 -8199
rect 43755 -8207 43761 -8191
rect 43778 -8207 43786 -8199
rect 43789 -8207 43795 -8191
rect 41309 -8250 41315 -8234
rect 41332 -8250 41340 -8242
rect 41343 -8250 41349 -8234
rect 40590 -8290 40598 -8279
rect 40769 -8284 40811 -8250
rect 40841 -8284 40883 -8250
rect 40913 -8284 40955 -8250
rect 41057 -8284 41099 -8250
rect 41129 -8284 41243 -8250
rect 41273 -8284 41315 -8250
rect 40601 -8324 40643 -8290
rect 40590 -8374 40598 -8363
rect 41166 -8367 41208 -8333
rect 40601 -8408 40643 -8374
rect 40590 -8457 40598 -8446
rect 40601 -8491 40643 -8457
rect 40831 -8517 40873 -8483
rect 40876 -8517 40884 -8472
rect 40953 -8534 40959 -8416
rect 40976 -8483 40984 -8472
rect 40987 -8483 40993 -8450
rect 41023 -8483 41029 -8450
rect 40987 -8517 41029 -8483
rect 41032 -8517 41040 -8472
rect 40987 -8568 40993 -8517
rect 41023 -8568 41029 -8517
rect 41057 -8534 41063 -8417
rect 41154 -8458 41155 -8417
rect 41166 -8451 41208 -8417
rect 41166 -8534 41208 -8500
rect 41309 -8534 41315 -8284
rect 41343 -8284 41385 -8250
rect 41870 -8274 41912 -8240
rect 41966 -8274 42008 -8240
rect 42062 -8274 42104 -8240
rect 43569 -8241 43611 -8207
rect 43633 -8241 43686 -8207
rect 43713 -8241 43761 -8207
rect 41332 -8333 41340 -8322
rect 41343 -8333 41349 -8284
rect 41582 -8293 41590 -8285
rect 41682 -8293 41690 -8285
rect 41509 -8327 41579 -8293
rect 41581 -8327 41623 -8293
rect 41693 -8327 41735 -8293
rect 42224 -8317 42266 -8283
rect 42320 -8317 42362 -8283
rect 42416 -8317 42458 -8283
rect 42512 -8317 42554 -8283
rect 42608 -8317 42650 -8283
rect 43633 -8324 43675 -8290
rect 43678 -8324 43686 -8279
rect 41343 -8367 41385 -8333
rect 41936 -8336 41944 -8328
rect 42036 -8336 42044 -8328
rect 41332 -8417 41340 -8406
rect 41343 -8417 41349 -8367
rect 41537 -8410 41579 -8376
rect 41582 -8410 41590 -8365
rect 41682 -8376 41690 -8365
rect 41863 -8370 41933 -8336
rect 41935 -8370 41977 -8336
rect 42047 -8370 42089 -8336
rect 42772 -8360 42814 -8326
rect 42868 -8360 42910 -8326
rect 42964 -8360 43006 -8326
rect 43060 -8360 43102 -8326
rect 43156 -8360 43198 -8326
rect 43252 -8360 43294 -8326
rect 43348 -8360 43390 -8326
rect 41693 -8410 41735 -8376
rect 42326 -8379 42334 -8371
rect 42403 -8379 42409 -8363
rect 42426 -8379 42434 -8371
rect 42437 -8379 42443 -8363
rect 41343 -8451 41385 -8417
rect 41332 -8500 41340 -8489
rect 41343 -8500 41349 -8451
rect 41537 -8494 41579 -8460
rect 41582 -8494 41590 -8449
rect 41682 -8460 41690 -8449
rect 41891 -8453 41933 -8419
rect 41936 -8453 41944 -8408
rect 42036 -8419 42044 -8408
rect 42217 -8413 42259 -8379
rect 42281 -8413 42334 -8379
rect 42361 -8413 42409 -8379
rect 42047 -8453 42089 -8419
rect 41693 -8494 41735 -8460
rect 41343 -8534 41385 -8500
rect 41343 -8568 41349 -8534
rect 39993 -8740 39999 -8706
rect 40289 -8723 40331 -8689
rect 40334 -8723 40342 -8681
rect 37740 -8906 37782 -8872
rect 37812 -8906 37854 -8872
rect 37884 -8906 37926 -8872
rect 38197 -8913 38239 -8879
rect 38242 -8913 38250 -8868
rect 38342 -8879 38350 -8868
rect 38353 -8913 38395 -8879
rect 38937 -8895 38979 -8861
rect 38982 -8895 38990 -8853
rect 36831 -8959 37314 -8925
rect 38165 -8949 38207 -8915
rect 38237 -8949 38279 -8915
rect 38551 -8956 38593 -8922
rect 38596 -8956 38604 -8911
rect 38696 -8922 38704 -8911
rect 39124 -8913 39137 -8845
rect 39165 -8879 39171 -8811
rect 39210 -8843 39216 -8775
rect 39244 -8809 39250 -8743
rect 39254 -8793 39296 -8759
rect 39457 -8838 39499 -8804
rect 39224 -8861 39232 -8853
rect 39235 -8895 39277 -8861
rect 39457 -8906 39499 -8872
rect 38707 -8956 38749 -8922
rect 36831 -8985 37301 -8959
rect 36835 -8993 37043 -8985
rect 36851 -9003 37027 -8993
rect 36577 -9140 36759 -9114
rect 36084 -9174 36126 -9140
rect 36180 -9174 36222 -9140
rect 36276 -9174 36318 -9140
rect 36372 -9174 36414 -9140
rect 36468 -9174 36510 -9140
rect 36564 -9174 36759 -9140
rect 36577 -9200 36759 -9174
rect 36777 -9174 36885 -9050
rect 37036 -9062 37043 -9051
rect 36655 -9870 36697 -9200
rect 36777 -9228 36787 -9174
rect 36462 -9936 36614 -9924
rect 36130 -9970 36614 -9936
rect 36462 -9971 36614 -9970
rect 36643 -9971 36697 -9870
rect 36789 -9971 36831 -9174
rect 36835 -9971 36842 -9174
rect 37047 -9971 37089 -9062
rect 37181 -9971 37223 -8985
rect 37434 -9002 37476 -8968
rect 37530 -9002 37572 -8968
rect 37626 -9002 37668 -8968
rect 37722 -9002 37764 -8968
rect 37818 -9002 37860 -8968
rect 37914 -9002 37956 -8968
rect 38010 -9002 38052 -8968
rect 38519 -8992 38561 -8958
rect 38591 -8992 38633 -8958
rect 38937 -8995 38979 -8961
rect 38982 -8995 38990 -8950
rect 39124 -9001 39132 -8913
rect 39506 -8922 39512 -8788
rect 39224 -8961 39232 -8950
rect 39540 -8956 39546 -8762
rect 39580 -8778 39588 -8767
rect 39576 -8809 39588 -8778
rect 39902 -8796 39944 -8762
rect 39235 -8995 39277 -8961
rect 38172 -9045 38214 -9011
rect 38268 -9045 38310 -9011
rect 38364 -9045 38406 -9011
rect 38873 -9035 38915 -9001
rect 38945 -9035 38987 -9001
rect 39017 -9035 39059 -9001
rect 39089 -9029 39132 -9001
rect 39435 -9025 39477 -8991
rect 39480 -9025 39488 -8980
rect 39576 -8992 39582 -8809
rect 39610 -8995 39616 -8812
rect 39089 -9035 39131 -9029
rect 38526 -9088 38568 -9054
rect 38622 -9088 38664 -9054
rect 38718 -9088 38760 -9054
rect 39622 -9076 39630 -8809
rect 39959 -8812 39960 -8742
rect 39993 -8819 39994 -8740
rect 40476 -8741 40489 -8673
rect 40517 -8707 40523 -8639
rect 40562 -8671 40568 -8603
rect 40596 -8637 40602 -8571
rect 40606 -8621 40648 -8587
rect 40807 -8666 40849 -8632
rect 40576 -8689 40584 -8681
rect 40587 -8723 40629 -8689
rect 40807 -8734 40849 -8700
rect 40476 -8753 40484 -8741
rect 40856 -8750 40862 -8616
rect 40251 -8819 40645 -8753
rect 40890 -8784 40896 -8590
rect 40930 -8606 40938 -8595
rect 40926 -8637 40938 -8606
rect 41252 -8624 41294 -8590
rect 39638 -8860 39680 -8826
rect 39987 -8830 40005 -8819
rect 39987 -8832 39994 -8830
rect 39638 -8928 39680 -8894
rect 39690 -8995 39696 -8860
rect 39921 -8874 39994 -8832
rect 40049 -8874 40645 -8819
rect 40785 -8853 40827 -8819
rect 40830 -8853 40838 -8808
rect 40926 -8820 40932 -8637
rect 40960 -8823 40966 -8640
rect 39921 -8877 40645 -8874
rect 39724 -8980 39730 -8892
rect 39841 -8942 39883 -8908
rect 39886 -8942 39894 -8900
rect 39722 -8991 39730 -8980
rect 39724 -9025 39730 -8991
rect 39733 -9025 39775 -8991
rect 39841 -9042 39883 -9008
rect 39886 -9042 39894 -8997
rect 39734 -9078 39776 -9044
rect 39806 -9078 39848 -9044
rect 39878 -9078 39920 -9044
rect 38880 -9131 38922 -9097
rect 38976 -9131 39018 -9097
rect 39072 -9131 39114 -9097
rect 39168 -9131 39210 -9097
rect 39264 -9131 39306 -9097
rect 39921 -9114 40073 -8877
rect 40251 -8899 40645 -8877
rect 40175 -8925 40645 -8899
rect 40972 -8904 40980 -8637
rect 41309 -8640 41310 -8570
rect 40988 -8688 41030 -8654
rect 41343 -8674 41344 -8568
rect 41537 -8577 41579 -8543
rect 41582 -8577 41590 -8532
rect 41682 -8543 41690 -8532
rect 41891 -8537 41933 -8503
rect 41936 -8537 41944 -8492
rect 42036 -8503 42044 -8492
rect 42281 -8496 42323 -8462
rect 42326 -8496 42334 -8451
rect 42047 -8537 42089 -8503
rect 41693 -8577 41735 -8543
rect 40988 -8756 41030 -8722
rect 41040 -8823 41046 -8688
rect 41602 -8691 41644 -8657
rect 41654 -8718 41660 -8641
rect 41074 -8808 41080 -8720
rect 41191 -8770 41233 -8736
rect 41236 -8770 41244 -8728
rect 41336 -8740 41344 -8729
rect 41347 -8774 41389 -8740
rect 41688 -8752 41694 -8607
rect 41891 -8620 41933 -8586
rect 41936 -8620 41944 -8575
rect 42036 -8586 42044 -8575
rect 42281 -8580 42323 -8546
rect 42326 -8580 42334 -8535
rect 42047 -8620 42089 -8586
rect 41956 -8734 41998 -8700
rect 42008 -8761 42014 -8684
rect 41072 -8819 41080 -8808
rect 41541 -8813 41583 -8779
rect 41586 -8813 41594 -8771
rect 41686 -8779 41694 -8771
rect 41697 -8813 41739 -8779
rect 42042 -8795 42048 -8650
rect 42281 -8663 42323 -8629
rect 42326 -8663 42334 -8618
rect 42403 -8679 42409 -8413
rect 42437 -8413 42479 -8379
rect 42482 -8413 42490 -8371
rect 42426 -8462 42434 -8451
rect 42437 -8462 42443 -8413
rect 42437 -8496 42479 -8462
rect 42482 -8496 42490 -8451
rect 42426 -8546 42434 -8535
rect 42437 -8546 42443 -8496
rect 42437 -8580 42479 -8546
rect 42482 -8580 42490 -8535
rect 42426 -8629 42434 -8618
rect 42437 -8629 42443 -8580
rect 42437 -8663 42479 -8629
rect 42482 -8663 42490 -8618
rect 42426 -8697 42434 -8671
rect 42437 -8713 42443 -8663
rect 42346 -8777 42388 -8743
rect 42403 -8804 42404 -8727
rect 42437 -8809 42438 -8713
rect 41074 -8853 41080 -8819
rect 41083 -8853 41125 -8819
rect 41191 -8870 41233 -8836
rect 41236 -8870 41244 -8825
rect 41336 -8832 41344 -8821
rect 41347 -8866 41389 -8832
rect 41895 -8856 41937 -8822
rect 41940 -8856 41948 -8814
rect 42040 -8822 42048 -8814
rect 42051 -8856 42093 -8822
rect 42468 -8845 42476 -8697
rect 42491 -8713 42495 -8363
rect 42525 -8679 42529 -8363
rect 42582 -8379 42590 -8371
rect 42531 -8413 42573 -8379
rect 42593 -8413 42645 -8379
rect 43303 -8422 43309 -8406
rect 43326 -8422 43334 -8414
rect 43337 -8422 43343 -8406
rect 43633 -8408 43675 -8374
rect 43678 -8408 43686 -8363
rect 42582 -8462 42590 -8451
rect 42763 -8456 42805 -8422
rect 42835 -8456 42877 -8422
rect 42907 -8456 42949 -8422
rect 43051 -8456 43093 -8422
rect 43123 -8456 43237 -8422
rect 43267 -8456 43309 -8422
rect 42593 -8496 42635 -8462
rect 42582 -8546 42590 -8535
rect 43160 -8539 43202 -8505
rect 42593 -8580 42635 -8546
rect 42582 -8629 42590 -8618
rect 42593 -8663 42635 -8629
rect 42825 -8689 42867 -8655
rect 42870 -8689 42878 -8644
rect 42947 -8706 42953 -8588
rect 42970 -8655 42978 -8644
rect 42981 -8655 42987 -8622
rect 43017 -8655 43023 -8622
rect 42981 -8689 43023 -8655
rect 43026 -8689 43034 -8644
rect 42981 -8740 42987 -8689
rect 43017 -8740 43023 -8689
rect 43051 -8706 43057 -8589
rect 43148 -8630 43149 -8589
rect 43160 -8623 43202 -8589
rect 43160 -8706 43202 -8672
rect 43303 -8706 43309 -8456
rect 43337 -8456 43379 -8422
rect 43326 -8505 43334 -8494
rect 43337 -8505 43343 -8456
rect 43633 -8491 43675 -8457
rect 43678 -8491 43686 -8446
rect 43337 -8539 43379 -8505
rect 43326 -8589 43334 -8578
rect 43337 -8589 43343 -8539
rect 43487 -8565 43595 -8499
rect 43755 -8507 43761 -8241
rect 43789 -8241 43831 -8207
rect 43834 -8241 43842 -8199
rect 43778 -8290 43786 -8279
rect 43789 -8290 43795 -8241
rect 43789 -8324 43831 -8290
rect 43834 -8324 43842 -8279
rect 43778 -8374 43786 -8363
rect 43789 -8374 43795 -8324
rect 43789 -8408 43831 -8374
rect 43834 -8408 43842 -8363
rect 43778 -8457 43786 -8446
rect 43789 -8457 43795 -8408
rect 43789 -8491 43831 -8457
rect 43834 -8491 43842 -8446
rect 43778 -8525 43786 -8499
rect 43789 -8541 43795 -8491
rect 43337 -8623 43379 -8589
rect 43698 -8605 43740 -8571
rect 43326 -8672 43334 -8661
rect 43337 -8672 43343 -8623
rect 43755 -8632 43756 -8555
rect 43789 -8637 43790 -8541
rect 43337 -8706 43379 -8672
rect 43820 -8673 43828 -8525
rect 43843 -8541 43847 -8191
rect 43877 -8507 43881 -8191
rect 43934 -8207 43942 -8199
rect 43883 -8241 43925 -8207
rect 43945 -8241 43997 -8207
rect 44860 -8231 44902 -8197
rect 44956 -8231 44998 -8197
rect 45052 -8231 45094 -8197
rect 47022 -8207 47030 -8199
rect 47099 -8207 47105 -8191
rect 47122 -8207 47130 -8199
rect 47133 -8207 47139 -8191
rect 44653 -8250 44659 -8234
rect 44676 -8250 44684 -8242
rect 44687 -8250 44693 -8234
rect 43934 -8290 43942 -8279
rect 44113 -8284 44155 -8250
rect 44185 -8284 44227 -8250
rect 44257 -8284 44299 -8250
rect 44401 -8284 44443 -8250
rect 44473 -8284 44587 -8250
rect 44617 -8284 44659 -8250
rect 43945 -8324 43987 -8290
rect 43934 -8374 43942 -8363
rect 44510 -8367 44552 -8333
rect 43945 -8408 43987 -8374
rect 43934 -8457 43942 -8446
rect 43945 -8491 43987 -8457
rect 44175 -8517 44217 -8483
rect 44220 -8517 44228 -8472
rect 44297 -8534 44303 -8416
rect 44320 -8483 44328 -8472
rect 44331 -8483 44337 -8450
rect 44367 -8483 44373 -8450
rect 44331 -8517 44373 -8483
rect 44376 -8517 44384 -8472
rect 44331 -8568 44337 -8517
rect 44367 -8568 44373 -8517
rect 44401 -8534 44407 -8417
rect 44498 -8458 44499 -8417
rect 44510 -8451 44552 -8417
rect 44510 -8534 44552 -8500
rect 44653 -8534 44659 -8284
rect 44687 -8284 44729 -8250
rect 45214 -8274 45256 -8240
rect 45310 -8274 45352 -8240
rect 45406 -8274 45448 -8240
rect 46913 -8241 46955 -8207
rect 46977 -8241 47030 -8207
rect 47057 -8241 47105 -8207
rect 44676 -8333 44684 -8322
rect 44687 -8333 44693 -8284
rect 44926 -8293 44934 -8285
rect 45026 -8293 45034 -8285
rect 44853 -8327 44923 -8293
rect 44925 -8327 44967 -8293
rect 45037 -8327 45079 -8293
rect 45568 -8317 45610 -8283
rect 45664 -8317 45706 -8283
rect 45760 -8317 45802 -8283
rect 45856 -8317 45898 -8283
rect 45952 -8317 45994 -8283
rect 46977 -8324 47019 -8290
rect 47022 -8324 47030 -8279
rect 44687 -8367 44729 -8333
rect 45280 -8336 45288 -8328
rect 45380 -8336 45388 -8328
rect 44676 -8417 44684 -8406
rect 44687 -8417 44693 -8367
rect 44881 -8410 44923 -8376
rect 44926 -8410 44934 -8365
rect 45026 -8376 45034 -8365
rect 45207 -8370 45277 -8336
rect 45279 -8370 45321 -8336
rect 45391 -8370 45433 -8336
rect 46116 -8360 46158 -8326
rect 46212 -8360 46254 -8326
rect 46308 -8360 46350 -8326
rect 46404 -8360 46446 -8326
rect 46500 -8360 46542 -8326
rect 46596 -8360 46638 -8326
rect 46692 -8360 46734 -8326
rect 45037 -8410 45079 -8376
rect 45670 -8379 45678 -8371
rect 45747 -8379 45753 -8363
rect 45770 -8379 45778 -8371
rect 45781 -8379 45787 -8363
rect 44687 -8451 44729 -8417
rect 44676 -8500 44684 -8489
rect 44687 -8500 44693 -8451
rect 44881 -8494 44923 -8460
rect 44926 -8494 44934 -8449
rect 45026 -8460 45034 -8449
rect 45235 -8453 45277 -8419
rect 45280 -8453 45288 -8408
rect 45380 -8419 45388 -8408
rect 45561 -8413 45603 -8379
rect 45625 -8413 45678 -8379
rect 45705 -8413 45753 -8379
rect 45391 -8453 45433 -8419
rect 45037 -8494 45079 -8460
rect 44687 -8534 44729 -8500
rect 44687 -8568 44693 -8534
rect 43337 -8740 43343 -8706
rect 43633 -8723 43675 -8689
rect 43678 -8723 43686 -8681
rect 41084 -8906 41126 -8872
rect 41156 -8906 41198 -8872
rect 41228 -8906 41270 -8872
rect 41541 -8913 41583 -8879
rect 41586 -8913 41594 -8868
rect 41686 -8879 41694 -8868
rect 41697 -8913 41739 -8879
rect 42281 -8895 42323 -8861
rect 42326 -8895 42334 -8853
rect 40175 -8959 40658 -8925
rect 41509 -8949 41551 -8915
rect 41581 -8949 41623 -8915
rect 41895 -8956 41937 -8922
rect 41940 -8956 41948 -8911
rect 42040 -8922 42048 -8911
rect 42468 -8913 42481 -8845
rect 42509 -8879 42515 -8811
rect 42554 -8843 42560 -8775
rect 42588 -8809 42594 -8743
rect 42598 -8793 42640 -8759
rect 42801 -8838 42843 -8804
rect 42568 -8861 42576 -8853
rect 42579 -8895 42621 -8861
rect 42801 -8906 42843 -8872
rect 42051 -8956 42093 -8922
rect 40175 -8985 40645 -8959
rect 40179 -8993 40387 -8985
rect 40195 -9003 40371 -8993
rect 39921 -9140 40103 -9114
rect 39428 -9174 39470 -9140
rect 39524 -9174 39566 -9140
rect 39620 -9174 39662 -9140
rect 39716 -9174 39758 -9140
rect 39812 -9174 39854 -9140
rect 39908 -9174 40103 -9140
rect 39921 -9200 40103 -9174
rect 40121 -9174 40229 -9050
rect 40380 -9062 40387 -9051
rect 39999 -9870 40041 -9200
rect 40121 -9228 40131 -9174
rect 39806 -9936 39958 -9924
rect 39474 -9970 39958 -9936
rect 39806 -9971 39958 -9970
rect 39987 -9971 40041 -9870
rect 40133 -9971 40175 -9174
rect 40179 -9971 40186 -9174
rect 40391 -9971 40433 -9062
rect 40525 -9971 40567 -8985
rect 40778 -9002 40820 -8968
rect 40874 -9002 40916 -8968
rect 40970 -9002 41012 -8968
rect 41066 -9002 41108 -8968
rect 41162 -9002 41204 -8968
rect 41258 -9002 41300 -8968
rect 41354 -9002 41396 -8968
rect 41863 -8992 41905 -8958
rect 41935 -8992 41977 -8958
rect 42281 -8995 42323 -8961
rect 42326 -8995 42334 -8950
rect 42468 -9001 42476 -8913
rect 42850 -8922 42856 -8788
rect 42568 -8961 42576 -8950
rect 42884 -8956 42890 -8762
rect 42924 -8778 42932 -8767
rect 42920 -8809 42932 -8778
rect 43246 -8796 43288 -8762
rect 42579 -8995 42621 -8961
rect 41516 -9045 41558 -9011
rect 41612 -9045 41654 -9011
rect 41708 -9045 41750 -9011
rect 42217 -9035 42259 -9001
rect 42289 -9035 42331 -9001
rect 42361 -9035 42403 -9001
rect 42433 -9029 42476 -9001
rect 42779 -9025 42821 -8991
rect 42824 -9025 42832 -8980
rect 42920 -8992 42926 -8809
rect 42954 -8995 42960 -8812
rect 42433 -9035 42475 -9029
rect 41870 -9088 41912 -9054
rect 41966 -9088 42008 -9054
rect 42062 -9088 42104 -9054
rect 42966 -9076 42974 -8809
rect 43303 -8812 43304 -8742
rect 43337 -8819 43338 -8740
rect 43820 -8741 43833 -8673
rect 43861 -8707 43867 -8639
rect 43906 -8671 43912 -8603
rect 43940 -8637 43946 -8571
rect 43950 -8621 43992 -8587
rect 44151 -8666 44193 -8632
rect 43920 -8689 43928 -8681
rect 43931 -8723 43973 -8689
rect 44151 -8734 44193 -8700
rect 43820 -8753 43828 -8741
rect 44200 -8750 44206 -8616
rect 43595 -8819 43989 -8753
rect 44234 -8784 44240 -8590
rect 44274 -8606 44282 -8595
rect 44270 -8637 44282 -8606
rect 44596 -8624 44638 -8590
rect 42982 -8860 43024 -8826
rect 43331 -8830 43349 -8819
rect 43331 -8832 43338 -8830
rect 42982 -8928 43024 -8894
rect 43034 -8995 43040 -8860
rect 43265 -8874 43338 -8832
rect 43393 -8874 43989 -8819
rect 44129 -8853 44171 -8819
rect 44174 -8853 44182 -8808
rect 44270 -8820 44276 -8637
rect 44304 -8823 44310 -8640
rect 43265 -8877 43989 -8874
rect 43068 -8980 43074 -8892
rect 43185 -8942 43227 -8908
rect 43230 -8942 43238 -8900
rect 43066 -8991 43074 -8980
rect 43068 -9025 43074 -8991
rect 43077 -9025 43119 -8991
rect 43185 -9042 43227 -9008
rect 43230 -9042 43238 -8997
rect 43078 -9078 43120 -9044
rect 43150 -9078 43192 -9044
rect 43222 -9078 43264 -9044
rect 42224 -9131 42266 -9097
rect 42320 -9131 42362 -9097
rect 42416 -9131 42458 -9097
rect 42512 -9131 42554 -9097
rect 42608 -9131 42650 -9097
rect 43265 -9114 43417 -8877
rect 43595 -8899 43989 -8877
rect 43519 -8925 43989 -8899
rect 44316 -8904 44324 -8637
rect 44653 -8640 44654 -8570
rect 44332 -8688 44374 -8654
rect 44687 -8674 44688 -8568
rect 44881 -8577 44923 -8543
rect 44926 -8577 44934 -8532
rect 45026 -8543 45034 -8532
rect 45235 -8537 45277 -8503
rect 45280 -8537 45288 -8492
rect 45380 -8503 45388 -8492
rect 45625 -8496 45667 -8462
rect 45670 -8496 45678 -8451
rect 45391 -8537 45433 -8503
rect 45037 -8577 45079 -8543
rect 44332 -8756 44374 -8722
rect 44384 -8823 44390 -8688
rect 44946 -8691 44988 -8657
rect 44998 -8718 45004 -8641
rect 44418 -8808 44424 -8720
rect 44535 -8770 44577 -8736
rect 44580 -8770 44588 -8728
rect 44680 -8740 44688 -8729
rect 44691 -8774 44733 -8740
rect 45032 -8752 45038 -8607
rect 45235 -8620 45277 -8586
rect 45280 -8620 45288 -8575
rect 45380 -8586 45388 -8575
rect 45625 -8580 45667 -8546
rect 45670 -8580 45678 -8535
rect 45391 -8620 45433 -8586
rect 45300 -8734 45342 -8700
rect 45352 -8761 45358 -8684
rect 44416 -8819 44424 -8808
rect 44885 -8813 44927 -8779
rect 44930 -8813 44938 -8771
rect 45030 -8779 45038 -8771
rect 45041 -8813 45083 -8779
rect 45386 -8795 45392 -8650
rect 45625 -8663 45667 -8629
rect 45670 -8663 45678 -8618
rect 45747 -8679 45753 -8413
rect 45781 -8413 45823 -8379
rect 45826 -8413 45834 -8371
rect 45770 -8462 45778 -8451
rect 45781 -8462 45787 -8413
rect 45781 -8496 45823 -8462
rect 45826 -8496 45834 -8451
rect 45770 -8546 45778 -8535
rect 45781 -8546 45787 -8496
rect 45781 -8580 45823 -8546
rect 45826 -8580 45834 -8535
rect 45770 -8629 45778 -8618
rect 45781 -8629 45787 -8580
rect 45781 -8663 45823 -8629
rect 45826 -8663 45834 -8618
rect 45770 -8697 45778 -8671
rect 45781 -8713 45787 -8663
rect 45690 -8777 45732 -8743
rect 45747 -8804 45748 -8727
rect 45781 -8809 45782 -8713
rect 44418 -8853 44424 -8819
rect 44427 -8853 44469 -8819
rect 44535 -8870 44577 -8836
rect 44580 -8870 44588 -8825
rect 44680 -8832 44688 -8821
rect 44691 -8866 44733 -8832
rect 45239 -8856 45281 -8822
rect 45284 -8856 45292 -8814
rect 45384 -8822 45392 -8814
rect 45395 -8856 45437 -8822
rect 45812 -8845 45820 -8697
rect 45835 -8713 45839 -8363
rect 45869 -8679 45873 -8363
rect 45926 -8379 45934 -8371
rect 45875 -8413 45917 -8379
rect 45937 -8413 45989 -8379
rect 46647 -8422 46653 -8406
rect 46670 -8422 46678 -8414
rect 46681 -8422 46687 -8406
rect 46977 -8408 47019 -8374
rect 47022 -8408 47030 -8363
rect 45926 -8462 45934 -8451
rect 46107 -8456 46149 -8422
rect 46179 -8456 46221 -8422
rect 46251 -8456 46293 -8422
rect 46395 -8456 46437 -8422
rect 46467 -8456 46581 -8422
rect 46611 -8456 46653 -8422
rect 45937 -8496 45979 -8462
rect 45926 -8546 45934 -8535
rect 46504 -8539 46546 -8505
rect 45937 -8580 45979 -8546
rect 45926 -8629 45934 -8618
rect 45937 -8663 45979 -8629
rect 46169 -8689 46211 -8655
rect 46214 -8689 46222 -8644
rect 46291 -8706 46297 -8588
rect 46314 -8655 46322 -8644
rect 46325 -8655 46331 -8622
rect 46361 -8655 46367 -8622
rect 46325 -8689 46367 -8655
rect 46370 -8689 46378 -8644
rect 46325 -8740 46331 -8689
rect 46361 -8740 46367 -8689
rect 46395 -8706 46401 -8589
rect 46492 -8630 46493 -8589
rect 46504 -8623 46546 -8589
rect 46504 -8706 46546 -8672
rect 46647 -8706 46653 -8456
rect 46681 -8456 46723 -8422
rect 46670 -8505 46678 -8494
rect 46681 -8505 46687 -8456
rect 46977 -8491 47019 -8457
rect 47022 -8491 47030 -8446
rect 46681 -8539 46723 -8505
rect 46670 -8589 46678 -8578
rect 46681 -8589 46687 -8539
rect 46831 -8565 46939 -8499
rect 47099 -8507 47105 -8241
rect 47133 -8241 47175 -8207
rect 47178 -8241 47186 -8199
rect 47122 -8290 47130 -8279
rect 47133 -8290 47139 -8241
rect 47133 -8324 47175 -8290
rect 47178 -8324 47186 -8279
rect 47122 -8374 47130 -8363
rect 47133 -8374 47139 -8324
rect 47133 -8408 47175 -8374
rect 47178 -8408 47186 -8363
rect 47122 -8457 47130 -8446
rect 47133 -8457 47139 -8408
rect 47133 -8491 47175 -8457
rect 47178 -8491 47186 -8446
rect 47122 -8525 47130 -8499
rect 47133 -8541 47139 -8491
rect 46681 -8623 46723 -8589
rect 47042 -8605 47084 -8571
rect 46670 -8672 46678 -8661
rect 46681 -8672 46687 -8623
rect 47099 -8632 47100 -8555
rect 47133 -8637 47134 -8541
rect 46681 -8706 46723 -8672
rect 47164 -8673 47172 -8525
rect 47187 -8541 47191 -8191
rect 47221 -8507 47225 -8191
rect 47278 -8207 47286 -8199
rect 47227 -8241 47269 -8207
rect 47289 -8241 47341 -8207
rect 48204 -8231 48246 -8197
rect 48300 -8231 48342 -8197
rect 48396 -8231 48438 -8197
rect 50366 -8207 50374 -8199
rect 50443 -8207 50449 -8191
rect 50466 -8207 50474 -8199
rect 50477 -8207 50483 -8191
rect 47997 -8250 48003 -8234
rect 48020 -8250 48028 -8242
rect 48031 -8250 48037 -8234
rect 47278 -8290 47286 -8279
rect 47457 -8284 47499 -8250
rect 47529 -8284 47571 -8250
rect 47601 -8284 47643 -8250
rect 47745 -8284 47787 -8250
rect 47817 -8284 47931 -8250
rect 47961 -8284 48003 -8250
rect 47289 -8324 47331 -8290
rect 47278 -8374 47286 -8363
rect 47854 -8367 47896 -8333
rect 47289 -8408 47331 -8374
rect 47278 -8457 47286 -8446
rect 47289 -8491 47331 -8457
rect 47519 -8517 47561 -8483
rect 47564 -8517 47572 -8472
rect 47641 -8534 47647 -8416
rect 47664 -8483 47672 -8472
rect 47675 -8483 47681 -8450
rect 47711 -8483 47717 -8450
rect 47675 -8517 47717 -8483
rect 47720 -8517 47728 -8472
rect 47675 -8568 47681 -8517
rect 47711 -8568 47717 -8517
rect 47745 -8534 47751 -8417
rect 47842 -8458 47843 -8417
rect 47854 -8451 47896 -8417
rect 47854 -8534 47896 -8500
rect 47997 -8534 48003 -8284
rect 48031 -8284 48073 -8250
rect 48558 -8274 48600 -8240
rect 48654 -8274 48696 -8240
rect 48750 -8274 48792 -8240
rect 50257 -8241 50299 -8207
rect 50321 -8241 50374 -8207
rect 50401 -8241 50449 -8207
rect 48020 -8333 48028 -8322
rect 48031 -8333 48037 -8284
rect 48270 -8293 48278 -8285
rect 48370 -8293 48378 -8285
rect 48197 -8327 48267 -8293
rect 48269 -8327 48311 -8293
rect 48381 -8327 48423 -8293
rect 48912 -8317 48954 -8283
rect 49008 -8317 49050 -8283
rect 49104 -8317 49146 -8283
rect 49200 -8317 49242 -8283
rect 49296 -8317 49338 -8283
rect 50321 -8324 50363 -8290
rect 50366 -8324 50374 -8279
rect 48031 -8367 48073 -8333
rect 48624 -8336 48632 -8328
rect 48724 -8336 48732 -8328
rect 48020 -8417 48028 -8406
rect 48031 -8417 48037 -8367
rect 48225 -8410 48267 -8376
rect 48270 -8410 48278 -8365
rect 48370 -8376 48378 -8365
rect 48551 -8370 48621 -8336
rect 48623 -8370 48665 -8336
rect 48735 -8370 48777 -8336
rect 49460 -8360 49502 -8326
rect 49556 -8360 49598 -8326
rect 49652 -8360 49694 -8326
rect 49748 -8360 49790 -8326
rect 49844 -8360 49886 -8326
rect 49940 -8360 49982 -8326
rect 50036 -8360 50078 -8326
rect 48381 -8410 48423 -8376
rect 49014 -8379 49022 -8371
rect 49091 -8379 49097 -8363
rect 49114 -8379 49122 -8371
rect 49125 -8379 49131 -8363
rect 48031 -8451 48073 -8417
rect 48020 -8500 48028 -8489
rect 48031 -8500 48037 -8451
rect 48225 -8494 48267 -8460
rect 48270 -8494 48278 -8449
rect 48370 -8460 48378 -8449
rect 48579 -8453 48621 -8419
rect 48624 -8453 48632 -8408
rect 48724 -8419 48732 -8408
rect 48905 -8413 48947 -8379
rect 48969 -8413 49022 -8379
rect 49049 -8413 49097 -8379
rect 48735 -8453 48777 -8419
rect 48381 -8494 48423 -8460
rect 48031 -8534 48073 -8500
rect 48031 -8568 48037 -8534
rect 46681 -8740 46687 -8706
rect 46977 -8723 47019 -8689
rect 47022 -8723 47030 -8681
rect 44428 -8906 44470 -8872
rect 44500 -8906 44542 -8872
rect 44572 -8906 44614 -8872
rect 44885 -8913 44927 -8879
rect 44930 -8913 44938 -8868
rect 45030 -8879 45038 -8868
rect 45041 -8913 45083 -8879
rect 45625 -8895 45667 -8861
rect 45670 -8895 45678 -8853
rect 43519 -8959 44002 -8925
rect 44853 -8949 44895 -8915
rect 44925 -8949 44967 -8915
rect 45239 -8956 45281 -8922
rect 45284 -8956 45292 -8911
rect 45384 -8922 45392 -8911
rect 45812 -8913 45825 -8845
rect 45853 -8879 45859 -8811
rect 45898 -8843 45904 -8775
rect 45932 -8809 45938 -8743
rect 45942 -8793 45984 -8759
rect 46145 -8838 46187 -8804
rect 45912 -8861 45920 -8853
rect 45923 -8895 45965 -8861
rect 46145 -8906 46187 -8872
rect 45395 -8956 45437 -8922
rect 43519 -8985 43989 -8959
rect 43523 -8993 43731 -8985
rect 43539 -9003 43715 -8993
rect 43265 -9140 43447 -9114
rect 42772 -9174 42814 -9140
rect 42868 -9174 42910 -9140
rect 42964 -9174 43006 -9140
rect 43060 -9174 43102 -9140
rect 43156 -9174 43198 -9140
rect 43252 -9174 43447 -9140
rect 43265 -9200 43447 -9174
rect 43465 -9174 43573 -9050
rect 43724 -9062 43731 -9051
rect 43343 -9870 43385 -9200
rect 43465 -9228 43475 -9174
rect 43150 -9936 43302 -9924
rect 42818 -9970 43302 -9936
rect 43150 -9971 43302 -9970
rect 43331 -9971 43385 -9870
rect 43477 -9971 43519 -9174
rect 43523 -9971 43530 -9174
rect 43735 -9971 43777 -9062
rect 43869 -9971 43911 -8985
rect 44122 -9002 44164 -8968
rect 44218 -9002 44260 -8968
rect 44314 -9002 44356 -8968
rect 44410 -9002 44452 -8968
rect 44506 -9002 44548 -8968
rect 44602 -9002 44644 -8968
rect 44698 -9002 44740 -8968
rect 45207 -8992 45249 -8958
rect 45279 -8992 45321 -8958
rect 45625 -8995 45667 -8961
rect 45670 -8995 45678 -8950
rect 45812 -9001 45820 -8913
rect 46194 -8922 46200 -8788
rect 45912 -8961 45920 -8950
rect 46228 -8956 46234 -8762
rect 46268 -8778 46276 -8767
rect 46264 -8809 46276 -8778
rect 46590 -8796 46632 -8762
rect 45923 -8995 45965 -8961
rect 44860 -9045 44902 -9011
rect 44956 -9045 44998 -9011
rect 45052 -9045 45094 -9011
rect 45561 -9035 45603 -9001
rect 45633 -9035 45675 -9001
rect 45705 -9035 45747 -9001
rect 45777 -9029 45820 -9001
rect 46123 -9025 46165 -8991
rect 46168 -9025 46176 -8980
rect 46264 -8992 46270 -8809
rect 46298 -8995 46304 -8812
rect 45777 -9035 45819 -9029
rect 45214 -9088 45256 -9054
rect 45310 -9088 45352 -9054
rect 45406 -9088 45448 -9054
rect 46310 -9076 46318 -8809
rect 46647 -8812 46648 -8742
rect 46681 -8819 46682 -8740
rect 47164 -8741 47177 -8673
rect 47205 -8707 47211 -8639
rect 47250 -8671 47256 -8603
rect 47284 -8637 47290 -8571
rect 47294 -8621 47336 -8587
rect 47495 -8666 47537 -8632
rect 47264 -8689 47272 -8681
rect 47275 -8723 47317 -8689
rect 47495 -8734 47537 -8700
rect 47164 -8753 47172 -8741
rect 47544 -8750 47550 -8616
rect 46939 -8819 47333 -8753
rect 47578 -8784 47584 -8590
rect 47618 -8606 47626 -8595
rect 47614 -8637 47626 -8606
rect 47940 -8624 47982 -8590
rect 46326 -8860 46368 -8826
rect 46675 -8830 46693 -8819
rect 46675 -8832 46682 -8830
rect 46326 -8928 46368 -8894
rect 46378 -8995 46384 -8860
rect 46609 -8874 46682 -8832
rect 46737 -8874 47333 -8819
rect 47473 -8853 47515 -8819
rect 47518 -8853 47526 -8808
rect 47614 -8820 47620 -8637
rect 47648 -8823 47654 -8640
rect 46609 -8877 47333 -8874
rect 46412 -8980 46418 -8892
rect 46529 -8942 46571 -8908
rect 46574 -8942 46582 -8900
rect 46410 -8991 46418 -8980
rect 46412 -9025 46418 -8991
rect 46421 -9025 46463 -8991
rect 46529 -9042 46571 -9008
rect 46574 -9042 46582 -8997
rect 46422 -9078 46464 -9044
rect 46494 -9078 46536 -9044
rect 46566 -9078 46608 -9044
rect 45568 -9131 45610 -9097
rect 45664 -9131 45706 -9097
rect 45760 -9131 45802 -9097
rect 45856 -9131 45898 -9097
rect 45952 -9131 45994 -9097
rect 46609 -9114 46761 -8877
rect 46939 -8899 47333 -8877
rect 46863 -8925 47333 -8899
rect 47660 -8904 47668 -8637
rect 47997 -8640 47998 -8570
rect 47676 -8688 47718 -8654
rect 48031 -8674 48032 -8568
rect 48225 -8577 48267 -8543
rect 48270 -8577 48278 -8532
rect 48370 -8543 48378 -8532
rect 48579 -8537 48621 -8503
rect 48624 -8537 48632 -8492
rect 48724 -8503 48732 -8492
rect 48969 -8496 49011 -8462
rect 49014 -8496 49022 -8451
rect 48735 -8537 48777 -8503
rect 48381 -8577 48423 -8543
rect 47676 -8756 47718 -8722
rect 47728 -8823 47734 -8688
rect 48290 -8691 48332 -8657
rect 48342 -8718 48348 -8641
rect 47762 -8808 47768 -8720
rect 47879 -8770 47921 -8736
rect 47924 -8770 47932 -8728
rect 48024 -8740 48032 -8729
rect 48035 -8774 48077 -8740
rect 48376 -8752 48382 -8607
rect 48579 -8620 48621 -8586
rect 48624 -8620 48632 -8575
rect 48724 -8586 48732 -8575
rect 48969 -8580 49011 -8546
rect 49014 -8580 49022 -8535
rect 48735 -8620 48777 -8586
rect 48644 -8734 48686 -8700
rect 48696 -8761 48702 -8684
rect 47760 -8819 47768 -8808
rect 48229 -8813 48271 -8779
rect 48274 -8813 48282 -8771
rect 48374 -8779 48382 -8771
rect 48385 -8813 48427 -8779
rect 48730 -8795 48736 -8650
rect 48969 -8663 49011 -8629
rect 49014 -8663 49022 -8618
rect 49091 -8679 49097 -8413
rect 49125 -8413 49167 -8379
rect 49170 -8413 49178 -8371
rect 49114 -8462 49122 -8451
rect 49125 -8462 49131 -8413
rect 49125 -8496 49167 -8462
rect 49170 -8496 49178 -8451
rect 49114 -8546 49122 -8535
rect 49125 -8546 49131 -8496
rect 49125 -8580 49167 -8546
rect 49170 -8580 49178 -8535
rect 49114 -8629 49122 -8618
rect 49125 -8629 49131 -8580
rect 49125 -8663 49167 -8629
rect 49170 -8663 49178 -8618
rect 49114 -8697 49122 -8671
rect 49125 -8713 49131 -8663
rect 49034 -8777 49076 -8743
rect 49091 -8804 49092 -8727
rect 49125 -8809 49126 -8713
rect 47762 -8853 47768 -8819
rect 47771 -8853 47813 -8819
rect 47879 -8870 47921 -8836
rect 47924 -8870 47932 -8825
rect 48024 -8832 48032 -8821
rect 48035 -8866 48077 -8832
rect 48583 -8856 48625 -8822
rect 48628 -8856 48636 -8814
rect 48728 -8822 48736 -8814
rect 48739 -8856 48781 -8822
rect 49156 -8845 49164 -8697
rect 49179 -8713 49183 -8363
rect 49213 -8679 49217 -8363
rect 49270 -8379 49278 -8371
rect 49219 -8413 49261 -8379
rect 49281 -8413 49333 -8379
rect 49991 -8422 49997 -8406
rect 50014 -8422 50022 -8414
rect 50025 -8422 50031 -8406
rect 50321 -8408 50363 -8374
rect 50366 -8408 50374 -8363
rect 49270 -8462 49278 -8451
rect 49451 -8456 49493 -8422
rect 49523 -8456 49565 -8422
rect 49595 -8456 49637 -8422
rect 49739 -8456 49781 -8422
rect 49811 -8456 49925 -8422
rect 49955 -8456 49997 -8422
rect 49281 -8496 49323 -8462
rect 49270 -8546 49278 -8535
rect 49848 -8539 49890 -8505
rect 49281 -8580 49323 -8546
rect 49270 -8629 49278 -8618
rect 49281 -8663 49323 -8629
rect 49513 -8689 49555 -8655
rect 49558 -8689 49566 -8644
rect 49635 -8706 49641 -8588
rect 49658 -8655 49666 -8644
rect 49669 -8655 49675 -8622
rect 49705 -8655 49711 -8622
rect 49669 -8689 49711 -8655
rect 49714 -8689 49722 -8644
rect 49669 -8740 49675 -8689
rect 49705 -8740 49711 -8689
rect 49739 -8706 49745 -8589
rect 49836 -8630 49837 -8589
rect 49848 -8623 49890 -8589
rect 49848 -8706 49890 -8672
rect 49991 -8706 49997 -8456
rect 50025 -8456 50067 -8422
rect 50014 -8505 50022 -8494
rect 50025 -8505 50031 -8456
rect 50321 -8491 50363 -8457
rect 50366 -8491 50374 -8446
rect 50025 -8539 50067 -8505
rect 50014 -8589 50022 -8578
rect 50025 -8589 50031 -8539
rect 50175 -8565 50283 -8499
rect 50443 -8507 50449 -8241
rect 50477 -8241 50519 -8207
rect 50522 -8241 50530 -8199
rect 50466 -8290 50474 -8279
rect 50477 -8290 50483 -8241
rect 50477 -8324 50519 -8290
rect 50522 -8324 50530 -8279
rect 50466 -8374 50474 -8363
rect 50477 -8374 50483 -8324
rect 50477 -8408 50519 -8374
rect 50522 -8408 50530 -8363
rect 50466 -8457 50474 -8446
rect 50477 -8457 50483 -8408
rect 50477 -8491 50519 -8457
rect 50522 -8491 50530 -8446
rect 50466 -8525 50474 -8499
rect 50477 -8541 50483 -8491
rect 50025 -8623 50067 -8589
rect 50386 -8605 50428 -8571
rect 50014 -8672 50022 -8661
rect 50025 -8672 50031 -8623
rect 50443 -8632 50444 -8555
rect 50477 -8637 50478 -8541
rect 50025 -8706 50067 -8672
rect 50508 -8673 50516 -8525
rect 50531 -8541 50535 -8191
rect 50565 -8507 50569 -8191
rect 50622 -8207 50630 -8199
rect 50571 -8241 50613 -8207
rect 50633 -8241 50685 -8207
rect 51548 -8231 51590 -8197
rect 51644 -8231 51686 -8197
rect 51740 -8231 51782 -8197
rect 53711 -8207 53718 -8199
rect 51341 -8250 51347 -8234
rect 51364 -8250 51372 -8242
rect 51375 -8250 51381 -8234
rect 50622 -8290 50630 -8279
rect 50801 -8284 50843 -8250
rect 50873 -8284 50915 -8250
rect 50945 -8284 50987 -8250
rect 51089 -8284 51131 -8250
rect 51161 -8284 51275 -8250
rect 51305 -8284 51347 -8250
rect 50633 -8324 50675 -8290
rect 50622 -8374 50630 -8363
rect 51198 -8367 51240 -8333
rect 50633 -8408 50675 -8374
rect 50622 -8457 50630 -8446
rect 50633 -8491 50675 -8457
rect 50863 -8517 50905 -8483
rect 50908 -8517 50916 -8472
rect 50985 -8534 50991 -8416
rect 51008 -8483 51016 -8472
rect 51019 -8483 51025 -8450
rect 51055 -8483 51061 -8450
rect 51019 -8517 51061 -8483
rect 51064 -8517 51072 -8472
rect 51019 -8568 51025 -8517
rect 51055 -8568 51061 -8517
rect 51089 -8534 51095 -8417
rect 51186 -8458 51187 -8417
rect 51198 -8451 51240 -8417
rect 51198 -8534 51240 -8500
rect 51341 -8534 51347 -8284
rect 51375 -8284 51417 -8250
rect 51902 -8274 51944 -8240
rect 51998 -8274 52040 -8240
rect 52094 -8274 52136 -8240
rect 53602 -8241 53643 -8207
rect 53666 -8241 53718 -8207
rect 53746 -8241 53787 -8207
rect 51364 -8333 51372 -8322
rect 51375 -8333 51381 -8284
rect 51614 -8293 51622 -8285
rect 51714 -8293 51722 -8285
rect 51541 -8327 51611 -8293
rect 51613 -8327 51655 -8293
rect 51725 -8327 51767 -8293
rect 52256 -8317 52298 -8283
rect 52352 -8317 52394 -8283
rect 52448 -8317 52490 -8283
rect 52544 -8317 52586 -8283
rect 52640 -8317 52682 -8283
rect 53666 -8324 53707 -8290
rect 53711 -8324 53718 -8279
rect 51375 -8367 51417 -8333
rect 51968 -8336 51976 -8328
rect 52068 -8336 52076 -8328
rect 51364 -8417 51372 -8406
rect 51375 -8417 51381 -8367
rect 51569 -8410 51611 -8376
rect 51614 -8410 51622 -8365
rect 51714 -8376 51722 -8365
rect 51895 -8370 51965 -8336
rect 51967 -8370 52009 -8336
rect 52079 -8370 52121 -8336
rect 52804 -8360 52846 -8326
rect 52900 -8360 52942 -8326
rect 52996 -8360 53038 -8326
rect 53092 -8360 53134 -8326
rect 53188 -8360 53230 -8326
rect 53284 -8360 53326 -8326
rect 53380 -8360 53422 -8326
rect 51725 -8410 51767 -8376
rect 52358 -8379 52366 -8371
rect 52435 -8379 52441 -8363
rect 52458 -8379 52466 -8371
rect 52469 -8379 52475 -8363
rect 51375 -8451 51417 -8417
rect 51364 -8500 51372 -8489
rect 51375 -8500 51381 -8451
rect 51569 -8494 51611 -8460
rect 51614 -8494 51622 -8449
rect 51714 -8460 51722 -8449
rect 51923 -8453 51965 -8419
rect 51968 -8453 51976 -8408
rect 52068 -8419 52076 -8408
rect 52249 -8413 52291 -8379
rect 52313 -8413 52366 -8379
rect 52393 -8413 52441 -8379
rect 52079 -8453 52121 -8419
rect 51725 -8494 51767 -8460
rect 51375 -8534 51417 -8500
rect 51375 -8568 51381 -8534
rect 50025 -8740 50031 -8706
rect 50321 -8723 50363 -8689
rect 50366 -8723 50374 -8681
rect 47772 -8906 47814 -8872
rect 47844 -8906 47886 -8872
rect 47916 -8906 47958 -8872
rect 48229 -8913 48271 -8879
rect 48274 -8913 48282 -8868
rect 48374 -8879 48382 -8868
rect 48385 -8913 48427 -8879
rect 48969 -8895 49011 -8861
rect 49014 -8895 49022 -8853
rect 46863 -8959 47346 -8925
rect 48197 -8949 48239 -8915
rect 48269 -8949 48311 -8915
rect 48583 -8956 48625 -8922
rect 48628 -8956 48636 -8911
rect 48728 -8922 48736 -8911
rect 49156 -8913 49169 -8845
rect 49197 -8879 49203 -8811
rect 49242 -8843 49248 -8775
rect 49276 -8809 49282 -8743
rect 49286 -8793 49328 -8759
rect 49489 -8838 49531 -8804
rect 49256 -8861 49264 -8853
rect 49267 -8895 49309 -8861
rect 49489 -8906 49531 -8872
rect 48739 -8956 48781 -8922
rect 46863 -8985 47333 -8959
rect 46867 -8993 47075 -8985
rect 46883 -9003 47059 -8993
rect 46609 -9140 46791 -9114
rect 46116 -9174 46158 -9140
rect 46212 -9174 46254 -9140
rect 46308 -9174 46350 -9140
rect 46404 -9174 46446 -9140
rect 46500 -9174 46542 -9140
rect 46596 -9174 46791 -9140
rect 46609 -9200 46791 -9174
rect 46809 -9174 46917 -9050
rect 47068 -9062 47075 -9051
rect 46687 -9870 46729 -9200
rect 46809 -9228 46819 -9174
rect 46494 -9936 46646 -9924
rect 46162 -9970 46646 -9936
rect 46494 -9971 46646 -9970
rect 46675 -9971 46729 -9870
rect 46821 -9971 46863 -9174
rect 46867 -9971 46874 -9174
rect 47079 -9971 47121 -9062
rect 47213 -9971 47255 -8985
rect 47466 -9002 47508 -8968
rect 47562 -9002 47604 -8968
rect 47658 -9002 47700 -8968
rect 47754 -9002 47796 -8968
rect 47850 -9002 47892 -8968
rect 47946 -9002 47988 -8968
rect 48042 -9002 48084 -8968
rect 48551 -8992 48593 -8958
rect 48623 -8992 48665 -8958
rect 48969 -8995 49011 -8961
rect 49014 -8995 49022 -8950
rect 49156 -9001 49164 -8913
rect 49538 -8922 49544 -8788
rect 49256 -8961 49264 -8950
rect 49572 -8956 49578 -8762
rect 49612 -8778 49620 -8767
rect 49608 -8809 49620 -8778
rect 49934 -8796 49976 -8762
rect 49267 -8995 49309 -8961
rect 48204 -9045 48246 -9011
rect 48300 -9045 48342 -9011
rect 48396 -9045 48438 -9011
rect 48905 -9035 48947 -9001
rect 48977 -9035 49019 -9001
rect 49049 -9035 49091 -9001
rect 49121 -9029 49164 -9001
rect 49467 -9025 49509 -8991
rect 49512 -9025 49520 -8980
rect 49608 -8992 49614 -8809
rect 49642 -8995 49648 -8812
rect 49121 -9035 49163 -9029
rect 48558 -9088 48600 -9054
rect 48654 -9088 48696 -9054
rect 48750 -9088 48792 -9054
rect 49654 -9076 49662 -8809
rect 49991 -8812 49992 -8742
rect 50025 -8819 50026 -8740
rect 50508 -8741 50521 -8673
rect 50549 -8707 50555 -8639
rect 50594 -8671 50600 -8603
rect 50628 -8637 50634 -8571
rect 50638 -8621 50680 -8587
rect 50839 -8666 50881 -8632
rect 50608 -8689 50616 -8681
rect 50619 -8723 50661 -8689
rect 50839 -8734 50881 -8700
rect 50508 -8753 50516 -8741
rect 50888 -8750 50894 -8616
rect 50283 -8819 50677 -8753
rect 50922 -8784 50928 -8590
rect 50962 -8606 50970 -8595
rect 50958 -8637 50970 -8606
rect 51284 -8624 51326 -8590
rect 49670 -8860 49712 -8826
rect 50019 -8830 50037 -8819
rect 50019 -8832 50026 -8830
rect 49670 -8928 49712 -8894
rect 49722 -8995 49728 -8860
rect 49953 -8874 50026 -8832
rect 50081 -8874 50677 -8819
rect 50817 -8853 50859 -8819
rect 50862 -8853 50870 -8808
rect 50958 -8820 50964 -8637
rect 50992 -8823 50998 -8640
rect 49953 -8877 50677 -8874
rect 49756 -8980 49762 -8892
rect 49873 -8942 49915 -8908
rect 49918 -8942 49926 -8900
rect 49754 -8991 49762 -8980
rect 49756 -9025 49762 -8991
rect 49765 -9025 49807 -8991
rect 49873 -9042 49915 -9008
rect 49918 -9042 49926 -8997
rect 49766 -9078 49808 -9044
rect 49838 -9078 49880 -9044
rect 49910 -9078 49952 -9044
rect 48912 -9131 48954 -9097
rect 49008 -9131 49050 -9097
rect 49104 -9131 49146 -9097
rect 49200 -9131 49242 -9097
rect 49296 -9131 49338 -9097
rect 49953 -9114 50105 -8877
rect 50283 -8899 50677 -8877
rect 50207 -8925 50677 -8899
rect 51004 -8904 51012 -8637
rect 51341 -8640 51342 -8570
rect 51020 -8688 51062 -8654
rect 51375 -8674 51376 -8568
rect 51569 -8577 51611 -8543
rect 51614 -8577 51622 -8532
rect 51714 -8543 51722 -8532
rect 51923 -8537 51965 -8503
rect 51968 -8537 51976 -8492
rect 52068 -8503 52076 -8492
rect 52313 -8496 52355 -8462
rect 52358 -8496 52366 -8451
rect 52079 -8537 52121 -8503
rect 51725 -8577 51767 -8543
rect 51020 -8756 51062 -8722
rect 51072 -8823 51078 -8688
rect 51634 -8691 51676 -8657
rect 51686 -8718 51692 -8641
rect 51106 -8808 51112 -8720
rect 51223 -8770 51265 -8736
rect 51268 -8770 51276 -8728
rect 51368 -8740 51376 -8729
rect 51379 -8774 51421 -8740
rect 51720 -8752 51726 -8607
rect 51923 -8620 51965 -8586
rect 51968 -8620 51976 -8575
rect 52068 -8586 52076 -8575
rect 52313 -8580 52355 -8546
rect 52358 -8580 52366 -8535
rect 52079 -8620 52121 -8586
rect 51988 -8734 52030 -8700
rect 52040 -8761 52046 -8684
rect 51104 -8819 51112 -8808
rect 51573 -8813 51615 -8779
rect 51618 -8813 51626 -8771
rect 51718 -8779 51726 -8771
rect 51729 -8813 51771 -8779
rect 52074 -8795 52080 -8650
rect 52313 -8663 52355 -8629
rect 52358 -8663 52366 -8618
rect 52435 -8679 52441 -8413
rect 52469 -8413 52511 -8379
rect 52514 -8413 52522 -8371
rect 52458 -8462 52466 -8451
rect 52469 -8462 52475 -8413
rect 52469 -8496 52511 -8462
rect 52514 -8496 52522 -8451
rect 52458 -8546 52466 -8535
rect 52469 -8546 52475 -8496
rect 52469 -8580 52511 -8546
rect 52514 -8580 52522 -8535
rect 52458 -8629 52466 -8618
rect 52469 -8629 52475 -8580
rect 52469 -8663 52511 -8629
rect 52514 -8663 52522 -8618
rect 52458 -8697 52466 -8671
rect 52469 -8713 52475 -8663
rect 52378 -8777 52420 -8743
rect 52435 -8804 52436 -8727
rect 52469 -8809 52470 -8713
rect 51106 -8853 51112 -8819
rect 51115 -8853 51157 -8819
rect 51223 -8870 51265 -8836
rect 51268 -8870 51276 -8825
rect 51368 -8832 51376 -8821
rect 51379 -8866 51421 -8832
rect 51927 -8856 51969 -8822
rect 51972 -8856 51980 -8814
rect 52072 -8822 52080 -8814
rect 52083 -8856 52125 -8822
rect 52500 -8845 52508 -8697
rect 52523 -8713 52527 -8363
rect 52557 -8679 52561 -8363
rect 52614 -8379 52622 -8371
rect 52563 -8413 52605 -8379
rect 52625 -8413 52677 -8379
rect 53335 -8422 53341 -8406
rect 53358 -8422 53366 -8414
rect 53369 -8422 53375 -8406
rect 53666 -8408 53707 -8374
rect 53711 -8408 53718 -8363
rect 52614 -8462 52622 -8451
rect 52795 -8456 52837 -8422
rect 52867 -8456 52909 -8422
rect 52939 -8456 52981 -8422
rect 53083 -8456 53125 -8422
rect 53155 -8456 53269 -8422
rect 53299 -8456 53341 -8422
rect 52625 -8496 52667 -8462
rect 52614 -8546 52622 -8535
rect 53192 -8539 53234 -8505
rect 52625 -8580 52667 -8546
rect 52614 -8629 52622 -8618
rect 52625 -8663 52667 -8629
rect 52857 -8689 52899 -8655
rect 52902 -8689 52910 -8644
rect 52979 -8706 52985 -8588
rect 53002 -8655 53010 -8644
rect 53013 -8655 53019 -8622
rect 53049 -8655 53055 -8622
rect 53013 -8689 53055 -8655
rect 53058 -8689 53066 -8644
rect 53013 -8740 53019 -8689
rect 53049 -8740 53055 -8689
rect 53083 -8706 53089 -8589
rect 53180 -8630 53181 -8589
rect 53192 -8623 53234 -8589
rect 53192 -8706 53234 -8672
rect 53335 -8706 53341 -8456
rect 53369 -8456 53411 -8422
rect 53358 -8505 53366 -8494
rect 53369 -8505 53375 -8456
rect 53666 -8491 53707 -8457
rect 53711 -8491 53718 -8446
rect 53369 -8539 53411 -8505
rect 53358 -8589 53366 -8578
rect 53369 -8589 53375 -8539
rect 53519 -8565 53628 -8499
rect 53788 -8507 53793 -8191
rect 53811 -8207 53818 -8199
rect 53822 -8207 53827 -8191
rect 53822 -8241 53863 -8207
rect 53867 -8241 53874 -8199
rect 53811 -8290 53818 -8279
rect 53822 -8290 53827 -8241
rect 53822 -8324 53863 -8290
rect 53867 -8324 53874 -8279
rect 53811 -8374 53818 -8363
rect 53822 -8374 53827 -8324
rect 53822 -8408 53863 -8374
rect 53867 -8408 53874 -8363
rect 53811 -8457 53818 -8446
rect 53822 -8457 53827 -8408
rect 53822 -8491 53863 -8457
rect 53867 -8491 53874 -8446
rect 53811 -8525 53818 -8499
rect 53822 -8541 53827 -8491
rect 53369 -8623 53411 -8589
rect 53731 -8605 53772 -8571
rect 53358 -8672 53366 -8661
rect 53369 -8672 53375 -8623
rect 53369 -8706 53411 -8672
rect 53853 -8673 53860 -8525
rect 53876 -8541 53879 -8191
rect 53910 -8507 53913 -8191
rect 53967 -8207 53974 -8199
rect 53916 -8241 53957 -8207
rect 53978 -8241 54029 -8207
rect 54893 -8231 54934 -8197
rect 54989 -8231 55030 -8197
rect 55085 -8231 55126 -8197
rect 57055 -8207 57062 -8199
rect 54686 -8250 54691 -8234
rect 54709 -8250 54716 -8242
rect 54720 -8250 54725 -8234
rect 53967 -8290 53974 -8279
rect 54146 -8284 54187 -8250
rect 54218 -8284 54259 -8250
rect 54290 -8284 54331 -8250
rect 54434 -8284 54475 -8250
rect 54506 -8284 54619 -8250
rect 54650 -8284 54691 -8250
rect 53978 -8324 54019 -8290
rect 53967 -8374 53974 -8363
rect 54543 -8367 54584 -8333
rect 53978 -8408 54019 -8374
rect 53967 -8457 53974 -8446
rect 53978 -8491 54019 -8457
rect 54208 -8517 54249 -8483
rect 54253 -8517 54260 -8472
rect 54330 -8534 54335 -8416
rect 54353 -8483 54360 -8472
rect 54364 -8483 54369 -8450
rect 54400 -8483 54405 -8450
rect 54364 -8517 54405 -8483
rect 54409 -8517 54416 -8472
rect 54364 -8568 54369 -8517
rect 54400 -8568 54405 -8517
rect 54434 -8534 54439 -8417
rect 54543 -8451 54584 -8417
rect 54543 -8534 54584 -8500
rect 54686 -8534 54691 -8284
rect 54720 -8284 54761 -8250
rect 55247 -8274 55288 -8240
rect 55343 -8274 55384 -8240
rect 55439 -8274 55480 -8240
rect 56946 -8241 56987 -8207
rect 57010 -8241 57062 -8207
rect 57090 -8241 57131 -8207
rect 54709 -8333 54716 -8322
rect 54720 -8333 54725 -8284
rect 54959 -8293 54966 -8285
rect 55059 -8293 55066 -8285
rect 54886 -8327 54955 -8293
rect 54958 -8327 54999 -8293
rect 55070 -8327 55111 -8293
rect 55601 -8317 55642 -8283
rect 55697 -8317 55738 -8283
rect 55793 -8317 55834 -8283
rect 55889 -8317 55930 -8283
rect 55985 -8317 56026 -8283
rect 57010 -8324 57051 -8290
rect 57055 -8324 57062 -8279
rect 54720 -8367 54761 -8333
rect 55313 -8336 55320 -8328
rect 55413 -8336 55420 -8328
rect 54709 -8417 54716 -8406
rect 54720 -8417 54725 -8367
rect 54914 -8410 54955 -8376
rect 54959 -8410 54966 -8365
rect 55059 -8376 55066 -8365
rect 55240 -8370 55309 -8336
rect 55312 -8370 55353 -8336
rect 55424 -8370 55465 -8336
rect 56149 -8360 56190 -8326
rect 56245 -8360 56286 -8326
rect 56341 -8360 56382 -8326
rect 56437 -8360 56478 -8326
rect 56533 -8360 56574 -8326
rect 56629 -8360 56670 -8326
rect 56725 -8360 56766 -8326
rect 55070 -8410 55111 -8376
rect 55703 -8379 55710 -8371
rect 54720 -8451 54761 -8417
rect 54709 -8500 54716 -8489
rect 54720 -8500 54725 -8451
rect 54914 -8494 54955 -8460
rect 54959 -8494 54966 -8449
rect 55059 -8460 55066 -8449
rect 55268 -8453 55309 -8419
rect 55313 -8453 55320 -8408
rect 55413 -8419 55420 -8408
rect 55594 -8413 55635 -8379
rect 55658 -8413 55710 -8379
rect 55738 -8413 55779 -8379
rect 55424 -8453 55465 -8419
rect 55070 -8494 55111 -8460
rect 54720 -8534 54761 -8500
rect 54720 -8568 54725 -8534
rect 53369 -8740 53375 -8706
rect 53666 -8723 53707 -8689
rect 53711 -8723 53718 -8681
rect 51116 -8906 51158 -8872
rect 51188 -8906 51230 -8872
rect 51260 -8906 51302 -8872
rect 51573 -8913 51615 -8879
rect 51618 -8913 51626 -8868
rect 51718 -8879 51726 -8868
rect 51729 -8913 51771 -8879
rect 52313 -8895 52355 -8861
rect 52358 -8895 52366 -8853
rect 50207 -8959 50690 -8925
rect 51541 -8949 51583 -8915
rect 51613 -8949 51655 -8915
rect 51927 -8956 51969 -8922
rect 51972 -8956 51980 -8911
rect 52072 -8922 52080 -8911
rect 52500 -8913 52513 -8845
rect 52541 -8879 52547 -8811
rect 52586 -8843 52592 -8775
rect 52620 -8809 52626 -8743
rect 52630 -8793 52672 -8759
rect 52833 -8838 52875 -8804
rect 52600 -8861 52608 -8853
rect 52611 -8895 52653 -8861
rect 52833 -8906 52875 -8872
rect 52083 -8956 52125 -8922
rect 50207 -8985 50677 -8959
rect 50211 -8993 50419 -8985
rect 50227 -9003 50403 -8993
rect 49953 -9140 50135 -9114
rect 49460 -9174 49502 -9140
rect 49556 -9174 49598 -9140
rect 49652 -9174 49694 -9140
rect 49748 -9174 49790 -9140
rect 49844 -9174 49886 -9140
rect 49940 -9174 50135 -9140
rect 49953 -9200 50135 -9174
rect 50153 -9174 50261 -9050
rect 50412 -9062 50419 -9051
rect 50031 -9870 50073 -9200
rect 50153 -9228 50163 -9174
rect 49838 -9936 49990 -9924
rect 49506 -9970 49990 -9936
rect 49838 -9971 49990 -9970
rect 50019 -9971 50073 -9870
rect 50165 -9971 50207 -9174
rect 50211 -9971 50218 -9174
rect 50423 -9971 50465 -9062
rect 50557 -9971 50599 -8985
rect 50810 -9002 50852 -8968
rect 50906 -9002 50948 -8968
rect 51002 -9002 51044 -8968
rect 51098 -9002 51140 -8968
rect 51194 -9002 51236 -8968
rect 51290 -9002 51332 -8968
rect 51386 -9002 51428 -8968
rect 51895 -8992 51937 -8958
rect 51967 -8992 52009 -8958
rect 52313 -8995 52355 -8961
rect 52358 -8995 52366 -8950
rect 52500 -9001 52508 -8913
rect 52882 -8922 52888 -8788
rect 52600 -8961 52608 -8950
rect 52916 -8956 52922 -8762
rect 52956 -8778 52964 -8767
rect 52952 -8809 52964 -8778
rect 53278 -8796 53320 -8762
rect 52611 -8995 52653 -8961
rect 51548 -9045 51590 -9011
rect 51644 -9045 51686 -9011
rect 51740 -9045 51782 -9011
rect 52249 -9035 52291 -9001
rect 52321 -9035 52363 -9001
rect 52393 -9035 52435 -9001
rect 52465 -9029 52508 -9001
rect 52811 -9025 52853 -8991
rect 52856 -9025 52864 -8980
rect 52952 -8992 52958 -8809
rect 52986 -8995 52992 -8812
rect 52465 -9035 52507 -9029
rect 51902 -9088 51944 -9054
rect 51998 -9088 52040 -9054
rect 52094 -9088 52136 -9054
rect 52998 -9076 53006 -8809
rect 53335 -8812 53336 -8742
rect 53369 -8819 53370 -8740
rect 53853 -8741 53865 -8673
rect 53894 -8707 53899 -8639
rect 53939 -8671 53944 -8603
rect 53973 -8637 53978 -8571
rect 54914 -8577 54955 -8543
rect 54959 -8577 54966 -8532
rect 55059 -8543 55066 -8532
rect 55268 -8537 55309 -8503
rect 55313 -8537 55320 -8492
rect 55413 -8503 55420 -8492
rect 55658 -8496 55699 -8462
rect 55703 -8496 55710 -8451
rect 55424 -8537 55465 -8503
rect 55070 -8577 55111 -8543
rect 53983 -8621 54024 -8587
rect 54184 -8666 54225 -8632
rect 53953 -8689 53960 -8681
rect 53964 -8723 54005 -8689
rect 54184 -8734 54225 -8700
rect 53853 -8753 53860 -8741
rect 54233 -8750 54238 -8616
rect 53628 -8819 54021 -8753
rect 54267 -8784 54272 -8590
rect 54307 -8606 54314 -8595
rect 54303 -8637 54314 -8606
rect 54629 -8624 54670 -8590
rect 53014 -8860 53056 -8826
rect 53363 -8830 53381 -8819
rect 53363 -8832 53370 -8830
rect 53014 -8928 53056 -8894
rect 53066 -8995 53072 -8860
rect 53297 -8874 53370 -8832
rect 53426 -8874 54021 -8819
rect 54162 -8853 54203 -8819
rect 54207 -8853 54214 -8808
rect 54303 -8820 54308 -8637
rect 54337 -8823 54342 -8640
rect 53297 -8877 54021 -8874
rect 53100 -8980 53106 -8892
rect 53217 -8942 53259 -8908
rect 53262 -8942 53270 -8900
rect 53098 -8991 53106 -8980
rect 53100 -9025 53106 -8991
rect 53109 -9025 53151 -8991
rect 53217 -9042 53259 -9008
rect 53262 -9042 53270 -8997
rect 53110 -9078 53152 -9044
rect 53182 -9078 53224 -9044
rect 53254 -9078 53296 -9044
rect 52256 -9131 52298 -9097
rect 52352 -9131 52394 -9097
rect 52448 -9131 52490 -9097
rect 52544 -9131 52586 -9097
rect 52640 -9131 52682 -9097
rect 53297 -9114 53449 -8877
rect 53628 -8899 54021 -8877
rect 53552 -8925 54021 -8899
rect 54349 -8904 54356 -8637
rect 54365 -8688 54406 -8654
rect 54365 -8756 54406 -8722
rect 54417 -8823 54422 -8688
rect 54979 -8691 55020 -8657
rect 55031 -8718 55036 -8641
rect 54451 -8808 54456 -8720
rect 54568 -8770 54609 -8736
rect 54613 -8770 54620 -8728
rect 54713 -8740 54720 -8729
rect 54724 -8774 54765 -8740
rect 55065 -8752 55070 -8607
rect 55268 -8620 55309 -8586
rect 55313 -8620 55320 -8575
rect 55413 -8586 55420 -8575
rect 55658 -8580 55699 -8546
rect 55703 -8580 55710 -8535
rect 55424 -8620 55465 -8586
rect 55333 -8734 55374 -8700
rect 55385 -8761 55390 -8684
rect 54449 -8819 54456 -8808
rect 54918 -8813 54959 -8779
rect 54963 -8813 54970 -8771
rect 55063 -8779 55070 -8771
rect 55074 -8813 55115 -8779
rect 55419 -8795 55424 -8650
rect 55658 -8663 55699 -8629
rect 55703 -8663 55710 -8618
rect 55780 -8679 55785 -8363
rect 55803 -8379 55810 -8371
rect 55814 -8379 55819 -8363
rect 55814 -8413 55855 -8379
rect 55859 -8413 55866 -8371
rect 55803 -8462 55810 -8451
rect 55814 -8462 55819 -8413
rect 55814 -8496 55855 -8462
rect 55859 -8496 55866 -8451
rect 55803 -8546 55810 -8535
rect 55814 -8546 55819 -8496
rect 55814 -8580 55855 -8546
rect 55859 -8580 55866 -8535
rect 55803 -8629 55810 -8618
rect 55814 -8629 55819 -8580
rect 55814 -8663 55855 -8629
rect 55859 -8663 55866 -8618
rect 55803 -8697 55810 -8671
rect 55814 -8713 55819 -8663
rect 55723 -8777 55764 -8743
rect 54451 -8853 54456 -8819
rect 54460 -8853 54501 -8819
rect 54568 -8870 54609 -8836
rect 54613 -8870 54620 -8825
rect 54713 -8832 54720 -8821
rect 54724 -8866 54765 -8832
rect 55272 -8856 55313 -8822
rect 55317 -8856 55324 -8814
rect 55417 -8822 55424 -8814
rect 55428 -8856 55469 -8822
rect 55845 -8845 55852 -8697
rect 55868 -8713 55871 -8363
rect 55902 -8679 55905 -8363
rect 55959 -8379 55966 -8371
rect 55908 -8413 55949 -8379
rect 55970 -8413 56021 -8379
rect 56680 -8422 56685 -8406
rect 56703 -8422 56710 -8414
rect 56714 -8422 56719 -8406
rect 57010 -8408 57051 -8374
rect 57055 -8408 57062 -8363
rect 55959 -8462 55966 -8451
rect 56140 -8456 56181 -8422
rect 56212 -8456 56253 -8422
rect 56284 -8456 56325 -8422
rect 56428 -8456 56469 -8422
rect 56500 -8456 56613 -8422
rect 56644 -8456 56685 -8422
rect 55970 -8496 56011 -8462
rect 55959 -8546 55966 -8535
rect 56537 -8539 56578 -8505
rect 55970 -8580 56011 -8546
rect 55959 -8629 55966 -8618
rect 55970 -8663 56011 -8629
rect 56202 -8689 56243 -8655
rect 56247 -8689 56254 -8644
rect 56324 -8706 56329 -8588
rect 56347 -8655 56354 -8644
rect 56358 -8655 56363 -8622
rect 56394 -8655 56399 -8622
rect 56358 -8689 56399 -8655
rect 56403 -8689 56410 -8644
rect 56358 -8740 56363 -8689
rect 56394 -8740 56399 -8689
rect 56428 -8706 56433 -8589
rect 56537 -8623 56578 -8589
rect 56537 -8706 56578 -8672
rect 56680 -8706 56685 -8456
rect 56714 -8456 56755 -8422
rect 56703 -8505 56710 -8494
rect 56714 -8505 56719 -8456
rect 57010 -8491 57051 -8457
rect 57055 -8491 57062 -8446
rect 56714 -8539 56755 -8505
rect 56703 -8589 56710 -8578
rect 56714 -8589 56719 -8539
rect 56863 -8565 56972 -8499
rect 57132 -8507 57137 -8191
rect 57155 -8207 57162 -8199
rect 57166 -8207 57171 -8191
rect 57166 -8241 57207 -8207
rect 57211 -8241 57218 -8199
rect 57155 -8290 57162 -8279
rect 57166 -8290 57171 -8241
rect 57166 -8324 57207 -8290
rect 57211 -8324 57218 -8279
rect 57155 -8374 57162 -8363
rect 57166 -8374 57171 -8324
rect 57166 -8408 57207 -8374
rect 57211 -8408 57218 -8363
rect 57155 -8457 57162 -8446
rect 57166 -8457 57171 -8408
rect 57166 -8491 57207 -8457
rect 57211 -8491 57218 -8446
rect 57155 -8525 57162 -8499
rect 57166 -8541 57171 -8491
rect 56714 -8623 56755 -8589
rect 57075 -8605 57116 -8571
rect 56703 -8672 56710 -8661
rect 56714 -8672 56719 -8623
rect 56714 -8706 56755 -8672
rect 57197 -8673 57204 -8525
rect 57220 -8541 57223 -8191
rect 57254 -8507 57257 -8191
rect 57311 -8207 57318 -8199
rect 57260 -8241 57301 -8207
rect 57322 -8241 57373 -8207
rect 58237 -8231 58278 -8197
rect 58333 -8231 58374 -8197
rect 58429 -8231 58470 -8197
rect 60399 -8207 60406 -8199
rect 58030 -8250 58035 -8234
rect 58053 -8250 58060 -8242
rect 58064 -8250 58069 -8234
rect 57311 -8290 57318 -8279
rect 57490 -8284 57531 -8250
rect 57562 -8284 57603 -8250
rect 57634 -8284 57675 -8250
rect 57778 -8284 57819 -8250
rect 57850 -8284 57963 -8250
rect 57994 -8284 58035 -8250
rect 57322 -8324 57363 -8290
rect 57311 -8374 57318 -8363
rect 57887 -8367 57928 -8333
rect 57322 -8408 57363 -8374
rect 57311 -8457 57318 -8446
rect 57322 -8491 57363 -8457
rect 57552 -8517 57593 -8483
rect 57597 -8517 57604 -8472
rect 57674 -8534 57679 -8416
rect 57697 -8483 57704 -8472
rect 57708 -8483 57713 -8450
rect 57744 -8483 57749 -8450
rect 57708 -8517 57749 -8483
rect 57753 -8517 57760 -8472
rect 57708 -8568 57713 -8517
rect 57744 -8568 57749 -8517
rect 57778 -8534 57783 -8417
rect 57887 -8451 57928 -8417
rect 57887 -8534 57928 -8500
rect 58030 -8534 58035 -8284
rect 58064 -8284 58105 -8250
rect 58591 -8274 58632 -8240
rect 58687 -8274 58728 -8240
rect 58783 -8274 58824 -8240
rect 60290 -8241 60331 -8207
rect 60354 -8241 60406 -8207
rect 60434 -8241 60475 -8207
rect 58053 -8333 58060 -8322
rect 58064 -8333 58069 -8284
rect 58303 -8293 58310 -8285
rect 58403 -8293 58410 -8285
rect 58230 -8327 58299 -8293
rect 58302 -8327 58343 -8293
rect 58414 -8327 58455 -8293
rect 58945 -8317 58986 -8283
rect 59041 -8317 59082 -8283
rect 59137 -8317 59178 -8283
rect 59233 -8317 59274 -8283
rect 59329 -8317 59370 -8283
rect 60354 -8324 60395 -8290
rect 60399 -8324 60406 -8279
rect 58064 -8367 58105 -8333
rect 58657 -8336 58664 -8328
rect 58757 -8336 58764 -8328
rect 58053 -8417 58060 -8406
rect 58064 -8417 58069 -8367
rect 58258 -8410 58299 -8376
rect 58303 -8410 58310 -8365
rect 58403 -8376 58410 -8365
rect 58584 -8370 58653 -8336
rect 58656 -8370 58697 -8336
rect 58768 -8370 58809 -8336
rect 59493 -8360 59534 -8326
rect 59589 -8360 59630 -8326
rect 59685 -8360 59726 -8326
rect 59781 -8360 59822 -8326
rect 59877 -8360 59918 -8326
rect 59973 -8360 60014 -8326
rect 60069 -8360 60110 -8326
rect 58414 -8410 58455 -8376
rect 59047 -8379 59054 -8371
rect 58064 -8451 58105 -8417
rect 58053 -8500 58060 -8489
rect 58064 -8500 58069 -8451
rect 58258 -8494 58299 -8460
rect 58303 -8494 58310 -8449
rect 58403 -8460 58410 -8449
rect 58612 -8453 58653 -8419
rect 58657 -8453 58664 -8408
rect 58757 -8419 58764 -8408
rect 58938 -8413 58979 -8379
rect 59002 -8413 59054 -8379
rect 59082 -8413 59123 -8379
rect 58768 -8453 58809 -8419
rect 58414 -8494 58455 -8460
rect 58064 -8534 58105 -8500
rect 58064 -8568 58069 -8534
rect 56714 -8740 56719 -8706
rect 57010 -8723 57051 -8689
rect 57055 -8723 57062 -8681
rect 57197 -8741 57209 -8673
rect 57238 -8707 57243 -8639
rect 57283 -8671 57288 -8603
rect 57317 -8637 57322 -8571
rect 58258 -8577 58299 -8543
rect 58303 -8577 58310 -8532
rect 58403 -8543 58410 -8532
rect 58612 -8537 58653 -8503
rect 58657 -8537 58664 -8492
rect 58757 -8503 58764 -8492
rect 59002 -8496 59043 -8462
rect 59047 -8496 59054 -8451
rect 58768 -8537 58809 -8503
rect 58414 -8577 58455 -8543
rect 57327 -8621 57368 -8587
rect 57528 -8666 57569 -8632
rect 57297 -8689 57304 -8681
rect 57308 -8723 57349 -8689
rect 57528 -8734 57569 -8700
rect 54461 -8906 54502 -8872
rect 54533 -8906 54574 -8872
rect 54605 -8906 54646 -8872
rect 54918 -8913 54959 -8879
rect 54963 -8913 54970 -8868
rect 55063 -8879 55070 -8868
rect 55074 -8913 55115 -8879
rect 55658 -8895 55699 -8861
rect 55703 -8895 55710 -8853
rect 53552 -8959 54034 -8925
rect 54886 -8949 54927 -8915
rect 54958 -8949 54999 -8915
rect 55272 -8956 55313 -8922
rect 55317 -8956 55324 -8911
rect 55417 -8922 55424 -8911
rect 55845 -8913 55857 -8845
rect 55886 -8879 55891 -8811
rect 55931 -8843 55936 -8775
rect 55965 -8809 55970 -8743
rect 57197 -8753 57204 -8741
rect 57577 -8750 57582 -8616
rect 55975 -8793 56016 -8759
rect 56178 -8838 56219 -8804
rect 55945 -8861 55952 -8853
rect 55956 -8895 55997 -8861
rect 56178 -8906 56219 -8872
rect 55428 -8956 55469 -8922
rect 53552 -8985 54021 -8959
rect 53555 -8993 53763 -8985
rect 53571 -9003 53747 -8993
rect 53297 -9140 53479 -9114
rect 52804 -9174 52846 -9140
rect 52900 -9174 52942 -9140
rect 52996 -9174 53038 -9140
rect 53092 -9174 53134 -9140
rect 53188 -9174 53230 -9140
rect 53284 -9174 53479 -9140
rect 53297 -9200 53479 -9174
rect 53497 -9174 53605 -9050
rect 53756 -9062 53763 -9051
rect 53375 -9870 53417 -9200
rect 53497 -9228 53507 -9174
rect 53182 -9936 53334 -9924
rect 52850 -9970 53334 -9936
rect 53182 -9971 53334 -9970
rect 53363 -9971 53417 -9870
rect 53509 -9971 53551 -9174
rect 53555 -9971 53562 -9174
rect 53767 -9971 53809 -9062
rect 53901 -9971 53943 -8985
rect 54155 -9002 54196 -8968
rect 54251 -9002 54292 -8968
rect 54347 -9002 54388 -8968
rect 54443 -9002 54484 -8968
rect 54539 -9002 54580 -8968
rect 54635 -9002 54676 -8968
rect 54731 -9002 54772 -8968
rect 55240 -8992 55281 -8958
rect 55312 -8992 55353 -8958
rect 55658 -8995 55699 -8961
rect 55703 -8995 55710 -8950
rect 55845 -9001 55852 -8913
rect 56227 -8922 56232 -8788
rect 55945 -8961 55952 -8950
rect 56261 -8956 56266 -8762
rect 56301 -8778 56308 -8767
rect 56297 -8809 56308 -8778
rect 56623 -8796 56664 -8762
rect 55956 -8995 55997 -8961
rect 54893 -9045 54934 -9011
rect 54989 -9045 55030 -9011
rect 55085 -9045 55126 -9011
rect 55594 -9035 55635 -9001
rect 55666 -9035 55707 -9001
rect 55738 -9035 55779 -9001
rect 55810 -9029 55852 -9001
rect 56156 -9025 56197 -8991
rect 56201 -9025 56208 -8980
rect 56297 -8992 56302 -8809
rect 56331 -8995 56336 -8812
rect 55810 -9035 55851 -9029
rect 55247 -9088 55288 -9054
rect 55343 -9088 55384 -9054
rect 55439 -9088 55480 -9054
rect 56343 -9076 56350 -8809
rect 56972 -8819 57365 -8753
rect 57611 -8784 57616 -8590
rect 57651 -8606 57658 -8595
rect 57647 -8637 57658 -8606
rect 57973 -8624 58014 -8590
rect 56359 -8860 56400 -8826
rect 56708 -8830 56725 -8819
rect 56708 -8832 56714 -8830
rect 56359 -8928 56400 -8894
rect 56411 -8995 56416 -8860
rect 56642 -8874 56714 -8832
rect 56770 -8874 57365 -8819
rect 57506 -8853 57547 -8819
rect 57551 -8853 57558 -8808
rect 57647 -8820 57652 -8637
rect 57681 -8823 57686 -8640
rect 56642 -8877 57365 -8874
rect 56445 -8980 56450 -8892
rect 56562 -8942 56603 -8908
rect 56607 -8942 56614 -8900
rect 56443 -8991 56450 -8980
rect 56445 -9025 56450 -8991
rect 56454 -9025 56495 -8991
rect 56562 -9042 56603 -9008
rect 56607 -9042 56614 -8997
rect 56455 -9078 56496 -9044
rect 56527 -9078 56568 -9044
rect 56599 -9078 56640 -9044
rect 55601 -9131 55642 -9097
rect 55697 -9131 55738 -9097
rect 55793 -9131 55834 -9097
rect 55889 -9131 55930 -9097
rect 55985 -9131 56026 -9097
rect 56642 -9114 56793 -8877
rect 56972 -8899 57365 -8877
rect 56896 -8925 57365 -8899
rect 57693 -8904 57700 -8637
rect 57709 -8688 57750 -8654
rect 57709 -8756 57750 -8722
rect 57761 -8823 57766 -8688
rect 58323 -8691 58364 -8657
rect 58375 -8718 58380 -8641
rect 57795 -8808 57800 -8720
rect 57912 -8770 57953 -8736
rect 57957 -8770 57964 -8728
rect 58057 -8740 58064 -8729
rect 58068 -8774 58109 -8740
rect 58409 -8752 58414 -8607
rect 58612 -8620 58653 -8586
rect 58657 -8620 58664 -8575
rect 58757 -8586 58764 -8575
rect 59002 -8580 59043 -8546
rect 59047 -8580 59054 -8535
rect 58768 -8620 58809 -8586
rect 58677 -8734 58718 -8700
rect 58729 -8761 58734 -8684
rect 57793 -8819 57800 -8808
rect 58262 -8813 58303 -8779
rect 58307 -8813 58314 -8771
rect 58407 -8779 58414 -8771
rect 58418 -8813 58459 -8779
rect 58763 -8795 58768 -8650
rect 59002 -8663 59043 -8629
rect 59047 -8663 59054 -8618
rect 59124 -8679 59129 -8363
rect 59147 -8379 59154 -8371
rect 59158 -8379 59163 -8363
rect 59158 -8413 59199 -8379
rect 59203 -8413 59210 -8371
rect 59147 -8462 59154 -8451
rect 59158 -8462 59163 -8413
rect 59158 -8496 59199 -8462
rect 59203 -8496 59210 -8451
rect 59147 -8546 59154 -8535
rect 59158 -8546 59163 -8496
rect 59158 -8580 59199 -8546
rect 59203 -8580 59210 -8535
rect 59147 -8629 59154 -8618
rect 59158 -8629 59163 -8580
rect 59158 -8663 59199 -8629
rect 59203 -8663 59210 -8618
rect 59147 -8697 59154 -8671
rect 59158 -8713 59163 -8663
rect 59067 -8777 59108 -8743
rect 57795 -8853 57800 -8819
rect 57804 -8853 57845 -8819
rect 57912 -8870 57953 -8836
rect 57957 -8870 57964 -8825
rect 58057 -8832 58064 -8821
rect 58068 -8866 58109 -8832
rect 58616 -8856 58657 -8822
rect 58661 -8856 58668 -8814
rect 58761 -8822 58768 -8814
rect 58772 -8856 58813 -8822
rect 59189 -8845 59196 -8697
rect 59212 -8713 59215 -8363
rect 59246 -8679 59249 -8363
rect 59303 -8379 59310 -8371
rect 59252 -8413 59293 -8379
rect 59314 -8413 59365 -8379
rect 60024 -8422 60029 -8406
rect 60047 -8422 60054 -8414
rect 60058 -8422 60063 -8406
rect 60354 -8408 60395 -8374
rect 60399 -8408 60406 -8363
rect 59303 -8462 59310 -8451
rect 59484 -8456 59525 -8422
rect 59556 -8456 59597 -8422
rect 59628 -8456 59669 -8422
rect 59772 -8456 59813 -8422
rect 59844 -8456 59957 -8422
rect 59988 -8456 60029 -8422
rect 59314 -8496 59355 -8462
rect 59303 -8546 59310 -8535
rect 59881 -8539 59922 -8505
rect 59314 -8580 59355 -8546
rect 59303 -8629 59310 -8618
rect 59314 -8663 59355 -8629
rect 59546 -8689 59587 -8655
rect 59591 -8689 59598 -8644
rect 59668 -8706 59673 -8588
rect 59691 -8655 59698 -8644
rect 59702 -8655 59707 -8622
rect 59738 -8655 59743 -8622
rect 59702 -8689 59743 -8655
rect 59747 -8689 59754 -8644
rect 59702 -8740 59707 -8689
rect 59738 -8740 59743 -8689
rect 59772 -8706 59777 -8589
rect 59881 -8623 59922 -8589
rect 59881 -8706 59922 -8672
rect 60024 -8706 60029 -8456
rect 60058 -8456 60099 -8422
rect 60047 -8505 60054 -8494
rect 60058 -8505 60063 -8456
rect 60354 -8491 60395 -8457
rect 60399 -8491 60406 -8446
rect 60058 -8539 60099 -8505
rect 60047 -8589 60054 -8578
rect 60058 -8589 60063 -8539
rect 60207 -8565 60316 -8499
rect 60476 -8507 60481 -8191
rect 60499 -8207 60506 -8199
rect 60510 -8207 60515 -8191
rect 60510 -8241 60551 -8207
rect 60555 -8241 60562 -8199
rect 60499 -8290 60506 -8279
rect 60510 -8290 60515 -8241
rect 60510 -8324 60551 -8290
rect 60555 -8324 60562 -8279
rect 60499 -8374 60506 -8363
rect 60510 -8374 60515 -8324
rect 60510 -8408 60551 -8374
rect 60555 -8408 60562 -8363
rect 60499 -8457 60506 -8446
rect 60510 -8457 60515 -8408
rect 60510 -8491 60551 -8457
rect 60555 -8491 60562 -8446
rect 60499 -8525 60506 -8499
rect 60510 -8541 60515 -8491
rect 60058 -8623 60099 -8589
rect 60419 -8605 60460 -8571
rect 60047 -8672 60054 -8661
rect 60058 -8672 60063 -8623
rect 60058 -8706 60099 -8672
rect 60541 -8673 60548 -8525
rect 60564 -8541 60567 -8191
rect 60598 -8507 60601 -8191
rect 60655 -8207 60662 -8199
rect 60604 -8241 60645 -8207
rect 60666 -8241 60717 -8207
rect 61581 -8231 61622 -8197
rect 61677 -8231 61718 -8197
rect 61773 -8231 61814 -8197
rect 63743 -8207 63750 -8199
rect 61374 -8250 61379 -8234
rect 61397 -8250 61404 -8242
rect 61408 -8250 61413 -8234
rect 60655 -8290 60662 -8279
rect 60834 -8284 60875 -8250
rect 60906 -8284 60947 -8250
rect 60978 -8284 61019 -8250
rect 61122 -8284 61163 -8250
rect 61194 -8284 61307 -8250
rect 61338 -8284 61379 -8250
rect 60666 -8324 60707 -8290
rect 60655 -8374 60662 -8363
rect 61231 -8367 61272 -8333
rect 60666 -8408 60707 -8374
rect 60655 -8457 60662 -8446
rect 60666 -8491 60707 -8457
rect 60896 -8517 60937 -8483
rect 60941 -8517 60948 -8472
rect 61018 -8534 61023 -8416
rect 61041 -8483 61048 -8472
rect 61052 -8483 61057 -8450
rect 61088 -8483 61093 -8450
rect 61052 -8517 61093 -8483
rect 61097 -8517 61104 -8472
rect 61052 -8568 61057 -8517
rect 61088 -8568 61093 -8517
rect 61122 -8534 61127 -8417
rect 61231 -8451 61272 -8417
rect 61231 -8534 61272 -8500
rect 61374 -8534 61379 -8284
rect 61408 -8284 61449 -8250
rect 61935 -8274 61976 -8240
rect 62031 -8274 62072 -8240
rect 62127 -8274 62168 -8240
rect 63634 -8241 63675 -8207
rect 63698 -8241 63750 -8207
rect 63778 -8241 63819 -8207
rect 61397 -8333 61404 -8322
rect 61408 -8333 61413 -8284
rect 61647 -8293 61654 -8285
rect 61747 -8293 61754 -8285
rect 61574 -8327 61643 -8293
rect 61646 -8327 61687 -8293
rect 61758 -8327 61799 -8293
rect 62289 -8317 62330 -8283
rect 62385 -8317 62426 -8283
rect 62481 -8317 62522 -8283
rect 62577 -8317 62618 -8283
rect 62673 -8317 62714 -8283
rect 63698 -8324 63739 -8290
rect 63743 -8324 63750 -8279
rect 61408 -8367 61449 -8333
rect 62001 -8336 62008 -8328
rect 62101 -8336 62108 -8328
rect 61397 -8417 61404 -8406
rect 61408 -8417 61413 -8367
rect 61602 -8410 61643 -8376
rect 61647 -8410 61654 -8365
rect 61747 -8376 61754 -8365
rect 61928 -8370 61997 -8336
rect 62000 -8370 62041 -8336
rect 62112 -8370 62153 -8336
rect 62837 -8360 62878 -8326
rect 62933 -8360 62974 -8326
rect 63029 -8360 63070 -8326
rect 63125 -8360 63166 -8326
rect 63221 -8360 63262 -8326
rect 63317 -8360 63358 -8326
rect 63413 -8360 63454 -8326
rect 61758 -8410 61799 -8376
rect 62391 -8379 62398 -8371
rect 61408 -8451 61449 -8417
rect 61397 -8500 61404 -8489
rect 61408 -8500 61413 -8451
rect 61602 -8494 61643 -8460
rect 61647 -8494 61654 -8449
rect 61747 -8460 61754 -8449
rect 61956 -8453 61997 -8419
rect 62001 -8453 62008 -8408
rect 62101 -8419 62108 -8408
rect 62282 -8413 62323 -8379
rect 62346 -8413 62398 -8379
rect 62426 -8413 62467 -8379
rect 62112 -8453 62153 -8419
rect 61758 -8494 61799 -8460
rect 61408 -8534 61449 -8500
rect 61408 -8568 61413 -8534
rect 60058 -8740 60063 -8706
rect 60354 -8723 60395 -8689
rect 60399 -8723 60406 -8681
rect 60541 -8741 60553 -8673
rect 60582 -8707 60587 -8639
rect 60627 -8671 60632 -8603
rect 60661 -8637 60666 -8571
rect 61602 -8577 61643 -8543
rect 61647 -8577 61654 -8532
rect 61747 -8543 61754 -8532
rect 61956 -8537 61997 -8503
rect 62001 -8537 62008 -8492
rect 62101 -8503 62108 -8492
rect 62346 -8496 62387 -8462
rect 62391 -8496 62398 -8451
rect 62112 -8537 62153 -8503
rect 61758 -8577 61799 -8543
rect 60671 -8621 60712 -8587
rect 60872 -8666 60913 -8632
rect 60641 -8689 60648 -8681
rect 60652 -8723 60693 -8689
rect 60872 -8734 60913 -8700
rect 57805 -8906 57846 -8872
rect 57877 -8906 57918 -8872
rect 57949 -8906 57990 -8872
rect 58262 -8913 58303 -8879
rect 58307 -8913 58314 -8868
rect 58407 -8879 58414 -8868
rect 58418 -8913 58459 -8879
rect 59002 -8895 59043 -8861
rect 59047 -8895 59054 -8853
rect 56896 -8959 57378 -8925
rect 58230 -8949 58271 -8915
rect 58302 -8949 58343 -8915
rect 58616 -8956 58657 -8922
rect 58661 -8956 58668 -8911
rect 58761 -8922 58768 -8911
rect 59189 -8913 59201 -8845
rect 59230 -8879 59235 -8811
rect 59275 -8843 59280 -8775
rect 59309 -8809 59314 -8743
rect 60541 -8753 60548 -8741
rect 60921 -8750 60926 -8616
rect 59319 -8793 59360 -8759
rect 59522 -8838 59563 -8804
rect 59289 -8861 59296 -8853
rect 59300 -8895 59341 -8861
rect 59522 -8906 59563 -8872
rect 58772 -8956 58813 -8922
rect 56896 -8985 57365 -8959
rect 56900 -8993 57107 -8985
rect 56916 -9003 57091 -8993
rect 56642 -9140 56823 -9114
rect 56149 -9174 56190 -9140
rect 56245 -9174 56286 -9140
rect 56341 -9174 56382 -9140
rect 56437 -9174 56478 -9140
rect 56533 -9174 56574 -9140
rect 56629 -9174 56823 -9140
rect 56642 -9200 56823 -9174
rect 56842 -9174 56949 -9050
rect 57101 -9062 57107 -9051
rect 56720 -9870 56761 -9200
rect 56842 -9228 56851 -9174
rect 56527 -9936 56678 -9924
rect 56195 -9970 56678 -9936
rect 56527 -9971 56678 -9970
rect 56708 -9971 56761 -9870
rect 56854 -9971 56895 -9174
rect 56900 -9971 56906 -9174
rect 57112 -9971 57153 -9062
rect 57246 -9971 57287 -8985
rect 57499 -9002 57540 -8968
rect 57595 -9002 57636 -8968
rect 57691 -9002 57732 -8968
rect 57787 -9002 57828 -8968
rect 57883 -9002 57924 -8968
rect 57979 -9002 58020 -8968
rect 58075 -9002 58116 -8968
rect 58584 -8992 58625 -8958
rect 58656 -8992 58697 -8958
rect 59002 -8995 59043 -8961
rect 59047 -8995 59054 -8950
rect 59189 -9001 59196 -8913
rect 59571 -8922 59576 -8788
rect 59289 -8961 59296 -8950
rect 59605 -8956 59610 -8762
rect 59645 -8778 59652 -8767
rect 59641 -8809 59652 -8778
rect 59967 -8796 60008 -8762
rect 59300 -8995 59341 -8961
rect 58237 -9045 58278 -9011
rect 58333 -9045 58374 -9011
rect 58429 -9045 58470 -9011
rect 58938 -9035 58979 -9001
rect 59010 -9035 59051 -9001
rect 59082 -9035 59123 -9001
rect 59154 -9029 59196 -9001
rect 59500 -9025 59541 -8991
rect 59545 -9025 59552 -8980
rect 59641 -8992 59646 -8809
rect 59675 -8995 59680 -8812
rect 59154 -9035 59195 -9029
rect 58591 -9088 58632 -9054
rect 58687 -9088 58728 -9054
rect 58783 -9088 58824 -9054
rect 59687 -9076 59694 -8809
rect 60316 -8819 60709 -8753
rect 60955 -8784 60960 -8590
rect 60995 -8606 61002 -8595
rect 60991 -8637 61002 -8606
rect 61317 -8624 61358 -8590
rect 59703 -8860 59744 -8826
rect 60052 -8830 60069 -8819
rect 60052 -8832 60058 -8830
rect 59703 -8928 59744 -8894
rect 59755 -8995 59760 -8860
rect 59986 -8874 60058 -8832
rect 60114 -8874 60709 -8819
rect 60850 -8853 60891 -8819
rect 60895 -8853 60902 -8808
rect 60991 -8820 60996 -8637
rect 61025 -8823 61030 -8640
rect 59986 -8877 60709 -8874
rect 59789 -8980 59794 -8892
rect 59906 -8942 59947 -8908
rect 59951 -8942 59958 -8900
rect 59787 -8991 59794 -8980
rect 59789 -9025 59794 -8991
rect 59798 -9025 59839 -8991
rect 59906 -9042 59947 -9008
rect 59951 -9042 59958 -8997
rect 59799 -9078 59840 -9044
rect 59871 -9078 59912 -9044
rect 59943 -9078 59984 -9044
rect 58945 -9131 58986 -9097
rect 59041 -9131 59082 -9097
rect 59137 -9131 59178 -9097
rect 59233 -9131 59274 -9097
rect 59329 -9131 59370 -9097
rect 59986 -9114 60137 -8877
rect 60316 -8899 60709 -8877
rect 60240 -8925 60709 -8899
rect 61037 -8904 61044 -8637
rect 61053 -8688 61094 -8654
rect 61053 -8756 61094 -8722
rect 61105 -8823 61110 -8688
rect 61667 -8691 61708 -8657
rect 61719 -8718 61724 -8641
rect 61139 -8808 61144 -8720
rect 61256 -8770 61297 -8736
rect 61301 -8770 61308 -8728
rect 61401 -8740 61408 -8729
rect 61412 -8774 61453 -8740
rect 61753 -8752 61758 -8607
rect 61956 -8620 61997 -8586
rect 62001 -8620 62008 -8575
rect 62101 -8586 62108 -8575
rect 62346 -8580 62387 -8546
rect 62391 -8580 62398 -8535
rect 62112 -8620 62153 -8586
rect 62021 -8734 62062 -8700
rect 62073 -8761 62078 -8684
rect 61137 -8819 61144 -8808
rect 61606 -8813 61647 -8779
rect 61651 -8813 61658 -8771
rect 61751 -8779 61758 -8771
rect 61762 -8813 61803 -8779
rect 62107 -8795 62112 -8650
rect 62346 -8663 62387 -8629
rect 62391 -8663 62398 -8618
rect 62468 -8679 62473 -8363
rect 62491 -8379 62498 -8371
rect 62502 -8379 62507 -8363
rect 62502 -8413 62543 -8379
rect 62547 -8413 62554 -8371
rect 62491 -8462 62498 -8451
rect 62502 -8462 62507 -8413
rect 62502 -8496 62543 -8462
rect 62547 -8496 62554 -8451
rect 62491 -8546 62498 -8535
rect 62502 -8546 62507 -8496
rect 62502 -8580 62543 -8546
rect 62547 -8580 62554 -8535
rect 62491 -8629 62498 -8618
rect 62502 -8629 62507 -8580
rect 62502 -8663 62543 -8629
rect 62547 -8663 62554 -8618
rect 62491 -8697 62498 -8671
rect 62502 -8713 62507 -8663
rect 62411 -8777 62452 -8743
rect 61139 -8853 61144 -8819
rect 61148 -8853 61189 -8819
rect 61256 -8870 61297 -8836
rect 61301 -8870 61308 -8825
rect 61401 -8832 61408 -8821
rect 61412 -8866 61453 -8832
rect 61960 -8856 62001 -8822
rect 62005 -8856 62012 -8814
rect 62105 -8822 62112 -8814
rect 62116 -8856 62157 -8822
rect 62533 -8845 62540 -8697
rect 62556 -8713 62559 -8363
rect 62590 -8679 62593 -8363
rect 62647 -8379 62654 -8371
rect 62596 -8413 62637 -8379
rect 62658 -8413 62709 -8379
rect 63368 -8422 63373 -8406
rect 63391 -8422 63398 -8414
rect 63402 -8422 63407 -8406
rect 63698 -8408 63739 -8374
rect 63743 -8408 63750 -8363
rect 62647 -8462 62654 -8451
rect 62828 -8456 62869 -8422
rect 62900 -8456 62941 -8422
rect 62972 -8456 63013 -8422
rect 63116 -8456 63157 -8422
rect 63188 -8456 63301 -8422
rect 63332 -8456 63373 -8422
rect 62658 -8496 62699 -8462
rect 62647 -8546 62654 -8535
rect 63225 -8539 63266 -8505
rect 62658 -8580 62699 -8546
rect 62647 -8629 62654 -8618
rect 62658 -8663 62699 -8629
rect 62890 -8689 62931 -8655
rect 62935 -8689 62942 -8644
rect 63012 -8706 63017 -8588
rect 63035 -8655 63042 -8644
rect 63046 -8655 63051 -8622
rect 63082 -8655 63087 -8622
rect 63046 -8689 63087 -8655
rect 63091 -8689 63098 -8644
rect 63046 -8740 63051 -8689
rect 63082 -8740 63087 -8689
rect 63116 -8706 63121 -8589
rect 63225 -8623 63266 -8589
rect 63225 -8706 63266 -8672
rect 63368 -8706 63373 -8456
rect 63402 -8456 63443 -8422
rect 63391 -8505 63398 -8494
rect 63402 -8505 63407 -8456
rect 63698 -8491 63739 -8457
rect 63743 -8491 63750 -8446
rect 63402 -8539 63443 -8505
rect 63391 -8589 63398 -8578
rect 63402 -8589 63407 -8539
rect 63551 -8565 63660 -8499
rect 63820 -8507 63825 -8191
rect 63843 -8207 63850 -8199
rect 63854 -8207 63859 -8191
rect 63854 -8241 63895 -8207
rect 63899 -8241 63906 -8199
rect 63843 -8290 63850 -8279
rect 63854 -8290 63859 -8241
rect 63854 -8324 63895 -8290
rect 63899 -8324 63906 -8279
rect 63843 -8374 63850 -8363
rect 63854 -8374 63859 -8324
rect 63854 -8408 63895 -8374
rect 63899 -8408 63906 -8363
rect 63843 -8457 63850 -8446
rect 63854 -8457 63859 -8408
rect 63854 -8491 63895 -8457
rect 63899 -8491 63906 -8446
rect 63843 -8525 63850 -8499
rect 63854 -8541 63859 -8491
rect 63402 -8623 63443 -8589
rect 63763 -8605 63804 -8571
rect 63391 -8672 63398 -8661
rect 63402 -8672 63407 -8623
rect 63402 -8706 63443 -8672
rect 63885 -8673 63892 -8525
rect 63908 -8541 63911 -8191
rect 63942 -8507 63945 -8191
rect 63999 -8207 64006 -8199
rect 63948 -8241 63989 -8207
rect 64010 -8241 64061 -8207
rect 64925 -8231 64966 -8197
rect 65021 -8231 65062 -8197
rect 65117 -8231 65158 -8197
rect 67087 -8207 67094 -8199
rect 64718 -8250 64723 -8234
rect 64741 -8250 64748 -8242
rect 64752 -8250 64757 -8234
rect 63999 -8290 64006 -8279
rect 64178 -8284 64219 -8250
rect 64250 -8284 64291 -8250
rect 64322 -8284 64363 -8250
rect 64466 -8284 64507 -8250
rect 64538 -8284 64651 -8250
rect 64682 -8284 64723 -8250
rect 64010 -8324 64051 -8290
rect 63999 -8374 64006 -8363
rect 64575 -8367 64616 -8333
rect 64010 -8408 64051 -8374
rect 63999 -8457 64006 -8446
rect 64010 -8491 64051 -8457
rect 64240 -8517 64281 -8483
rect 64285 -8517 64292 -8472
rect 64362 -8534 64367 -8416
rect 64385 -8483 64392 -8472
rect 64396 -8483 64401 -8450
rect 64432 -8483 64437 -8450
rect 64396 -8517 64437 -8483
rect 64441 -8517 64448 -8472
rect 64396 -8568 64401 -8517
rect 64432 -8568 64437 -8517
rect 64466 -8534 64471 -8417
rect 64575 -8451 64616 -8417
rect 64575 -8534 64616 -8500
rect 64718 -8534 64723 -8284
rect 64752 -8284 64793 -8250
rect 65279 -8274 65320 -8240
rect 65375 -8274 65416 -8240
rect 65471 -8274 65512 -8240
rect 66978 -8241 67019 -8207
rect 67042 -8241 67094 -8207
rect 67122 -8241 67163 -8207
rect 64741 -8333 64748 -8322
rect 64752 -8333 64757 -8284
rect 64991 -8293 64998 -8285
rect 65091 -8293 65098 -8285
rect 64918 -8327 64987 -8293
rect 64990 -8327 65031 -8293
rect 65102 -8327 65143 -8293
rect 65633 -8317 65674 -8283
rect 65729 -8317 65770 -8283
rect 65825 -8317 65866 -8283
rect 65921 -8317 65962 -8283
rect 66017 -8317 66058 -8283
rect 67042 -8324 67083 -8290
rect 67087 -8324 67094 -8279
rect 64752 -8367 64793 -8333
rect 65345 -8336 65352 -8328
rect 65445 -8336 65452 -8328
rect 64741 -8417 64748 -8406
rect 64752 -8417 64757 -8367
rect 64946 -8410 64987 -8376
rect 64991 -8410 64998 -8365
rect 65091 -8376 65098 -8365
rect 65272 -8370 65341 -8336
rect 65344 -8370 65385 -8336
rect 65456 -8370 65497 -8336
rect 66181 -8360 66222 -8326
rect 66277 -8360 66318 -8326
rect 66373 -8360 66414 -8326
rect 66469 -8360 66510 -8326
rect 66565 -8360 66606 -8326
rect 66661 -8360 66702 -8326
rect 66757 -8360 66798 -8326
rect 65102 -8410 65143 -8376
rect 65735 -8379 65742 -8371
rect 64752 -8451 64793 -8417
rect 64741 -8500 64748 -8489
rect 64752 -8500 64757 -8451
rect 64946 -8494 64987 -8460
rect 64991 -8494 64998 -8449
rect 65091 -8460 65098 -8449
rect 65300 -8453 65341 -8419
rect 65345 -8453 65352 -8408
rect 65445 -8419 65452 -8408
rect 65626 -8413 65667 -8379
rect 65690 -8413 65742 -8379
rect 65770 -8413 65811 -8379
rect 65456 -8453 65497 -8419
rect 65102 -8494 65143 -8460
rect 64752 -8534 64793 -8500
rect 64752 -8568 64757 -8534
rect 63402 -8740 63407 -8706
rect 63698 -8723 63739 -8689
rect 63743 -8723 63750 -8681
rect 63885 -8741 63897 -8673
rect 63926 -8707 63931 -8639
rect 63971 -8671 63976 -8603
rect 64005 -8637 64010 -8571
rect 64946 -8577 64987 -8543
rect 64991 -8577 64998 -8532
rect 65091 -8543 65098 -8532
rect 65300 -8537 65341 -8503
rect 65345 -8537 65352 -8492
rect 65445 -8503 65452 -8492
rect 65690 -8496 65731 -8462
rect 65735 -8496 65742 -8451
rect 65456 -8537 65497 -8503
rect 65102 -8577 65143 -8543
rect 64015 -8621 64056 -8587
rect 64216 -8666 64257 -8632
rect 63985 -8689 63992 -8681
rect 63996 -8723 64037 -8689
rect 64216 -8734 64257 -8700
rect 61149 -8906 61190 -8872
rect 61221 -8906 61262 -8872
rect 61293 -8906 61334 -8872
rect 61606 -8913 61647 -8879
rect 61651 -8913 61658 -8868
rect 61751 -8879 61758 -8868
rect 61762 -8913 61803 -8879
rect 62346 -8895 62387 -8861
rect 62391 -8895 62398 -8853
rect 60240 -8959 60722 -8925
rect 61574 -8949 61615 -8915
rect 61646 -8949 61687 -8915
rect 61960 -8956 62001 -8922
rect 62005 -8956 62012 -8911
rect 62105 -8922 62112 -8911
rect 62533 -8913 62545 -8845
rect 62574 -8879 62579 -8811
rect 62619 -8843 62624 -8775
rect 62653 -8809 62658 -8743
rect 63885 -8753 63892 -8741
rect 64265 -8750 64270 -8616
rect 62663 -8793 62704 -8759
rect 62866 -8838 62907 -8804
rect 62633 -8861 62640 -8853
rect 62644 -8895 62685 -8861
rect 62866 -8906 62907 -8872
rect 62116 -8956 62157 -8922
rect 60240 -8985 60709 -8959
rect 60244 -8993 60451 -8985
rect 60260 -9003 60435 -8993
rect 59986 -9140 60167 -9114
rect 59493 -9174 59534 -9140
rect 59589 -9174 59630 -9140
rect 59685 -9174 59726 -9140
rect 59781 -9174 59822 -9140
rect 59877 -9174 59918 -9140
rect 59973 -9174 60167 -9140
rect 59986 -9200 60167 -9174
rect 60186 -9174 60293 -9050
rect 60445 -9062 60451 -9051
rect 60064 -9870 60105 -9200
rect 60186 -9228 60195 -9174
rect 59871 -9936 60022 -9924
rect 59539 -9970 60022 -9936
rect 59871 -9971 60022 -9970
rect 60052 -9971 60105 -9870
rect 60198 -9971 60239 -9174
rect 60244 -9971 60250 -9174
rect 60456 -9971 60497 -9062
rect 60590 -9971 60631 -8985
rect 60843 -9002 60884 -8968
rect 60939 -9002 60980 -8968
rect 61035 -9002 61076 -8968
rect 61131 -9002 61172 -8968
rect 61227 -9002 61268 -8968
rect 61323 -9002 61364 -8968
rect 61419 -9002 61460 -8968
rect 61928 -8992 61969 -8958
rect 62000 -8992 62041 -8958
rect 62346 -8995 62387 -8961
rect 62391 -8995 62398 -8950
rect 62533 -9001 62540 -8913
rect 62915 -8922 62920 -8788
rect 62633 -8961 62640 -8950
rect 62949 -8956 62954 -8762
rect 62989 -8778 62996 -8767
rect 62985 -8809 62996 -8778
rect 63311 -8796 63352 -8762
rect 62644 -8995 62685 -8961
rect 61581 -9045 61622 -9011
rect 61677 -9045 61718 -9011
rect 61773 -9045 61814 -9011
rect 62282 -9035 62323 -9001
rect 62354 -9035 62395 -9001
rect 62426 -9035 62467 -9001
rect 62498 -9029 62540 -9001
rect 62844 -9025 62885 -8991
rect 62889 -9025 62896 -8980
rect 62985 -8992 62990 -8809
rect 63019 -8995 63024 -8812
rect 62498 -9035 62539 -9029
rect 61935 -9088 61976 -9054
rect 62031 -9088 62072 -9054
rect 62127 -9088 62168 -9054
rect 63031 -9076 63038 -8809
rect 63660 -8819 64053 -8753
rect 64299 -8784 64304 -8590
rect 64339 -8606 64346 -8595
rect 64335 -8637 64346 -8606
rect 64661 -8624 64702 -8590
rect 63047 -8860 63088 -8826
rect 63396 -8830 63413 -8819
rect 63396 -8832 63402 -8830
rect 63047 -8928 63088 -8894
rect 63099 -8995 63104 -8860
rect 63330 -8874 63402 -8832
rect 63458 -8874 64053 -8819
rect 64194 -8853 64235 -8819
rect 64239 -8853 64246 -8808
rect 64335 -8820 64340 -8637
rect 64369 -8823 64374 -8640
rect 63330 -8877 64053 -8874
rect 63133 -8980 63138 -8892
rect 63250 -8942 63291 -8908
rect 63295 -8942 63302 -8900
rect 63131 -8991 63138 -8980
rect 63133 -9025 63138 -8991
rect 63142 -9025 63183 -8991
rect 63250 -9042 63291 -9008
rect 63295 -9042 63302 -8997
rect 63143 -9078 63184 -9044
rect 63215 -9078 63256 -9044
rect 63287 -9078 63328 -9044
rect 62289 -9131 62330 -9097
rect 62385 -9131 62426 -9097
rect 62481 -9131 62522 -9097
rect 62577 -9131 62618 -9097
rect 62673 -9131 62714 -9097
rect 63330 -9114 63481 -8877
rect 63660 -8899 64053 -8877
rect 63584 -8925 64053 -8899
rect 64381 -8904 64388 -8637
rect 64397 -8688 64438 -8654
rect 64397 -8756 64438 -8722
rect 64449 -8823 64454 -8688
rect 65011 -8691 65052 -8657
rect 65063 -8718 65068 -8641
rect 64483 -8808 64488 -8720
rect 64600 -8770 64641 -8736
rect 64645 -8770 64652 -8728
rect 64745 -8740 64752 -8729
rect 64756 -8774 64797 -8740
rect 65097 -8752 65102 -8607
rect 65300 -8620 65341 -8586
rect 65345 -8620 65352 -8575
rect 65445 -8586 65452 -8575
rect 65690 -8580 65731 -8546
rect 65735 -8580 65742 -8535
rect 65456 -8620 65497 -8586
rect 65365 -8734 65406 -8700
rect 65417 -8761 65422 -8684
rect 64481 -8819 64488 -8808
rect 64950 -8813 64991 -8779
rect 64995 -8813 65002 -8771
rect 65095 -8779 65102 -8771
rect 65106 -8813 65147 -8779
rect 65451 -8795 65456 -8650
rect 65690 -8663 65731 -8629
rect 65735 -8663 65742 -8618
rect 65812 -8679 65817 -8363
rect 65835 -8379 65842 -8371
rect 65846 -8379 65851 -8363
rect 65846 -8413 65887 -8379
rect 65891 -8413 65898 -8371
rect 65835 -8462 65842 -8451
rect 65846 -8462 65851 -8413
rect 65846 -8496 65887 -8462
rect 65891 -8496 65898 -8451
rect 65835 -8546 65842 -8535
rect 65846 -8546 65851 -8496
rect 65846 -8580 65887 -8546
rect 65891 -8580 65898 -8535
rect 65835 -8629 65842 -8618
rect 65846 -8629 65851 -8580
rect 65846 -8663 65887 -8629
rect 65891 -8663 65898 -8618
rect 65835 -8697 65842 -8671
rect 65846 -8713 65851 -8663
rect 65755 -8777 65796 -8743
rect 64483 -8853 64488 -8819
rect 64492 -8853 64533 -8819
rect 64600 -8870 64641 -8836
rect 64645 -8870 64652 -8825
rect 64745 -8832 64752 -8821
rect 64756 -8866 64797 -8832
rect 65304 -8856 65345 -8822
rect 65349 -8856 65356 -8814
rect 65449 -8822 65456 -8814
rect 65460 -8856 65501 -8822
rect 65877 -8845 65884 -8697
rect 65900 -8713 65903 -8363
rect 65934 -8679 65937 -8363
rect 65991 -8379 65998 -8371
rect 65940 -8413 65981 -8379
rect 66002 -8413 66053 -8379
rect 66712 -8422 66717 -8406
rect 66735 -8422 66742 -8414
rect 66746 -8422 66751 -8406
rect 67042 -8408 67083 -8374
rect 67087 -8408 67094 -8363
rect 65991 -8462 65998 -8451
rect 66172 -8456 66213 -8422
rect 66244 -8456 66285 -8422
rect 66316 -8456 66357 -8422
rect 66460 -8456 66501 -8422
rect 66532 -8456 66645 -8422
rect 66676 -8456 66717 -8422
rect 66002 -8496 66043 -8462
rect 65991 -8546 65998 -8535
rect 66569 -8539 66610 -8505
rect 66002 -8580 66043 -8546
rect 65991 -8629 65998 -8618
rect 66002 -8663 66043 -8629
rect 66234 -8689 66275 -8655
rect 66279 -8689 66286 -8644
rect 66356 -8706 66361 -8588
rect 66379 -8655 66386 -8644
rect 66390 -8655 66395 -8622
rect 66426 -8655 66431 -8622
rect 66390 -8689 66431 -8655
rect 66435 -8689 66442 -8644
rect 66390 -8740 66395 -8689
rect 66426 -8740 66431 -8689
rect 66460 -8706 66465 -8589
rect 66569 -8623 66610 -8589
rect 66569 -8706 66610 -8672
rect 66712 -8706 66717 -8456
rect 66746 -8456 66787 -8422
rect 66735 -8505 66742 -8494
rect 66746 -8505 66751 -8456
rect 67042 -8491 67083 -8457
rect 67087 -8491 67094 -8446
rect 66746 -8539 66787 -8505
rect 66735 -8589 66742 -8578
rect 66746 -8589 66751 -8539
rect 66895 -8565 67004 -8499
rect 67164 -8507 67169 -8191
rect 67187 -8207 67194 -8199
rect 67198 -8207 67203 -8191
rect 67198 -8241 67239 -8207
rect 67243 -8241 67250 -8199
rect 67187 -8290 67194 -8279
rect 67198 -8290 67203 -8241
rect 67198 -8324 67239 -8290
rect 67243 -8324 67250 -8279
rect 67187 -8374 67194 -8363
rect 67198 -8374 67203 -8324
rect 67198 -8408 67239 -8374
rect 67243 -8408 67250 -8363
rect 67187 -8457 67194 -8446
rect 67198 -8457 67203 -8408
rect 67198 -8491 67239 -8457
rect 67243 -8491 67250 -8446
rect 67187 -8525 67194 -8499
rect 67198 -8541 67203 -8491
rect 66746 -8623 66787 -8589
rect 67107 -8605 67148 -8571
rect 66735 -8672 66742 -8661
rect 66746 -8672 66751 -8623
rect 66746 -8706 66787 -8672
rect 67229 -8673 67236 -8525
rect 67252 -8541 67255 -8191
rect 67286 -8507 67289 -8191
rect 67343 -8207 67350 -8199
rect 67292 -8241 67333 -8207
rect 67354 -8241 67405 -8207
rect 68269 -8231 68310 -8197
rect 68365 -8231 68406 -8197
rect 68461 -8231 68502 -8197
rect 70431 -8207 70438 -8199
rect 68062 -8250 68067 -8234
rect 68085 -8250 68092 -8242
rect 68096 -8250 68101 -8234
rect 67343 -8290 67350 -8279
rect 67522 -8284 67563 -8250
rect 67594 -8284 67635 -8250
rect 67666 -8284 67707 -8250
rect 67810 -8284 67851 -8250
rect 67882 -8284 67995 -8250
rect 68026 -8284 68067 -8250
rect 67354 -8324 67395 -8290
rect 67343 -8374 67350 -8363
rect 67919 -8367 67960 -8333
rect 67354 -8408 67395 -8374
rect 67343 -8457 67350 -8446
rect 67354 -8491 67395 -8457
rect 67584 -8517 67625 -8483
rect 67629 -8517 67636 -8472
rect 67706 -8534 67711 -8416
rect 67729 -8483 67736 -8472
rect 67740 -8483 67745 -8450
rect 67776 -8483 67781 -8450
rect 67740 -8517 67781 -8483
rect 67785 -8517 67792 -8472
rect 67740 -8568 67745 -8517
rect 67776 -8568 67781 -8517
rect 67810 -8534 67815 -8417
rect 67919 -8451 67960 -8417
rect 67919 -8534 67960 -8500
rect 68062 -8534 68067 -8284
rect 68096 -8284 68137 -8250
rect 68623 -8274 68664 -8240
rect 68719 -8274 68760 -8240
rect 68815 -8274 68856 -8240
rect 70322 -8241 70363 -8207
rect 70386 -8241 70438 -8207
rect 70466 -8241 70507 -8207
rect 68085 -8333 68092 -8322
rect 68096 -8333 68101 -8284
rect 68335 -8293 68342 -8285
rect 68435 -8293 68442 -8285
rect 68262 -8327 68331 -8293
rect 68334 -8327 68375 -8293
rect 68446 -8327 68487 -8293
rect 68977 -8317 69018 -8283
rect 69073 -8317 69114 -8283
rect 69169 -8317 69210 -8283
rect 69265 -8317 69306 -8283
rect 69361 -8317 69402 -8283
rect 70386 -8324 70427 -8290
rect 70431 -8324 70438 -8279
rect 68096 -8367 68137 -8333
rect 68689 -8336 68696 -8328
rect 68789 -8336 68796 -8328
rect 68085 -8417 68092 -8406
rect 68096 -8417 68101 -8367
rect 68290 -8410 68331 -8376
rect 68335 -8410 68342 -8365
rect 68435 -8376 68442 -8365
rect 68616 -8370 68685 -8336
rect 68688 -8370 68729 -8336
rect 68800 -8370 68841 -8336
rect 69525 -8360 69566 -8326
rect 69621 -8360 69662 -8326
rect 69717 -8360 69758 -8326
rect 69813 -8360 69854 -8326
rect 69909 -8360 69950 -8326
rect 70005 -8360 70046 -8326
rect 70101 -8360 70142 -8326
rect 68446 -8410 68487 -8376
rect 69079 -8379 69086 -8371
rect 68096 -8451 68137 -8417
rect 68085 -8500 68092 -8489
rect 68096 -8500 68101 -8451
rect 68290 -8494 68331 -8460
rect 68335 -8494 68342 -8449
rect 68435 -8460 68442 -8449
rect 68644 -8453 68685 -8419
rect 68689 -8453 68696 -8408
rect 68789 -8419 68796 -8408
rect 68970 -8413 69011 -8379
rect 69034 -8413 69086 -8379
rect 69114 -8413 69155 -8379
rect 68800 -8453 68841 -8419
rect 68446 -8494 68487 -8460
rect 68096 -8534 68137 -8500
rect 68096 -8568 68101 -8534
rect 66746 -8740 66751 -8706
rect 67042 -8723 67083 -8689
rect 67087 -8723 67094 -8681
rect 67229 -8741 67241 -8673
rect 67270 -8707 67275 -8639
rect 67315 -8671 67320 -8603
rect 67349 -8637 67354 -8571
rect 68290 -8577 68331 -8543
rect 68335 -8577 68342 -8532
rect 68435 -8543 68442 -8532
rect 68644 -8537 68685 -8503
rect 68689 -8537 68696 -8492
rect 68789 -8503 68796 -8492
rect 69034 -8496 69075 -8462
rect 69079 -8496 69086 -8451
rect 68800 -8537 68841 -8503
rect 68446 -8577 68487 -8543
rect 67359 -8621 67400 -8587
rect 67560 -8666 67601 -8632
rect 67329 -8689 67336 -8681
rect 67340 -8723 67381 -8689
rect 67560 -8734 67601 -8700
rect 64493 -8906 64534 -8872
rect 64565 -8906 64606 -8872
rect 64637 -8906 64678 -8872
rect 64950 -8913 64991 -8879
rect 64995 -8913 65002 -8868
rect 65095 -8879 65102 -8868
rect 65106 -8913 65147 -8879
rect 65690 -8895 65731 -8861
rect 65735 -8895 65742 -8853
rect 63584 -8959 64066 -8925
rect 64918 -8949 64959 -8915
rect 64990 -8949 65031 -8915
rect 65304 -8956 65345 -8922
rect 65349 -8956 65356 -8911
rect 65449 -8922 65456 -8911
rect 65877 -8913 65889 -8845
rect 65918 -8879 65923 -8811
rect 65963 -8843 65968 -8775
rect 65997 -8809 66002 -8743
rect 67229 -8753 67236 -8741
rect 67609 -8750 67614 -8616
rect 66007 -8793 66048 -8759
rect 66210 -8838 66251 -8804
rect 65977 -8861 65984 -8853
rect 65988 -8895 66029 -8861
rect 66210 -8906 66251 -8872
rect 65460 -8956 65501 -8922
rect 63584 -8985 64053 -8959
rect 63588 -8993 63795 -8985
rect 63604 -9003 63779 -8993
rect 63330 -9140 63511 -9114
rect 62837 -9174 62878 -9140
rect 62933 -9174 62974 -9140
rect 63029 -9174 63070 -9140
rect 63125 -9174 63166 -9140
rect 63221 -9174 63262 -9140
rect 63317 -9174 63511 -9140
rect 63330 -9200 63511 -9174
rect 63530 -9174 63637 -9050
rect 63789 -9062 63795 -9051
rect 63408 -9870 63449 -9200
rect 63530 -9228 63539 -9174
rect 63215 -9936 63366 -9924
rect 62883 -9970 63366 -9936
rect 63215 -9971 63366 -9970
rect 63396 -9971 63449 -9870
rect 63542 -9971 63583 -9174
rect 63588 -9971 63594 -9174
rect 63800 -9971 63841 -9062
rect 63934 -9971 63975 -8985
rect 64187 -9002 64228 -8968
rect 64283 -9002 64324 -8968
rect 64379 -9002 64420 -8968
rect 64475 -9002 64516 -8968
rect 64571 -9002 64612 -8968
rect 64667 -9002 64708 -8968
rect 64763 -9002 64804 -8968
rect 65272 -8992 65313 -8958
rect 65344 -8992 65385 -8958
rect 65690 -8995 65731 -8961
rect 65735 -8995 65742 -8950
rect 65877 -9001 65884 -8913
rect 66259 -8922 66264 -8788
rect 65977 -8961 65984 -8950
rect 66293 -8956 66298 -8762
rect 66333 -8778 66340 -8767
rect 66329 -8809 66340 -8778
rect 66655 -8796 66696 -8762
rect 65988 -8995 66029 -8961
rect 64925 -9045 64966 -9011
rect 65021 -9045 65062 -9011
rect 65117 -9045 65158 -9011
rect 65626 -9035 65667 -9001
rect 65698 -9035 65739 -9001
rect 65770 -9035 65811 -9001
rect 65842 -9029 65884 -9001
rect 66188 -9025 66229 -8991
rect 66233 -9025 66240 -8980
rect 66329 -8992 66334 -8809
rect 66363 -8995 66368 -8812
rect 65842 -9035 65883 -9029
rect 65279 -9088 65320 -9054
rect 65375 -9088 65416 -9054
rect 65471 -9088 65512 -9054
rect 66375 -9076 66382 -8809
rect 67004 -8819 67397 -8753
rect 67643 -8784 67648 -8590
rect 67683 -8606 67690 -8595
rect 67679 -8637 67690 -8606
rect 68005 -8624 68046 -8590
rect 66391 -8860 66432 -8826
rect 66740 -8830 66757 -8819
rect 66740 -8832 66746 -8830
rect 66391 -8928 66432 -8894
rect 66443 -8995 66448 -8860
rect 66674 -8874 66746 -8832
rect 66802 -8874 67397 -8819
rect 67538 -8853 67579 -8819
rect 67583 -8853 67590 -8808
rect 67679 -8820 67684 -8637
rect 67713 -8823 67718 -8640
rect 66674 -8877 67397 -8874
rect 66477 -8980 66482 -8892
rect 66594 -8942 66635 -8908
rect 66639 -8942 66646 -8900
rect 66475 -8991 66482 -8980
rect 66477 -9025 66482 -8991
rect 66486 -9025 66527 -8991
rect 66594 -9042 66635 -9008
rect 66639 -9042 66646 -8997
rect 66487 -9078 66528 -9044
rect 66559 -9078 66600 -9044
rect 66631 -9078 66672 -9044
rect 65633 -9131 65674 -9097
rect 65729 -9131 65770 -9097
rect 65825 -9131 65866 -9097
rect 65921 -9131 65962 -9097
rect 66017 -9131 66058 -9097
rect 66674 -9114 66825 -8877
rect 67004 -8899 67397 -8877
rect 66928 -8925 67397 -8899
rect 67725 -8904 67732 -8637
rect 67741 -8688 67782 -8654
rect 67741 -8756 67782 -8722
rect 67793 -8823 67798 -8688
rect 68355 -8691 68396 -8657
rect 68407 -8718 68412 -8641
rect 67827 -8808 67832 -8720
rect 67944 -8770 67985 -8736
rect 67989 -8770 67996 -8728
rect 68089 -8740 68096 -8729
rect 68100 -8774 68141 -8740
rect 68441 -8752 68446 -8607
rect 68644 -8620 68685 -8586
rect 68689 -8620 68696 -8575
rect 68789 -8586 68796 -8575
rect 69034 -8580 69075 -8546
rect 69079 -8580 69086 -8535
rect 68800 -8620 68841 -8586
rect 68709 -8734 68750 -8700
rect 68761 -8761 68766 -8684
rect 67825 -8819 67832 -8808
rect 68294 -8813 68335 -8779
rect 68339 -8813 68346 -8771
rect 68439 -8779 68446 -8771
rect 68450 -8813 68491 -8779
rect 68795 -8795 68800 -8650
rect 69034 -8663 69075 -8629
rect 69079 -8663 69086 -8618
rect 69156 -8679 69161 -8363
rect 69179 -8379 69186 -8371
rect 69190 -8379 69195 -8363
rect 69190 -8413 69231 -8379
rect 69235 -8413 69242 -8371
rect 69179 -8462 69186 -8451
rect 69190 -8462 69195 -8413
rect 69190 -8496 69231 -8462
rect 69235 -8496 69242 -8451
rect 69179 -8546 69186 -8535
rect 69190 -8546 69195 -8496
rect 69190 -8580 69231 -8546
rect 69235 -8580 69242 -8535
rect 69179 -8629 69186 -8618
rect 69190 -8629 69195 -8580
rect 69190 -8663 69231 -8629
rect 69235 -8663 69242 -8618
rect 69179 -8697 69186 -8671
rect 69190 -8713 69195 -8663
rect 69099 -8777 69140 -8743
rect 67827 -8853 67832 -8819
rect 67836 -8853 67877 -8819
rect 67944 -8870 67985 -8836
rect 67989 -8870 67996 -8825
rect 68089 -8832 68096 -8821
rect 68100 -8866 68141 -8832
rect 68648 -8856 68689 -8822
rect 68693 -8856 68700 -8814
rect 68793 -8822 68800 -8814
rect 68804 -8856 68845 -8822
rect 69221 -8845 69228 -8697
rect 69244 -8713 69247 -8363
rect 69278 -8679 69281 -8363
rect 69335 -8379 69342 -8371
rect 69284 -8413 69325 -8379
rect 69346 -8413 69397 -8379
rect 70056 -8422 70061 -8406
rect 70079 -8422 70086 -8414
rect 70090 -8422 70095 -8406
rect 70386 -8408 70427 -8374
rect 70431 -8408 70438 -8363
rect 69335 -8462 69342 -8451
rect 69516 -8456 69557 -8422
rect 69588 -8456 69629 -8422
rect 69660 -8456 69701 -8422
rect 69804 -8456 69845 -8422
rect 69876 -8456 69989 -8422
rect 70020 -8456 70061 -8422
rect 69346 -8496 69387 -8462
rect 69335 -8546 69342 -8535
rect 69913 -8539 69954 -8505
rect 69346 -8580 69387 -8546
rect 69335 -8629 69342 -8618
rect 69346 -8663 69387 -8629
rect 69578 -8689 69619 -8655
rect 69623 -8689 69630 -8644
rect 69700 -8706 69705 -8588
rect 69723 -8655 69730 -8644
rect 69734 -8655 69739 -8622
rect 69770 -8655 69775 -8622
rect 69734 -8689 69775 -8655
rect 69779 -8689 69786 -8644
rect 69734 -8740 69739 -8689
rect 69770 -8740 69775 -8689
rect 69804 -8706 69809 -8589
rect 69913 -8623 69954 -8589
rect 69913 -8706 69954 -8672
rect 70056 -8706 70061 -8456
rect 70090 -8456 70131 -8422
rect 70079 -8505 70086 -8494
rect 70090 -8505 70095 -8456
rect 70386 -8491 70427 -8457
rect 70431 -8491 70438 -8446
rect 70090 -8539 70131 -8505
rect 70079 -8589 70086 -8578
rect 70090 -8589 70095 -8539
rect 70239 -8565 70348 -8499
rect 70508 -8507 70513 -8191
rect 70531 -8207 70538 -8199
rect 70542 -8207 70547 -8191
rect 70542 -8241 70583 -8207
rect 70587 -8241 70594 -8199
rect 70531 -8290 70538 -8279
rect 70542 -8290 70547 -8241
rect 70542 -8324 70583 -8290
rect 70587 -8324 70594 -8279
rect 70531 -8374 70538 -8363
rect 70542 -8374 70547 -8324
rect 70542 -8408 70583 -8374
rect 70587 -8408 70594 -8363
rect 70531 -8457 70538 -8446
rect 70542 -8457 70547 -8408
rect 70542 -8491 70583 -8457
rect 70587 -8491 70594 -8446
rect 70531 -8525 70538 -8499
rect 70542 -8541 70547 -8491
rect 70090 -8623 70131 -8589
rect 70451 -8605 70492 -8571
rect 70079 -8672 70086 -8661
rect 70090 -8672 70095 -8623
rect 70090 -8706 70131 -8672
rect 70573 -8673 70580 -8525
rect 70596 -8541 70599 -8191
rect 70630 -8507 70633 -8191
rect 70687 -8207 70694 -8199
rect 70636 -8241 70677 -8207
rect 70698 -8241 70749 -8207
rect 71613 -8231 71654 -8197
rect 71709 -8231 71750 -8197
rect 71805 -8231 71846 -8197
rect 73775 -8207 73782 -8199
rect 71406 -8250 71411 -8234
rect 71429 -8250 71436 -8242
rect 71440 -8250 71445 -8234
rect 70687 -8290 70694 -8279
rect 70866 -8284 70907 -8250
rect 70938 -8284 70979 -8250
rect 71010 -8284 71051 -8250
rect 71154 -8284 71195 -8250
rect 71226 -8284 71339 -8250
rect 71370 -8284 71411 -8250
rect 70698 -8324 70739 -8290
rect 70687 -8374 70694 -8363
rect 71263 -8367 71304 -8333
rect 70698 -8408 70739 -8374
rect 70687 -8457 70694 -8446
rect 70698 -8491 70739 -8457
rect 70928 -8517 70969 -8483
rect 70973 -8517 70980 -8472
rect 71050 -8534 71055 -8416
rect 71073 -8483 71080 -8472
rect 71084 -8483 71089 -8450
rect 71120 -8483 71125 -8450
rect 71084 -8517 71125 -8483
rect 71129 -8517 71136 -8472
rect 71084 -8568 71089 -8517
rect 71120 -8568 71125 -8517
rect 71154 -8534 71159 -8417
rect 71263 -8451 71304 -8417
rect 71263 -8534 71304 -8500
rect 71406 -8534 71411 -8284
rect 71440 -8284 71481 -8250
rect 71967 -8274 72008 -8240
rect 72063 -8274 72104 -8240
rect 72159 -8274 72200 -8240
rect 73666 -8241 73707 -8207
rect 73730 -8241 73782 -8207
rect 73810 -8241 73851 -8207
rect 71429 -8333 71436 -8322
rect 71440 -8333 71445 -8284
rect 71679 -8293 71686 -8285
rect 71779 -8293 71786 -8285
rect 71606 -8327 71675 -8293
rect 71678 -8327 71719 -8293
rect 71790 -8327 71831 -8293
rect 72321 -8317 72362 -8283
rect 72417 -8317 72458 -8283
rect 72513 -8317 72554 -8283
rect 72609 -8317 72650 -8283
rect 72705 -8317 72746 -8283
rect 73730 -8324 73771 -8290
rect 73775 -8324 73782 -8279
rect 71440 -8367 71481 -8333
rect 72033 -8336 72040 -8328
rect 72133 -8336 72140 -8328
rect 71429 -8417 71436 -8406
rect 71440 -8417 71445 -8367
rect 71634 -8410 71675 -8376
rect 71679 -8410 71686 -8365
rect 71779 -8376 71786 -8365
rect 71960 -8370 72029 -8336
rect 72032 -8370 72073 -8336
rect 72144 -8370 72185 -8336
rect 72869 -8360 72910 -8326
rect 72965 -8360 73006 -8326
rect 73061 -8360 73102 -8326
rect 73157 -8360 73198 -8326
rect 73253 -8360 73294 -8326
rect 73349 -8360 73390 -8326
rect 73445 -8360 73486 -8326
rect 71790 -8410 71831 -8376
rect 72423 -8379 72430 -8371
rect 71440 -8451 71481 -8417
rect 71429 -8500 71436 -8489
rect 71440 -8500 71445 -8451
rect 71634 -8494 71675 -8460
rect 71679 -8494 71686 -8449
rect 71779 -8460 71786 -8449
rect 71988 -8453 72029 -8419
rect 72033 -8453 72040 -8408
rect 72133 -8419 72140 -8408
rect 72314 -8413 72355 -8379
rect 72378 -8413 72430 -8379
rect 72458 -8413 72499 -8379
rect 72144 -8453 72185 -8419
rect 71790 -8494 71831 -8460
rect 71440 -8534 71481 -8500
rect 71440 -8568 71445 -8534
rect 70090 -8740 70095 -8706
rect 70386 -8723 70427 -8689
rect 70431 -8723 70438 -8681
rect 70573 -8741 70585 -8673
rect 70614 -8707 70619 -8639
rect 70659 -8671 70664 -8603
rect 70693 -8637 70698 -8571
rect 71634 -8577 71675 -8543
rect 71679 -8577 71686 -8532
rect 71779 -8543 71786 -8532
rect 71988 -8537 72029 -8503
rect 72033 -8537 72040 -8492
rect 72133 -8503 72140 -8492
rect 72378 -8496 72419 -8462
rect 72423 -8496 72430 -8451
rect 72144 -8537 72185 -8503
rect 71790 -8577 71831 -8543
rect 70703 -8621 70744 -8587
rect 70904 -8666 70945 -8632
rect 70673 -8689 70680 -8681
rect 70684 -8723 70725 -8689
rect 70904 -8734 70945 -8700
rect 67837 -8906 67878 -8872
rect 67909 -8906 67950 -8872
rect 67981 -8906 68022 -8872
rect 68294 -8913 68335 -8879
rect 68339 -8913 68346 -8868
rect 68439 -8879 68446 -8868
rect 68450 -8913 68491 -8879
rect 69034 -8895 69075 -8861
rect 69079 -8895 69086 -8853
rect 66928 -8959 67410 -8925
rect 68262 -8949 68303 -8915
rect 68334 -8949 68375 -8915
rect 68648 -8956 68689 -8922
rect 68693 -8956 68700 -8911
rect 68793 -8922 68800 -8911
rect 69221 -8913 69233 -8845
rect 69262 -8879 69267 -8811
rect 69307 -8843 69312 -8775
rect 69341 -8809 69346 -8743
rect 70573 -8753 70580 -8741
rect 70953 -8750 70958 -8616
rect 69351 -8793 69392 -8759
rect 69554 -8838 69595 -8804
rect 69321 -8861 69328 -8853
rect 69332 -8895 69373 -8861
rect 69554 -8906 69595 -8872
rect 68804 -8956 68845 -8922
rect 66928 -8985 67397 -8959
rect 66932 -8993 67139 -8985
rect 66948 -9003 67123 -8993
rect 66674 -9140 66855 -9114
rect 66181 -9174 66222 -9140
rect 66277 -9174 66318 -9140
rect 66373 -9174 66414 -9140
rect 66469 -9174 66510 -9140
rect 66565 -9174 66606 -9140
rect 66661 -9174 66855 -9140
rect 66674 -9200 66855 -9174
rect 66874 -9174 66981 -9050
rect 67133 -9062 67139 -9051
rect 66752 -9870 66793 -9200
rect 66874 -9228 66883 -9174
rect 66559 -9936 66710 -9924
rect 66227 -9970 66710 -9936
rect 66559 -9971 66710 -9970
rect 66740 -9971 66793 -9870
rect 66886 -9971 66927 -9174
rect 66932 -9971 66938 -9174
rect 67144 -9971 67185 -9062
rect 67278 -9971 67319 -8985
rect 67531 -9002 67572 -8968
rect 67627 -9002 67668 -8968
rect 67723 -9002 67764 -8968
rect 67819 -9002 67860 -8968
rect 67915 -9002 67956 -8968
rect 68011 -9002 68052 -8968
rect 68107 -9002 68148 -8968
rect 68616 -8992 68657 -8958
rect 68688 -8992 68729 -8958
rect 69034 -8995 69075 -8961
rect 69079 -8995 69086 -8950
rect 69221 -9001 69228 -8913
rect 69603 -8922 69608 -8788
rect 69321 -8961 69328 -8950
rect 69637 -8956 69642 -8762
rect 69677 -8778 69684 -8767
rect 69673 -8809 69684 -8778
rect 69999 -8796 70040 -8762
rect 69332 -8995 69373 -8961
rect 68269 -9045 68310 -9011
rect 68365 -9045 68406 -9011
rect 68461 -9045 68502 -9011
rect 68970 -9035 69011 -9001
rect 69042 -9035 69083 -9001
rect 69114 -9035 69155 -9001
rect 69186 -9029 69228 -9001
rect 69532 -9025 69573 -8991
rect 69577 -9025 69584 -8980
rect 69673 -8992 69678 -8809
rect 69707 -8995 69712 -8812
rect 69186 -9035 69227 -9029
rect 68623 -9088 68664 -9054
rect 68719 -9088 68760 -9054
rect 68815 -9088 68856 -9054
rect 69719 -9076 69726 -8809
rect 70348 -8819 70741 -8753
rect 70987 -8784 70992 -8590
rect 71027 -8606 71034 -8595
rect 71023 -8637 71034 -8606
rect 71349 -8624 71390 -8590
rect 69735 -8860 69776 -8826
rect 70084 -8830 70101 -8819
rect 70084 -8832 70090 -8830
rect 69735 -8928 69776 -8894
rect 69787 -8995 69792 -8860
rect 70018 -8874 70090 -8832
rect 70146 -8874 70741 -8819
rect 70882 -8853 70923 -8819
rect 70927 -8853 70934 -8808
rect 71023 -8820 71028 -8637
rect 71057 -8823 71062 -8640
rect 70018 -8877 70741 -8874
rect 69821 -8980 69826 -8892
rect 69938 -8942 69979 -8908
rect 69983 -8942 69990 -8900
rect 69819 -8991 69826 -8980
rect 69821 -9025 69826 -8991
rect 69830 -9025 69871 -8991
rect 69938 -9042 69979 -9008
rect 69983 -9042 69990 -8997
rect 69831 -9078 69872 -9044
rect 69903 -9078 69944 -9044
rect 69975 -9078 70016 -9044
rect 68977 -9131 69018 -9097
rect 69073 -9131 69114 -9097
rect 69169 -9131 69210 -9097
rect 69265 -9131 69306 -9097
rect 69361 -9131 69402 -9097
rect 70018 -9114 70169 -8877
rect 70348 -8899 70741 -8877
rect 70272 -8925 70741 -8899
rect 71069 -8904 71076 -8637
rect 71085 -8688 71126 -8654
rect 71085 -8756 71126 -8722
rect 71137 -8823 71142 -8688
rect 71699 -8691 71740 -8657
rect 71751 -8718 71756 -8641
rect 71171 -8808 71176 -8720
rect 71288 -8770 71329 -8736
rect 71333 -8770 71340 -8728
rect 71433 -8740 71440 -8729
rect 71444 -8774 71485 -8740
rect 71785 -8752 71790 -8607
rect 71988 -8620 72029 -8586
rect 72033 -8620 72040 -8575
rect 72133 -8586 72140 -8575
rect 72378 -8580 72419 -8546
rect 72423 -8580 72430 -8535
rect 72144 -8620 72185 -8586
rect 72053 -8734 72094 -8700
rect 72105 -8761 72110 -8684
rect 71169 -8819 71176 -8808
rect 71638 -8813 71679 -8779
rect 71683 -8813 71690 -8771
rect 71783 -8779 71790 -8771
rect 71794 -8813 71835 -8779
rect 72139 -8795 72144 -8650
rect 72378 -8663 72419 -8629
rect 72423 -8663 72430 -8618
rect 72500 -8679 72505 -8363
rect 72523 -8379 72530 -8371
rect 72534 -8379 72539 -8363
rect 72534 -8413 72575 -8379
rect 72579 -8413 72586 -8371
rect 72523 -8462 72530 -8451
rect 72534 -8462 72539 -8413
rect 72534 -8496 72575 -8462
rect 72579 -8496 72586 -8451
rect 72523 -8546 72530 -8535
rect 72534 -8546 72539 -8496
rect 72534 -8580 72575 -8546
rect 72579 -8580 72586 -8535
rect 72523 -8629 72530 -8618
rect 72534 -8629 72539 -8580
rect 72534 -8663 72575 -8629
rect 72579 -8663 72586 -8618
rect 72523 -8697 72530 -8671
rect 72534 -8713 72539 -8663
rect 72443 -8777 72484 -8743
rect 71171 -8853 71176 -8819
rect 71180 -8853 71221 -8819
rect 71288 -8870 71329 -8836
rect 71333 -8870 71340 -8825
rect 71433 -8832 71440 -8821
rect 71444 -8866 71485 -8832
rect 71992 -8856 72033 -8822
rect 72037 -8856 72044 -8814
rect 72137 -8822 72144 -8814
rect 72148 -8856 72189 -8822
rect 72565 -8845 72572 -8697
rect 72588 -8713 72591 -8363
rect 72622 -8679 72625 -8363
rect 72679 -8379 72686 -8371
rect 72628 -8413 72669 -8379
rect 72690 -8413 72741 -8379
rect 73400 -8422 73405 -8406
rect 73423 -8422 73430 -8414
rect 73434 -8422 73439 -8406
rect 73730 -8408 73771 -8374
rect 73775 -8408 73782 -8363
rect 72679 -8462 72686 -8451
rect 72860 -8456 72901 -8422
rect 72932 -8456 72973 -8422
rect 73004 -8456 73045 -8422
rect 73148 -8456 73189 -8422
rect 73220 -8456 73333 -8422
rect 73364 -8456 73405 -8422
rect 72690 -8496 72731 -8462
rect 72679 -8546 72686 -8535
rect 73257 -8539 73298 -8505
rect 72690 -8580 72731 -8546
rect 72679 -8629 72686 -8618
rect 72690 -8663 72731 -8629
rect 72922 -8689 72963 -8655
rect 72967 -8689 72974 -8644
rect 73044 -8706 73049 -8588
rect 73067 -8655 73074 -8644
rect 73078 -8655 73083 -8622
rect 73114 -8655 73119 -8622
rect 73078 -8689 73119 -8655
rect 73123 -8689 73130 -8644
rect 73078 -8740 73083 -8689
rect 73114 -8740 73119 -8689
rect 73148 -8706 73153 -8589
rect 73257 -8623 73298 -8589
rect 73257 -8706 73298 -8672
rect 73400 -8706 73405 -8456
rect 73434 -8456 73475 -8422
rect 73423 -8505 73430 -8494
rect 73434 -8505 73439 -8456
rect 73730 -8491 73771 -8457
rect 73775 -8491 73782 -8446
rect 73434 -8539 73475 -8505
rect 73423 -8589 73430 -8578
rect 73434 -8589 73439 -8539
rect 73583 -8565 73692 -8499
rect 73852 -8507 73857 -8191
rect 73875 -8207 73882 -8199
rect 73886 -8207 73891 -8191
rect 73886 -8241 73927 -8207
rect 73931 -8241 73938 -8199
rect 73875 -8290 73882 -8279
rect 73886 -8290 73891 -8241
rect 73886 -8324 73927 -8290
rect 73931 -8324 73938 -8279
rect 73875 -8374 73882 -8363
rect 73886 -8374 73891 -8324
rect 73886 -8408 73927 -8374
rect 73931 -8408 73938 -8363
rect 73875 -8457 73882 -8446
rect 73886 -8457 73891 -8408
rect 73886 -8491 73927 -8457
rect 73931 -8491 73938 -8446
rect 73875 -8525 73882 -8499
rect 73886 -8541 73891 -8491
rect 73434 -8623 73475 -8589
rect 73795 -8605 73836 -8571
rect 73423 -8672 73430 -8661
rect 73434 -8672 73439 -8623
rect 73434 -8706 73475 -8672
rect 73917 -8673 73924 -8525
rect 73940 -8541 73943 -8191
rect 73974 -8507 73977 -8191
rect 74031 -8207 74038 -8199
rect 73980 -8241 74021 -8207
rect 74042 -8241 74093 -8207
rect 74957 -8231 74998 -8197
rect 75053 -8231 75094 -8197
rect 75149 -8231 75190 -8197
rect 77119 -8207 77126 -8199
rect 74750 -8250 74755 -8234
rect 74773 -8250 74780 -8242
rect 74784 -8250 74789 -8234
rect 74031 -8290 74038 -8279
rect 74210 -8284 74251 -8250
rect 74282 -8284 74323 -8250
rect 74354 -8284 74395 -8250
rect 74498 -8284 74539 -8250
rect 74570 -8284 74683 -8250
rect 74714 -8284 74755 -8250
rect 74042 -8324 74083 -8290
rect 74031 -8374 74038 -8363
rect 74607 -8367 74648 -8333
rect 74042 -8408 74083 -8374
rect 74031 -8457 74038 -8446
rect 74042 -8491 74083 -8457
rect 74272 -8517 74313 -8483
rect 74317 -8517 74324 -8472
rect 74394 -8534 74399 -8416
rect 74417 -8483 74424 -8472
rect 74428 -8483 74433 -8450
rect 74464 -8483 74469 -8450
rect 74428 -8517 74469 -8483
rect 74473 -8517 74480 -8472
rect 74428 -8568 74433 -8517
rect 74464 -8568 74469 -8517
rect 74498 -8534 74503 -8417
rect 74607 -8451 74648 -8417
rect 74607 -8534 74648 -8500
rect 74750 -8534 74755 -8284
rect 74784 -8284 74825 -8250
rect 75311 -8274 75352 -8240
rect 75407 -8274 75448 -8240
rect 75503 -8274 75544 -8240
rect 77010 -8241 77051 -8207
rect 77074 -8241 77126 -8207
rect 77154 -8241 77195 -8207
rect 74773 -8333 74780 -8322
rect 74784 -8333 74789 -8284
rect 75023 -8293 75030 -8285
rect 75123 -8293 75130 -8285
rect 74950 -8327 75019 -8293
rect 75022 -8327 75063 -8293
rect 75134 -8327 75175 -8293
rect 75665 -8317 75706 -8283
rect 75761 -8317 75802 -8283
rect 75857 -8317 75898 -8283
rect 75953 -8317 75994 -8283
rect 76049 -8317 76090 -8283
rect 77074 -8324 77115 -8290
rect 77119 -8324 77126 -8279
rect 74784 -8367 74825 -8333
rect 75377 -8336 75384 -8328
rect 75477 -8336 75484 -8328
rect 74773 -8417 74780 -8406
rect 74784 -8417 74789 -8367
rect 74978 -8410 75019 -8376
rect 75023 -8410 75030 -8365
rect 75123 -8376 75130 -8365
rect 75304 -8370 75373 -8336
rect 75376 -8370 75417 -8336
rect 75488 -8370 75529 -8336
rect 76213 -8360 76254 -8326
rect 76309 -8360 76350 -8326
rect 76405 -8360 76446 -8326
rect 76501 -8360 76542 -8326
rect 76597 -8360 76638 -8326
rect 76693 -8360 76734 -8326
rect 76789 -8360 76830 -8326
rect 75134 -8410 75175 -8376
rect 75767 -8379 75774 -8371
rect 74784 -8451 74825 -8417
rect 74773 -8500 74780 -8489
rect 74784 -8500 74789 -8451
rect 74978 -8494 75019 -8460
rect 75023 -8494 75030 -8449
rect 75123 -8460 75130 -8449
rect 75332 -8453 75373 -8419
rect 75377 -8453 75384 -8408
rect 75477 -8419 75484 -8408
rect 75658 -8413 75699 -8379
rect 75722 -8413 75774 -8379
rect 75802 -8413 75843 -8379
rect 75488 -8453 75529 -8419
rect 75134 -8494 75175 -8460
rect 74784 -8534 74825 -8500
rect 74784 -8568 74789 -8534
rect 73434 -8740 73439 -8706
rect 73730 -8723 73771 -8689
rect 73775 -8723 73782 -8681
rect 73917 -8741 73929 -8673
rect 73958 -8707 73963 -8639
rect 74003 -8671 74008 -8603
rect 74037 -8637 74042 -8571
rect 74978 -8577 75019 -8543
rect 75023 -8577 75030 -8532
rect 75123 -8543 75130 -8532
rect 75332 -8537 75373 -8503
rect 75377 -8537 75384 -8492
rect 75477 -8503 75484 -8492
rect 75722 -8496 75763 -8462
rect 75767 -8496 75774 -8451
rect 75488 -8537 75529 -8503
rect 75134 -8577 75175 -8543
rect 74047 -8621 74088 -8587
rect 74248 -8666 74289 -8632
rect 74017 -8689 74024 -8681
rect 74028 -8723 74069 -8689
rect 74248 -8734 74289 -8700
rect 71181 -8906 71222 -8872
rect 71253 -8906 71294 -8872
rect 71325 -8906 71366 -8872
rect 71638 -8913 71679 -8879
rect 71683 -8913 71690 -8868
rect 71783 -8879 71790 -8868
rect 71794 -8913 71835 -8879
rect 72378 -8895 72419 -8861
rect 72423 -8895 72430 -8853
rect 70272 -8959 70754 -8925
rect 71606 -8949 71647 -8915
rect 71678 -8949 71719 -8915
rect 71992 -8956 72033 -8922
rect 72037 -8956 72044 -8911
rect 72137 -8922 72144 -8911
rect 72565 -8913 72577 -8845
rect 72606 -8879 72611 -8811
rect 72651 -8843 72656 -8775
rect 72685 -8809 72690 -8743
rect 73917 -8753 73924 -8741
rect 74297 -8750 74302 -8616
rect 72695 -8793 72736 -8759
rect 72898 -8838 72939 -8804
rect 72665 -8861 72672 -8853
rect 72676 -8895 72717 -8861
rect 72898 -8906 72939 -8872
rect 72148 -8956 72189 -8922
rect 70272 -8985 70741 -8959
rect 70276 -8993 70483 -8985
rect 70292 -9003 70467 -8993
rect 70018 -9140 70199 -9114
rect 69525 -9174 69566 -9140
rect 69621 -9174 69662 -9140
rect 69717 -9174 69758 -9140
rect 69813 -9174 69854 -9140
rect 69909 -9174 69950 -9140
rect 70005 -9174 70199 -9140
rect 70018 -9200 70199 -9174
rect 70218 -9174 70325 -9050
rect 70477 -9062 70483 -9051
rect 70096 -9870 70137 -9200
rect 70218 -9228 70227 -9174
rect 69903 -9936 70054 -9924
rect 69571 -9970 70054 -9936
rect 69903 -9971 70054 -9970
rect 70084 -9971 70137 -9870
rect 70230 -9971 70271 -9174
rect 70276 -9971 70282 -9174
rect 70488 -9971 70529 -9062
rect 70622 -9971 70663 -8985
rect 70875 -9002 70916 -8968
rect 70971 -9002 71012 -8968
rect 71067 -9002 71108 -8968
rect 71163 -9002 71204 -8968
rect 71259 -9002 71300 -8968
rect 71355 -9002 71396 -8968
rect 71451 -9002 71492 -8968
rect 71960 -8992 72001 -8958
rect 72032 -8992 72073 -8958
rect 72378 -8995 72419 -8961
rect 72423 -8995 72430 -8950
rect 72565 -9001 72572 -8913
rect 72947 -8922 72952 -8788
rect 72665 -8961 72672 -8950
rect 72981 -8956 72986 -8762
rect 73021 -8778 73028 -8767
rect 73017 -8809 73028 -8778
rect 73343 -8796 73384 -8762
rect 72676 -8995 72717 -8961
rect 71613 -9045 71654 -9011
rect 71709 -9045 71750 -9011
rect 71805 -9045 71846 -9011
rect 72314 -9035 72355 -9001
rect 72386 -9035 72427 -9001
rect 72458 -9035 72499 -9001
rect 72530 -9029 72572 -9001
rect 72876 -9025 72917 -8991
rect 72921 -9025 72928 -8980
rect 73017 -8992 73022 -8809
rect 73051 -8995 73056 -8812
rect 72530 -9035 72571 -9029
rect 71967 -9088 72008 -9054
rect 72063 -9088 72104 -9054
rect 72159 -9088 72200 -9054
rect 73063 -9076 73070 -8809
rect 73692 -8819 74085 -8753
rect 74331 -8784 74336 -8590
rect 74371 -8606 74378 -8595
rect 74367 -8637 74378 -8606
rect 74693 -8624 74734 -8590
rect 73079 -8860 73120 -8826
rect 73428 -8830 73445 -8819
rect 73428 -8832 73434 -8830
rect 73079 -8928 73120 -8894
rect 73131 -8995 73136 -8860
rect 73362 -8874 73434 -8832
rect 73490 -8874 74085 -8819
rect 74226 -8853 74267 -8819
rect 74271 -8853 74278 -8808
rect 74367 -8820 74372 -8637
rect 74401 -8823 74406 -8640
rect 73362 -8877 74085 -8874
rect 73165 -8980 73170 -8892
rect 73282 -8942 73323 -8908
rect 73327 -8942 73334 -8900
rect 73163 -8991 73170 -8980
rect 73165 -9025 73170 -8991
rect 73174 -9025 73215 -8991
rect 73282 -9042 73323 -9008
rect 73327 -9042 73334 -8997
rect 73175 -9078 73216 -9044
rect 73247 -9078 73288 -9044
rect 73319 -9078 73360 -9044
rect 72321 -9131 72362 -9097
rect 72417 -9131 72458 -9097
rect 72513 -9131 72554 -9097
rect 72609 -9131 72650 -9097
rect 72705 -9131 72746 -9097
rect 73362 -9114 73513 -8877
rect 73692 -8899 74085 -8877
rect 73616 -8925 74085 -8899
rect 74413 -8904 74420 -8637
rect 74429 -8688 74470 -8654
rect 74429 -8756 74470 -8722
rect 74481 -8823 74486 -8688
rect 75043 -8691 75084 -8657
rect 75095 -8718 75100 -8641
rect 74515 -8808 74520 -8720
rect 74632 -8770 74673 -8736
rect 74677 -8770 74684 -8728
rect 74777 -8740 74784 -8729
rect 74788 -8774 74829 -8740
rect 75129 -8752 75134 -8607
rect 75332 -8620 75373 -8586
rect 75377 -8620 75384 -8575
rect 75477 -8586 75484 -8575
rect 75722 -8580 75763 -8546
rect 75767 -8580 75774 -8535
rect 75488 -8620 75529 -8586
rect 75397 -8734 75438 -8700
rect 75449 -8761 75454 -8684
rect 74513 -8819 74520 -8808
rect 74982 -8813 75023 -8779
rect 75027 -8813 75034 -8771
rect 75127 -8779 75134 -8771
rect 75138 -8813 75179 -8779
rect 75483 -8795 75488 -8650
rect 75722 -8663 75763 -8629
rect 75767 -8663 75774 -8618
rect 75844 -8679 75849 -8363
rect 75867 -8379 75874 -8371
rect 75878 -8379 75883 -8363
rect 75878 -8413 75919 -8379
rect 75923 -8413 75930 -8371
rect 75867 -8462 75874 -8451
rect 75878 -8462 75883 -8413
rect 75878 -8496 75919 -8462
rect 75923 -8496 75930 -8451
rect 75867 -8546 75874 -8535
rect 75878 -8546 75883 -8496
rect 75878 -8580 75919 -8546
rect 75923 -8580 75930 -8535
rect 75867 -8629 75874 -8618
rect 75878 -8629 75883 -8580
rect 75878 -8663 75919 -8629
rect 75923 -8663 75930 -8618
rect 75867 -8697 75874 -8671
rect 75878 -8713 75883 -8663
rect 75787 -8777 75828 -8743
rect 74515 -8853 74520 -8819
rect 74524 -8853 74565 -8819
rect 74632 -8870 74673 -8836
rect 74677 -8870 74684 -8825
rect 74777 -8832 74784 -8821
rect 74788 -8866 74829 -8832
rect 75336 -8856 75377 -8822
rect 75381 -8856 75388 -8814
rect 75481 -8822 75488 -8814
rect 75492 -8856 75533 -8822
rect 75909 -8845 75916 -8697
rect 75932 -8713 75935 -8363
rect 75966 -8679 75969 -8363
rect 76023 -8379 76030 -8371
rect 75972 -8413 76013 -8379
rect 76034 -8413 76085 -8379
rect 76744 -8422 76749 -8406
rect 76767 -8422 76774 -8414
rect 76778 -8422 76783 -8406
rect 77074 -8408 77115 -8374
rect 77119 -8408 77126 -8363
rect 76023 -8462 76030 -8451
rect 76204 -8456 76245 -8422
rect 76276 -8456 76317 -8422
rect 76348 -8456 76389 -8422
rect 76492 -8456 76533 -8422
rect 76564 -8456 76677 -8422
rect 76708 -8456 76749 -8422
rect 76034 -8496 76075 -8462
rect 76023 -8546 76030 -8535
rect 76601 -8539 76642 -8505
rect 76034 -8580 76075 -8546
rect 76023 -8629 76030 -8618
rect 76034 -8663 76075 -8629
rect 76266 -8689 76307 -8655
rect 76311 -8689 76318 -8644
rect 76388 -8706 76393 -8588
rect 76411 -8655 76418 -8644
rect 76422 -8655 76427 -8622
rect 76458 -8655 76463 -8622
rect 76422 -8689 76463 -8655
rect 76467 -8689 76474 -8644
rect 76422 -8740 76427 -8689
rect 76458 -8740 76463 -8689
rect 76492 -8706 76497 -8589
rect 76601 -8623 76642 -8589
rect 76601 -8706 76642 -8672
rect 76744 -8706 76749 -8456
rect 76778 -8456 76819 -8422
rect 76767 -8505 76774 -8494
rect 76778 -8505 76783 -8456
rect 77074 -8491 77115 -8457
rect 77119 -8491 77126 -8446
rect 76778 -8539 76819 -8505
rect 76767 -8589 76774 -8578
rect 76778 -8589 76783 -8539
rect 76927 -8565 77036 -8499
rect 77196 -8507 77201 -8191
rect 77219 -8207 77226 -8199
rect 77230 -8207 77235 -8191
rect 77230 -8241 77271 -8207
rect 77275 -8241 77282 -8199
rect 77219 -8290 77226 -8279
rect 77230 -8290 77235 -8241
rect 77230 -8324 77271 -8290
rect 77275 -8324 77282 -8279
rect 77219 -8374 77226 -8363
rect 77230 -8374 77235 -8324
rect 77230 -8408 77271 -8374
rect 77275 -8408 77282 -8363
rect 77219 -8457 77226 -8446
rect 77230 -8457 77235 -8408
rect 77230 -8491 77271 -8457
rect 77275 -8491 77282 -8446
rect 77219 -8525 77226 -8499
rect 77230 -8541 77235 -8491
rect 76778 -8623 76819 -8589
rect 77139 -8605 77180 -8571
rect 76767 -8672 76774 -8661
rect 76778 -8672 76783 -8623
rect 76778 -8706 76819 -8672
rect 77261 -8673 77268 -8525
rect 77284 -8541 77287 -8191
rect 77318 -8507 77321 -8191
rect 77375 -8207 77382 -8199
rect 77324 -8241 77365 -8207
rect 77386 -8241 77437 -8207
rect 78301 -8231 78342 -8197
rect 78397 -8231 78438 -8197
rect 78493 -8231 78534 -8197
rect 80463 -8207 80470 -8199
rect 78094 -8250 78099 -8234
rect 78117 -8250 78124 -8242
rect 78128 -8250 78133 -8234
rect 77375 -8290 77382 -8279
rect 77554 -8284 77595 -8250
rect 77626 -8284 77667 -8250
rect 77698 -8284 77739 -8250
rect 77842 -8284 77883 -8250
rect 77914 -8284 78027 -8250
rect 78058 -8284 78099 -8250
rect 77386 -8324 77427 -8290
rect 77375 -8374 77382 -8363
rect 77951 -8367 77992 -8333
rect 77386 -8408 77427 -8374
rect 77375 -8457 77382 -8446
rect 77386 -8491 77427 -8457
rect 77616 -8517 77657 -8483
rect 77661 -8517 77668 -8472
rect 77738 -8534 77743 -8416
rect 77761 -8483 77768 -8472
rect 77772 -8483 77777 -8450
rect 77808 -8483 77813 -8450
rect 77772 -8517 77813 -8483
rect 77817 -8517 77824 -8472
rect 77772 -8568 77777 -8517
rect 77808 -8568 77813 -8517
rect 77842 -8534 77847 -8417
rect 77951 -8451 77992 -8417
rect 77951 -8534 77992 -8500
rect 78094 -8534 78099 -8284
rect 78128 -8284 78169 -8250
rect 78655 -8274 78696 -8240
rect 78751 -8274 78792 -8240
rect 78847 -8274 78888 -8240
rect 80354 -8241 80395 -8207
rect 80418 -8241 80470 -8207
rect 80498 -8241 80539 -8207
rect 78117 -8333 78124 -8322
rect 78128 -8333 78133 -8284
rect 78367 -8293 78374 -8285
rect 78467 -8293 78474 -8285
rect 78294 -8327 78363 -8293
rect 78366 -8327 78407 -8293
rect 78478 -8327 78519 -8293
rect 79009 -8317 79050 -8283
rect 79105 -8317 79146 -8283
rect 79201 -8317 79242 -8283
rect 79297 -8317 79338 -8283
rect 79393 -8317 79434 -8283
rect 80418 -8324 80459 -8290
rect 80463 -8324 80470 -8279
rect 78128 -8367 78169 -8333
rect 78721 -8336 78728 -8328
rect 78821 -8336 78828 -8328
rect 78117 -8417 78124 -8406
rect 78128 -8417 78133 -8367
rect 78322 -8410 78363 -8376
rect 78367 -8410 78374 -8365
rect 78467 -8376 78474 -8365
rect 78648 -8370 78717 -8336
rect 78720 -8370 78761 -8336
rect 78832 -8370 78873 -8336
rect 79557 -8360 79598 -8326
rect 79653 -8360 79694 -8326
rect 79749 -8360 79790 -8326
rect 79845 -8360 79886 -8326
rect 79941 -8360 79982 -8326
rect 80037 -8360 80078 -8326
rect 80133 -8360 80174 -8326
rect 78478 -8410 78519 -8376
rect 79111 -8379 79118 -8371
rect 78128 -8451 78169 -8417
rect 78117 -8500 78124 -8489
rect 78128 -8500 78133 -8451
rect 78322 -8494 78363 -8460
rect 78367 -8494 78374 -8449
rect 78467 -8460 78474 -8449
rect 78676 -8453 78717 -8419
rect 78721 -8453 78728 -8408
rect 78821 -8419 78828 -8408
rect 79002 -8413 79043 -8379
rect 79066 -8413 79118 -8379
rect 79146 -8413 79187 -8379
rect 78832 -8453 78873 -8419
rect 78478 -8494 78519 -8460
rect 78128 -8534 78169 -8500
rect 78128 -8568 78133 -8534
rect 76778 -8740 76783 -8706
rect 77074 -8723 77115 -8689
rect 77119 -8723 77126 -8681
rect 77261 -8741 77273 -8673
rect 77302 -8707 77307 -8639
rect 77347 -8671 77352 -8603
rect 77381 -8637 77386 -8571
rect 78322 -8577 78363 -8543
rect 78367 -8577 78374 -8532
rect 78467 -8543 78474 -8532
rect 78676 -8537 78717 -8503
rect 78721 -8537 78728 -8492
rect 78821 -8503 78828 -8492
rect 79066 -8496 79107 -8462
rect 79111 -8496 79118 -8451
rect 78832 -8537 78873 -8503
rect 78478 -8577 78519 -8543
rect 77391 -8621 77432 -8587
rect 77592 -8666 77633 -8632
rect 77361 -8689 77368 -8681
rect 77372 -8723 77413 -8689
rect 77592 -8734 77633 -8700
rect 74525 -8906 74566 -8872
rect 74597 -8906 74638 -8872
rect 74669 -8906 74710 -8872
rect 74982 -8913 75023 -8879
rect 75027 -8913 75034 -8868
rect 75127 -8879 75134 -8868
rect 75138 -8913 75179 -8879
rect 75722 -8895 75763 -8861
rect 75767 -8895 75774 -8853
rect 73616 -8959 74098 -8925
rect 74950 -8949 74991 -8915
rect 75022 -8949 75063 -8915
rect 75336 -8956 75377 -8922
rect 75381 -8956 75388 -8911
rect 75481 -8922 75488 -8911
rect 75909 -8913 75921 -8845
rect 75950 -8879 75955 -8811
rect 75995 -8843 76000 -8775
rect 76029 -8809 76034 -8743
rect 77261 -8753 77268 -8741
rect 77641 -8750 77646 -8616
rect 76039 -8793 76080 -8759
rect 76242 -8838 76283 -8804
rect 76009 -8861 76016 -8853
rect 76020 -8895 76061 -8861
rect 76242 -8906 76283 -8872
rect 75492 -8956 75533 -8922
rect 73616 -8985 74085 -8959
rect 73620 -8993 73827 -8985
rect 73636 -9003 73811 -8993
rect 73362 -9140 73543 -9114
rect 72869 -9174 72910 -9140
rect 72965 -9174 73006 -9140
rect 73061 -9174 73102 -9140
rect 73157 -9174 73198 -9140
rect 73253 -9174 73294 -9140
rect 73349 -9174 73543 -9140
rect 73362 -9200 73543 -9174
rect 73562 -9174 73669 -9050
rect 73821 -9062 73827 -9051
rect 73440 -9870 73481 -9200
rect 73562 -9228 73571 -9174
rect 73247 -9936 73398 -9924
rect 72915 -9970 73398 -9936
rect 73247 -9971 73398 -9970
rect 73428 -9971 73481 -9870
rect 73574 -9971 73615 -9174
rect 73620 -9971 73626 -9174
rect 73832 -9971 73873 -9062
rect 73966 -9971 74007 -8985
rect 74219 -9002 74260 -8968
rect 74315 -9002 74356 -8968
rect 74411 -9002 74452 -8968
rect 74507 -9002 74548 -8968
rect 74603 -9002 74644 -8968
rect 74699 -9002 74740 -8968
rect 74795 -9002 74836 -8968
rect 75304 -8992 75345 -8958
rect 75376 -8992 75417 -8958
rect 75722 -8995 75763 -8961
rect 75767 -8995 75774 -8950
rect 75909 -9001 75916 -8913
rect 76291 -8922 76296 -8788
rect 76009 -8961 76016 -8950
rect 76325 -8956 76330 -8762
rect 76365 -8778 76372 -8767
rect 76361 -8809 76372 -8778
rect 76687 -8796 76728 -8762
rect 76020 -8995 76061 -8961
rect 74957 -9045 74998 -9011
rect 75053 -9045 75094 -9011
rect 75149 -9045 75190 -9011
rect 75658 -9035 75699 -9001
rect 75730 -9035 75771 -9001
rect 75802 -9035 75843 -9001
rect 75874 -9029 75916 -9001
rect 76220 -9025 76261 -8991
rect 76265 -9025 76272 -8980
rect 76361 -8992 76366 -8809
rect 76395 -8995 76400 -8812
rect 75874 -9035 75915 -9029
rect 75311 -9088 75352 -9054
rect 75407 -9088 75448 -9054
rect 75503 -9088 75544 -9054
rect 76407 -9076 76414 -8809
rect 77036 -8819 77429 -8753
rect 77675 -8784 77680 -8590
rect 77715 -8606 77722 -8595
rect 77711 -8637 77722 -8606
rect 78037 -8624 78078 -8590
rect 76423 -8860 76464 -8826
rect 76772 -8830 76789 -8819
rect 76772 -8832 76778 -8830
rect 76423 -8928 76464 -8894
rect 76475 -8995 76480 -8860
rect 76706 -8874 76778 -8832
rect 76834 -8874 77429 -8819
rect 77570 -8853 77611 -8819
rect 77615 -8853 77622 -8808
rect 77711 -8820 77716 -8637
rect 77745 -8823 77750 -8640
rect 76706 -8877 77429 -8874
rect 76509 -8980 76514 -8892
rect 76626 -8942 76667 -8908
rect 76671 -8942 76678 -8900
rect 76507 -8991 76514 -8980
rect 76509 -9025 76514 -8991
rect 76518 -9025 76559 -8991
rect 76626 -9042 76667 -9008
rect 76671 -9042 76678 -8997
rect 76519 -9078 76560 -9044
rect 76591 -9078 76632 -9044
rect 76663 -9078 76704 -9044
rect 75665 -9131 75706 -9097
rect 75761 -9131 75802 -9097
rect 75857 -9131 75898 -9097
rect 75953 -9131 75994 -9097
rect 76049 -9131 76090 -9097
rect 76706 -9114 76857 -8877
rect 77036 -8899 77429 -8877
rect 76960 -8925 77429 -8899
rect 77757 -8904 77764 -8637
rect 77773 -8688 77814 -8654
rect 77773 -8756 77814 -8722
rect 77825 -8823 77830 -8688
rect 78387 -8691 78428 -8657
rect 78439 -8718 78444 -8641
rect 77859 -8808 77864 -8720
rect 77976 -8770 78017 -8736
rect 78021 -8770 78028 -8728
rect 78121 -8740 78128 -8729
rect 78132 -8774 78173 -8740
rect 78473 -8752 78478 -8607
rect 78676 -8620 78717 -8586
rect 78721 -8620 78728 -8575
rect 78821 -8586 78828 -8575
rect 79066 -8580 79107 -8546
rect 79111 -8580 79118 -8535
rect 78832 -8620 78873 -8586
rect 78741 -8734 78782 -8700
rect 78793 -8761 78798 -8684
rect 77857 -8819 77864 -8808
rect 78326 -8813 78367 -8779
rect 78371 -8813 78378 -8771
rect 78471 -8779 78478 -8771
rect 78482 -8813 78523 -8779
rect 78827 -8795 78832 -8650
rect 79066 -8663 79107 -8629
rect 79111 -8663 79118 -8618
rect 79188 -8679 79193 -8363
rect 79211 -8379 79218 -8371
rect 79222 -8379 79227 -8363
rect 79222 -8413 79263 -8379
rect 79267 -8413 79274 -8371
rect 79211 -8462 79218 -8451
rect 79222 -8462 79227 -8413
rect 79222 -8496 79263 -8462
rect 79267 -8496 79274 -8451
rect 79211 -8546 79218 -8535
rect 79222 -8546 79227 -8496
rect 79222 -8580 79263 -8546
rect 79267 -8580 79274 -8535
rect 79211 -8629 79218 -8618
rect 79222 -8629 79227 -8580
rect 79222 -8663 79263 -8629
rect 79267 -8663 79274 -8618
rect 79211 -8697 79218 -8671
rect 79222 -8713 79227 -8663
rect 79131 -8777 79172 -8743
rect 77859 -8853 77864 -8819
rect 77868 -8853 77909 -8819
rect 77976 -8870 78017 -8836
rect 78021 -8870 78028 -8825
rect 78121 -8832 78128 -8821
rect 78132 -8866 78173 -8832
rect 78680 -8856 78721 -8822
rect 78725 -8856 78732 -8814
rect 78825 -8822 78832 -8814
rect 78836 -8856 78877 -8822
rect 79253 -8845 79260 -8697
rect 79276 -8713 79279 -8363
rect 79310 -8679 79313 -8363
rect 79367 -8379 79374 -8371
rect 79316 -8413 79357 -8379
rect 79378 -8413 79429 -8379
rect 80088 -8422 80093 -8406
rect 80111 -8422 80118 -8414
rect 80122 -8422 80127 -8406
rect 80418 -8408 80459 -8374
rect 80463 -8408 80470 -8363
rect 79367 -8462 79374 -8451
rect 79548 -8456 79589 -8422
rect 79620 -8456 79661 -8422
rect 79692 -8456 79733 -8422
rect 79836 -8456 79877 -8422
rect 79908 -8456 80021 -8422
rect 80052 -8456 80093 -8422
rect 79378 -8496 79419 -8462
rect 79367 -8546 79374 -8535
rect 79945 -8539 79986 -8505
rect 79378 -8580 79419 -8546
rect 79367 -8629 79374 -8618
rect 79378 -8663 79419 -8629
rect 79610 -8689 79651 -8655
rect 79655 -8689 79662 -8644
rect 79732 -8706 79737 -8588
rect 79755 -8655 79762 -8644
rect 79766 -8655 79771 -8622
rect 79802 -8655 79807 -8622
rect 79766 -8689 79807 -8655
rect 79811 -8689 79818 -8644
rect 79766 -8740 79771 -8689
rect 79802 -8740 79807 -8689
rect 79836 -8706 79841 -8589
rect 79945 -8623 79986 -8589
rect 79945 -8706 79986 -8672
rect 80088 -8706 80093 -8456
rect 80122 -8456 80163 -8422
rect 80111 -8505 80118 -8494
rect 80122 -8505 80127 -8456
rect 80418 -8491 80459 -8457
rect 80463 -8491 80470 -8446
rect 80122 -8539 80163 -8505
rect 80111 -8589 80118 -8578
rect 80122 -8589 80127 -8539
rect 80271 -8565 80380 -8499
rect 80540 -8507 80545 -8191
rect 80563 -8207 80570 -8199
rect 80574 -8207 80579 -8191
rect 80574 -8241 80615 -8207
rect 80619 -8241 80626 -8199
rect 80563 -8290 80570 -8279
rect 80574 -8290 80579 -8241
rect 80574 -8324 80615 -8290
rect 80619 -8324 80626 -8279
rect 80563 -8374 80570 -8363
rect 80574 -8374 80579 -8324
rect 80574 -8408 80615 -8374
rect 80619 -8408 80626 -8363
rect 80563 -8457 80570 -8446
rect 80574 -8457 80579 -8408
rect 80574 -8491 80615 -8457
rect 80619 -8491 80626 -8446
rect 80563 -8525 80570 -8499
rect 80574 -8541 80579 -8491
rect 80122 -8623 80163 -8589
rect 80483 -8605 80524 -8571
rect 80111 -8672 80118 -8661
rect 80122 -8672 80127 -8623
rect 80122 -8706 80163 -8672
rect 80605 -8673 80612 -8525
rect 80628 -8541 80631 -8191
rect 80662 -8507 80665 -8191
rect 80719 -8207 80726 -8199
rect 80668 -8241 80709 -8207
rect 80730 -8241 80781 -8207
rect 81645 -8231 81686 -8197
rect 81741 -8231 81782 -8197
rect 81837 -8231 81878 -8197
rect 83807 -8207 83814 -8199
rect 81438 -8250 81443 -8234
rect 81461 -8250 81468 -8242
rect 81472 -8250 81477 -8234
rect 80719 -8290 80726 -8279
rect 80898 -8284 80939 -8250
rect 80970 -8284 81011 -8250
rect 81042 -8284 81083 -8250
rect 81186 -8284 81227 -8250
rect 81258 -8284 81371 -8250
rect 81402 -8284 81443 -8250
rect 80730 -8324 80771 -8290
rect 80719 -8374 80726 -8363
rect 81295 -8367 81336 -8333
rect 80730 -8408 80771 -8374
rect 80719 -8457 80726 -8446
rect 80730 -8491 80771 -8457
rect 80960 -8517 81001 -8483
rect 81005 -8517 81012 -8472
rect 81082 -8534 81087 -8416
rect 81105 -8483 81112 -8472
rect 81116 -8483 81121 -8450
rect 81152 -8483 81157 -8450
rect 81116 -8517 81157 -8483
rect 81161 -8517 81168 -8472
rect 81116 -8568 81121 -8517
rect 81152 -8568 81157 -8517
rect 81186 -8534 81191 -8417
rect 81295 -8451 81336 -8417
rect 81295 -8534 81336 -8500
rect 81438 -8534 81443 -8284
rect 81472 -8284 81513 -8250
rect 81999 -8274 82040 -8240
rect 82095 -8274 82136 -8240
rect 82191 -8274 82232 -8240
rect 83698 -8241 83739 -8207
rect 83762 -8241 83814 -8207
rect 83842 -8241 83883 -8207
rect 81461 -8333 81468 -8322
rect 81472 -8333 81477 -8284
rect 81711 -8293 81718 -8285
rect 81811 -8293 81818 -8285
rect 81638 -8327 81707 -8293
rect 81710 -8327 81751 -8293
rect 81822 -8327 81863 -8293
rect 82353 -8317 82394 -8283
rect 82449 -8317 82490 -8283
rect 82545 -8317 82586 -8283
rect 82641 -8317 82682 -8283
rect 82737 -8317 82778 -8283
rect 83762 -8324 83803 -8290
rect 83807 -8324 83814 -8279
rect 81472 -8367 81513 -8333
rect 82065 -8336 82072 -8328
rect 82165 -8336 82172 -8328
rect 81461 -8417 81468 -8406
rect 81472 -8417 81477 -8367
rect 81666 -8410 81707 -8376
rect 81711 -8410 81718 -8365
rect 81811 -8376 81818 -8365
rect 81992 -8370 82061 -8336
rect 82064 -8370 82105 -8336
rect 82176 -8370 82217 -8336
rect 82901 -8360 82942 -8326
rect 82997 -8360 83038 -8326
rect 83093 -8360 83134 -8326
rect 83189 -8360 83230 -8326
rect 83285 -8360 83326 -8326
rect 83381 -8360 83422 -8326
rect 83477 -8360 83518 -8326
rect 81822 -8410 81863 -8376
rect 82455 -8379 82462 -8371
rect 81472 -8451 81513 -8417
rect 81461 -8500 81468 -8489
rect 81472 -8500 81477 -8451
rect 81666 -8494 81707 -8460
rect 81711 -8494 81718 -8449
rect 81811 -8460 81818 -8449
rect 82020 -8453 82061 -8419
rect 82065 -8453 82072 -8408
rect 82165 -8419 82172 -8408
rect 82346 -8413 82387 -8379
rect 82410 -8413 82462 -8379
rect 82490 -8413 82531 -8379
rect 82176 -8453 82217 -8419
rect 81822 -8494 81863 -8460
rect 81472 -8534 81513 -8500
rect 81472 -8568 81477 -8534
rect 80122 -8740 80127 -8706
rect 80418 -8723 80459 -8689
rect 80463 -8723 80470 -8681
rect 80605 -8741 80617 -8673
rect 80646 -8707 80651 -8639
rect 80691 -8671 80696 -8603
rect 80725 -8637 80730 -8571
rect 81666 -8577 81707 -8543
rect 81711 -8577 81718 -8532
rect 81811 -8543 81818 -8532
rect 82020 -8537 82061 -8503
rect 82065 -8537 82072 -8492
rect 82165 -8503 82172 -8492
rect 82410 -8496 82451 -8462
rect 82455 -8496 82462 -8451
rect 82176 -8537 82217 -8503
rect 81822 -8577 81863 -8543
rect 80735 -8621 80776 -8587
rect 80936 -8666 80977 -8632
rect 80705 -8689 80712 -8681
rect 80716 -8723 80757 -8689
rect 80936 -8734 80977 -8700
rect 77869 -8906 77910 -8872
rect 77941 -8906 77982 -8872
rect 78013 -8906 78054 -8872
rect 78326 -8913 78367 -8879
rect 78371 -8913 78378 -8868
rect 78471 -8879 78478 -8868
rect 78482 -8913 78523 -8879
rect 79066 -8895 79107 -8861
rect 79111 -8895 79118 -8853
rect 76960 -8959 77442 -8925
rect 78294 -8949 78335 -8915
rect 78366 -8949 78407 -8915
rect 78680 -8956 78721 -8922
rect 78725 -8956 78732 -8911
rect 78825 -8922 78832 -8911
rect 79253 -8913 79265 -8845
rect 79294 -8879 79299 -8811
rect 79339 -8843 79344 -8775
rect 79373 -8809 79378 -8743
rect 80605 -8753 80612 -8741
rect 80985 -8750 80990 -8616
rect 79383 -8793 79424 -8759
rect 79586 -8838 79627 -8804
rect 79353 -8861 79360 -8853
rect 79364 -8895 79405 -8861
rect 79586 -8906 79627 -8872
rect 78836 -8956 78877 -8922
rect 76960 -8985 77429 -8959
rect 76964 -8993 77171 -8985
rect 76980 -9003 77155 -8993
rect 76706 -9140 76887 -9114
rect 76213 -9174 76254 -9140
rect 76309 -9174 76350 -9140
rect 76405 -9174 76446 -9140
rect 76501 -9174 76542 -9140
rect 76597 -9174 76638 -9140
rect 76693 -9174 76887 -9140
rect 76706 -9200 76887 -9174
rect 76906 -9174 77013 -9050
rect 77165 -9062 77171 -9051
rect 76784 -9870 76825 -9200
rect 76906 -9228 76915 -9174
rect 76591 -9936 76742 -9924
rect 76259 -9970 76742 -9936
rect 76591 -9971 76742 -9970
rect 76772 -9971 76825 -9870
rect 76918 -9971 76959 -9174
rect 76964 -9971 76970 -9174
rect 77176 -9971 77217 -9062
rect 77310 -9971 77351 -8985
rect 77563 -9002 77604 -8968
rect 77659 -9002 77700 -8968
rect 77755 -9002 77796 -8968
rect 77851 -9002 77892 -8968
rect 77947 -9002 77988 -8968
rect 78043 -9002 78084 -8968
rect 78139 -9002 78180 -8968
rect 78648 -8992 78689 -8958
rect 78720 -8992 78761 -8958
rect 79066 -8995 79107 -8961
rect 79111 -8995 79118 -8950
rect 79253 -9001 79260 -8913
rect 79635 -8922 79640 -8788
rect 79353 -8961 79360 -8950
rect 79669 -8956 79674 -8762
rect 79709 -8778 79716 -8767
rect 79705 -8809 79716 -8778
rect 80031 -8796 80072 -8762
rect 79364 -8995 79405 -8961
rect 78301 -9045 78342 -9011
rect 78397 -9045 78438 -9011
rect 78493 -9045 78534 -9011
rect 79002 -9035 79043 -9001
rect 79074 -9035 79115 -9001
rect 79146 -9035 79187 -9001
rect 79218 -9029 79260 -9001
rect 79564 -9025 79605 -8991
rect 79609 -9025 79616 -8980
rect 79705 -8992 79710 -8809
rect 79739 -8995 79744 -8812
rect 79218 -9035 79259 -9029
rect 78655 -9088 78696 -9054
rect 78751 -9088 78792 -9054
rect 78847 -9088 78888 -9054
rect 79751 -9076 79758 -8809
rect 80380 -8819 80773 -8753
rect 81019 -8784 81024 -8590
rect 81059 -8606 81066 -8595
rect 81055 -8637 81066 -8606
rect 81381 -8624 81422 -8590
rect 79767 -8860 79808 -8826
rect 80116 -8830 80133 -8819
rect 80116 -8832 80122 -8830
rect 79767 -8928 79808 -8894
rect 79819 -8995 79824 -8860
rect 80050 -8874 80122 -8832
rect 80178 -8874 80773 -8819
rect 80914 -8853 80955 -8819
rect 80959 -8853 80966 -8808
rect 81055 -8820 81060 -8637
rect 81089 -8823 81094 -8640
rect 80050 -8877 80773 -8874
rect 79853 -8980 79858 -8892
rect 79970 -8942 80011 -8908
rect 80015 -8942 80022 -8900
rect 79851 -8991 79858 -8980
rect 79853 -9025 79858 -8991
rect 79862 -9025 79903 -8991
rect 79970 -9042 80011 -9008
rect 80015 -9042 80022 -8997
rect 79863 -9078 79904 -9044
rect 79935 -9078 79976 -9044
rect 80007 -9078 80048 -9044
rect 79009 -9131 79050 -9097
rect 79105 -9131 79146 -9097
rect 79201 -9131 79242 -9097
rect 79297 -9131 79338 -9097
rect 79393 -9131 79434 -9097
rect 80050 -9114 80201 -8877
rect 80380 -8899 80773 -8877
rect 80304 -8925 80773 -8899
rect 81101 -8904 81108 -8637
rect 81117 -8688 81158 -8654
rect 81117 -8756 81158 -8722
rect 81169 -8823 81174 -8688
rect 81731 -8691 81772 -8657
rect 81783 -8718 81788 -8641
rect 81203 -8808 81208 -8720
rect 81320 -8770 81361 -8736
rect 81365 -8770 81372 -8728
rect 81465 -8740 81472 -8729
rect 81476 -8774 81517 -8740
rect 81817 -8752 81822 -8607
rect 82020 -8620 82061 -8586
rect 82065 -8620 82072 -8575
rect 82165 -8586 82172 -8575
rect 82410 -8580 82451 -8546
rect 82455 -8580 82462 -8535
rect 82176 -8620 82217 -8586
rect 82085 -8734 82126 -8700
rect 82137 -8761 82142 -8684
rect 81201 -8819 81208 -8808
rect 81670 -8813 81711 -8779
rect 81715 -8813 81722 -8771
rect 81815 -8779 81822 -8771
rect 81826 -8813 81867 -8779
rect 82171 -8795 82176 -8650
rect 82410 -8663 82451 -8629
rect 82455 -8663 82462 -8618
rect 82532 -8679 82537 -8363
rect 82555 -8379 82562 -8371
rect 82566 -8379 82571 -8363
rect 82566 -8413 82607 -8379
rect 82611 -8413 82618 -8371
rect 82555 -8462 82562 -8451
rect 82566 -8462 82571 -8413
rect 82566 -8496 82607 -8462
rect 82611 -8496 82618 -8451
rect 82555 -8546 82562 -8535
rect 82566 -8546 82571 -8496
rect 82566 -8580 82607 -8546
rect 82611 -8580 82618 -8535
rect 82555 -8629 82562 -8618
rect 82566 -8629 82571 -8580
rect 82566 -8663 82607 -8629
rect 82611 -8663 82618 -8618
rect 82555 -8697 82562 -8671
rect 82566 -8713 82571 -8663
rect 82475 -8777 82516 -8743
rect 81203 -8853 81208 -8819
rect 81212 -8853 81253 -8819
rect 81320 -8870 81361 -8836
rect 81365 -8870 81372 -8825
rect 81465 -8832 81472 -8821
rect 81476 -8866 81517 -8832
rect 82024 -8856 82065 -8822
rect 82069 -8856 82076 -8814
rect 82169 -8822 82176 -8814
rect 82180 -8856 82221 -8822
rect 82597 -8845 82604 -8697
rect 82620 -8713 82623 -8363
rect 82654 -8679 82657 -8363
rect 82711 -8379 82718 -8371
rect 82660 -8413 82701 -8379
rect 82722 -8413 82773 -8379
rect 83432 -8422 83437 -8406
rect 83455 -8422 83462 -8414
rect 83466 -8422 83471 -8406
rect 83762 -8408 83803 -8374
rect 83807 -8408 83814 -8363
rect 82711 -8462 82718 -8451
rect 82892 -8456 82933 -8422
rect 82964 -8456 83005 -8422
rect 83036 -8456 83077 -8422
rect 83180 -8456 83221 -8422
rect 83252 -8456 83365 -8422
rect 83396 -8456 83437 -8422
rect 82722 -8496 82763 -8462
rect 82711 -8546 82718 -8535
rect 83289 -8539 83330 -8505
rect 82722 -8580 82763 -8546
rect 82711 -8629 82718 -8618
rect 82722 -8663 82763 -8629
rect 82954 -8689 82995 -8655
rect 82999 -8689 83006 -8644
rect 83076 -8706 83081 -8588
rect 83099 -8655 83106 -8644
rect 83110 -8655 83115 -8622
rect 83146 -8655 83151 -8622
rect 83110 -8689 83151 -8655
rect 83155 -8689 83162 -8644
rect 83110 -8740 83115 -8689
rect 83146 -8740 83151 -8689
rect 83180 -8706 83185 -8589
rect 83289 -8623 83330 -8589
rect 83289 -8706 83330 -8672
rect 83432 -8706 83437 -8456
rect 83466 -8456 83507 -8422
rect 83455 -8505 83462 -8494
rect 83466 -8505 83471 -8456
rect 83762 -8491 83803 -8457
rect 83807 -8491 83814 -8446
rect 83466 -8539 83507 -8505
rect 83455 -8589 83462 -8578
rect 83466 -8589 83471 -8539
rect 83615 -8565 83724 -8499
rect 83884 -8507 83889 -8191
rect 83907 -8207 83914 -8199
rect 83918 -8207 83923 -8191
rect 83918 -8241 83959 -8207
rect 83963 -8241 83970 -8199
rect 83907 -8290 83914 -8279
rect 83918 -8290 83923 -8241
rect 83918 -8324 83959 -8290
rect 83963 -8324 83970 -8279
rect 83907 -8374 83914 -8363
rect 83918 -8374 83923 -8324
rect 83918 -8408 83959 -8374
rect 83963 -8408 83970 -8363
rect 83907 -8457 83914 -8446
rect 83918 -8457 83923 -8408
rect 83918 -8491 83959 -8457
rect 83963 -8491 83970 -8446
rect 83907 -8525 83914 -8499
rect 83918 -8541 83923 -8491
rect 83466 -8623 83507 -8589
rect 83827 -8605 83868 -8571
rect 83455 -8672 83462 -8661
rect 83466 -8672 83471 -8623
rect 83466 -8706 83507 -8672
rect 83949 -8673 83956 -8525
rect 83972 -8541 83975 -8191
rect 84006 -8507 84009 -8191
rect 84063 -8207 84070 -8199
rect 84012 -8241 84053 -8207
rect 84074 -8241 84125 -8207
rect 84989 -8231 85030 -8197
rect 85085 -8231 85126 -8197
rect 85181 -8231 85222 -8197
rect 87151 -8207 87158 -8199
rect 84782 -8250 84787 -8234
rect 84805 -8250 84812 -8242
rect 84816 -8250 84821 -8234
rect 84063 -8290 84070 -8279
rect 84242 -8284 84283 -8250
rect 84314 -8284 84355 -8250
rect 84386 -8284 84427 -8250
rect 84530 -8284 84571 -8250
rect 84602 -8284 84715 -8250
rect 84746 -8284 84787 -8250
rect 84074 -8324 84115 -8290
rect 84063 -8374 84070 -8363
rect 84639 -8367 84680 -8333
rect 84074 -8408 84115 -8374
rect 84063 -8457 84070 -8446
rect 84074 -8491 84115 -8457
rect 84304 -8517 84345 -8483
rect 84349 -8517 84356 -8472
rect 84426 -8534 84431 -8416
rect 84449 -8483 84456 -8472
rect 84460 -8483 84465 -8450
rect 84496 -8483 84501 -8450
rect 84460 -8517 84501 -8483
rect 84505 -8517 84512 -8472
rect 84460 -8568 84465 -8517
rect 84496 -8568 84501 -8517
rect 84530 -8534 84535 -8417
rect 84639 -8451 84680 -8417
rect 84639 -8534 84680 -8500
rect 84782 -8534 84787 -8284
rect 84816 -8284 84857 -8250
rect 85343 -8274 85384 -8240
rect 85439 -8274 85480 -8240
rect 85535 -8274 85576 -8240
rect 87042 -8241 87083 -8207
rect 87106 -8241 87158 -8207
rect 87186 -8241 87227 -8207
rect 84805 -8333 84812 -8322
rect 84816 -8333 84821 -8284
rect 85055 -8293 85062 -8285
rect 85155 -8293 85162 -8285
rect 84982 -8327 85051 -8293
rect 85054 -8327 85095 -8293
rect 85166 -8327 85207 -8293
rect 85697 -8317 85738 -8283
rect 85793 -8317 85834 -8283
rect 85889 -8317 85930 -8283
rect 85985 -8317 86026 -8283
rect 86081 -8317 86122 -8283
rect 87106 -8324 87147 -8290
rect 87151 -8324 87158 -8279
rect 84816 -8367 84857 -8333
rect 85409 -8336 85416 -8328
rect 85509 -8336 85516 -8328
rect 84805 -8417 84812 -8406
rect 84816 -8417 84821 -8367
rect 85010 -8410 85051 -8376
rect 85055 -8410 85062 -8365
rect 85155 -8376 85162 -8365
rect 85336 -8370 85405 -8336
rect 85408 -8370 85449 -8336
rect 85520 -8370 85561 -8336
rect 86245 -8360 86286 -8326
rect 86341 -8360 86382 -8326
rect 86437 -8360 86478 -8326
rect 86533 -8360 86574 -8326
rect 86629 -8360 86670 -8326
rect 86725 -8360 86766 -8326
rect 86821 -8360 86862 -8326
rect 85166 -8410 85207 -8376
rect 85799 -8379 85806 -8371
rect 84816 -8451 84857 -8417
rect 84805 -8500 84812 -8489
rect 84816 -8500 84821 -8451
rect 85010 -8494 85051 -8460
rect 85055 -8494 85062 -8449
rect 85155 -8460 85162 -8449
rect 85364 -8453 85405 -8419
rect 85409 -8453 85416 -8408
rect 85509 -8419 85516 -8408
rect 85690 -8413 85731 -8379
rect 85754 -8413 85806 -8379
rect 85834 -8413 85875 -8379
rect 85520 -8453 85561 -8419
rect 85166 -8494 85207 -8460
rect 84816 -8534 84857 -8500
rect 84816 -8568 84821 -8534
rect 83466 -8740 83471 -8706
rect 83762 -8723 83803 -8689
rect 83807 -8723 83814 -8681
rect 83949 -8741 83961 -8673
rect 83990 -8707 83995 -8639
rect 84035 -8671 84040 -8603
rect 84069 -8637 84074 -8571
rect 85010 -8577 85051 -8543
rect 85055 -8577 85062 -8532
rect 85155 -8543 85162 -8532
rect 85364 -8537 85405 -8503
rect 85409 -8537 85416 -8492
rect 85509 -8503 85516 -8492
rect 85754 -8496 85795 -8462
rect 85799 -8496 85806 -8451
rect 85520 -8537 85561 -8503
rect 85166 -8577 85207 -8543
rect 84079 -8621 84120 -8587
rect 84280 -8666 84321 -8632
rect 84049 -8689 84056 -8681
rect 84060 -8723 84101 -8689
rect 84280 -8734 84321 -8700
rect 81213 -8906 81254 -8872
rect 81285 -8906 81326 -8872
rect 81357 -8906 81398 -8872
rect 81670 -8913 81711 -8879
rect 81715 -8913 81722 -8868
rect 81815 -8879 81822 -8868
rect 81826 -8913 81867 -8879
rect 82410 -8895 82451 -8861
rect 82455 -8895 82462 -8853
rect 80304 -8959 80786 -8925
rect 81638 -8949 81679 -8915
rect 81710 -8949 81751 -8915
rect 82024 -8956 82065 -8922
rect 82069 -8956 82076 -8911
rect 82169 -8922 82176 -8911
rect 82597 -8913 82609 -8845
rect 82638 -8879 82643 -8811
rect 82683 -8843 82688 -8775
rect 82717 -8809 82722 -8743
rect 83949 -8753 83956 -8741
rect 84329 -8750 84334 -8616
rect 82727 -8793 82768 -8759
rect 82930 -8838 82971 -8804
rect 82697 -8861 82704 -8853
rect 82708 -8895 82749 -8861
rect 82930 -8906 82971 -8872
rect 82180 -8956 82221 -8922
rect 80304 -8985 80773 -8959
rect 80308 -8993 80515 -8985
rect 80324 -9003 80499 -8993
rect 80050 -9140 80231 -9114
rect 79557 -9174 79598 -9140
rect 79653 -9174 79694 -9140
rect 79749 -9174 79790 -9140
rect 79845 -9174 79886 -9140
rect 79941 -9174 79982 -9140
rect 80037 -9174 80231 -9140
rect 80050 -9200 80231 -9174
rect 80250 -9174 80357 -9050
rect 80509 -9062 80515 -9051
rect 80128 -9870 80169 -9200
rect 80250 -9228 80259 -9174
rect 79935 -9936 80086 -9924
rect 79603 -9970 80086 -9936
rect 79935 -9971 80086 -9970
rect 80116 -9971 80169 -9870
rect 80262 -9971 80303 -9174
rect 80308 -9971 80314 -9174
rect 80520 -9971 80561 -9062
rect 80654 -9971 80695 -8985
rect 80907 -9002 80948 -8968
rect 81003 -9002 81044 -8968
rect 81099 -9002 81140 -8968
rect 81195 -9002 81236 -8968
rect 81291 -9002 81332 -8968
rect 81387 -9002 81428 -8968
rect 81483 -9002 81524 -8968
rect 81992 -8992 82033 -8958
rect 82064 -8992 82105 -8958
rect 82410 -8995 82451 -8961
rect 82455 -8995 82462 -8950
rect 82597 -9001 82604 -8913
rect 82979 -8922 82984 -8788
rect 82697 -8961 82704 -8950
rect 83013 -8956 83018 -8762
rect 83053 -8778 83060 -8767
rect 83049 -8809 83060 -8778
rect 83375 -8796 83416 -8762
rect 82708 -8995 82749 -8961
rect 81645 -9045 81686 -9011
rect 81741 -9045 81782 -9011
rect 81837 -9045 81878 -9011
rect 82346 -9035 82387 -9001
rect 82418 -9035 82459 -9001
rect 82490 -9035 82531 -9001
rect 82562 -9029 82604 -9001
rect 82908 -9025 82949 -8991
rect 82953 -9025 82960 -8980
rect 83049 -8992 83054 -8809
rect 83083 -8995 83088 -8812
rect 82562 -9035 82603 -9029
rect 81999 -9088 82040 -9054
rect 82095 -9088 82136 -9054
rect 82191 -9088 82232 -9054
rect 83095 -9076 83102 -8809
rect 83724 -8819 84117 -8753
rect 84363 -8784 84368 -8590
rect 84403 -8606 84410 -8595
rect 84399 -8637 84410 -8606
rect 84725 -8624 84766 -8590
rect 83111 -8860 83152 -8826
rect 83460 -8830 83477 -8819
rect 83460 -8832 83466 -8830
rect 83111 -8928 83152 -8894
rect 83163 -8995 83168 -8860
rect 83394 -8874 83466 -8832
rect 83522 -8874 84117 -8819
rect 84258 -8853 84299 -8819
rect 84303 -8853 84310 -8808
rect 84399 -8820 84404 -8637
rect 84433 -8823 84438 -8640
rect 83394 -8877 84117 -8874
rect 83197 -8980 83202 -8892
rect 83314 -8942 83355 -8908
rect 83359 -8942 83366 -8900
rect 83195 -8991 83202 -8980
rect 83197 -9025 83202 -8991
rect 83206 -9025 83247 -8991
rect 83314 -9042 83355 -9008
rect 83359 -9042 83366 -8997
rect 83207 -9078 83248 -9044
rect 83279 -9078 83320 -9044
rect 83351 -9078 83392 -9044
rect 82353 -9131 82394 -9097
rect 82449 -9131 82490 -9097
rect 82545 -9131 82586 -9097
rect 82641 -9131 82682 -9097
rect 82737 -9131 82778 -9097
rect 83394 -9114 83545 -8877
rect 83724 -8899 84117 -8877
rect 83648 -8925 84117 -8899
rect 84445 -8904 84452 -8637
rect 84461 -8688 84502 -8654
rect 84461 -8756 84502 -8722
rect 84513 -8823 84518 -8688
rect 85075 -8691 85116 -8657
rect 85127 -8718 85132 -8641
rect 84547 -8808 84552 -8720
rect 84664 -8770 84705 -8736
rect 84709 -8770 84716 -8728
rect 84809 -8740 84816 -8729
rect 84820 -8774 84861 -8740
rect 85161 -8752 85166 -8607
rect 85364 -8620 85405 -8586
rect 85409 -8620 85416 -8575
rect 85509 -8586 85516 -8575
rect 85754 -8580 85795 -8546
rect 85799 -8580 85806 -8535
rect 85520 -8620 85561 -8586
rect 85429 -8734 85470 -8700
rect 85481 -8761 85486 -8684
rect 84545 -8819 84552 -8808
rect 85014 -8813 85055 -8779
rect 85059 -8813 85066 -8771
rect 85159 -8779 85166 -8771
rect 85170 -8813 85211 -8779
rect 85515 -8795 85520 -8650
rect 85754 -8663 85795 -8629
rect 85799 -8663 85806 -8618
rect 85876 -8679 85881 -8363
rect 85899 -8379 85906 -8371
rect 85910 -8379 85915 -8363
rect 85910 -8413 85951 -8379
rect 85955 -8413 85962 -8371
rect 85899 -8462 85906 -8451
rect 85910 -8462 85915 -8413
rect 85910 -8496 85951 -8462
rect 85955 -8496 85962 -8451
rect 85899 -8546 85906 -8535
rect 85910 -8546 85915 -8496
rect 85910 -8580 85951 -8546
rect 85955 -8580 85962 -8535
rect 85899 -8629 85906 -8618
rect 85910 -8629 85915 -8580
rect 85910 -8663 85951 -8629
rect 85955 -8663 85962 -8618
rect 85899 -8697 85906 -8671
rect 85910 -8713 85915 -8663
rect 85819 -8777 85860 -8743
rect 84547 -8853 84552 -8819
rect 84556 -8853 84597 -8819
rect 84664 -8870 84705 -8836
rect 84709 -8870 84716 -8825
rect 84809 -8832 84816 -8821
rect 84820 -8866 84861 -8832
rect 85368 -8856 85409 -8822
rect 85413 -8856 85420 -8814
rect 85513 -8822 85520 -8814
rect 85524 -8856 85565 -8822
rect 85941 -8845 85948 -8697
rect 85964 -8713 85967 -8363
rect 85998 -8679 86001 -8363
rect 86055 -8379 86062 -8371
rect 86004 -8413 86045 -8379
rect 86066 -8413 86117 -8379
rect 86776 -8422 86781 -8406
rect 86799 -8422 86806 -8414
rect 86810 -8422 86815 -8406
rect 87106 -8408 87147 -8374
rect 87151 -8408 87158 -8363
rect 86055 -8462 86062 -8451
rect 86236 -8456 86277 -8422
rect 86308 -8456 86349 -8422
rect 86380 -8456 86421 -8422
rect 86524 -8456 86565 -8422
rect 86596 -8456 86709 -8422
rect 86740 -8456 86781 -8422
rect 86066 -8496 86107 -8462
rect 86055 -8546 86062 -8535
rect 86633 -8539 86674 -8505
rect 86066 -8580 86107 -8546
rect 86055 -8629 86062 -8618
rect 86066 -8663 86107 -8629
rect 86298 -8689 86339 -8655
rect 86343 -8689 86350 -8644
rect 86420 -8706 86425 -8588
rect 86443 -8655 86450 -8644
rect 86454 -8655 86459 -8622
rect 86490 -8655 86495 -8622
rect 86454 -8689 86495 -8655
rect 86499 -8689 86506 -8644
rect 86454 -8740 86459 -8689
rect 86490 -8740 86495 -8689
rect 86524 -8706 86529 -8589
rect 86633 -8623 86674 -8589
rect 86633 -8706 86674 -8672
rect 86776 -8706 86781 -8456
rect 86810 -8456 86851 -8422
rect 86799 -8505 86806 -8494
rect 86810 -8505 86815 -8456
rect 87106 -8491 87147 -8457
rect 87151 -8491 87158 -8446
rect 86810 -8539 86851 -8505
rect 86799 -8589 86806 -8578
rect 86810 -8589 86815 -8539
rect 86959 -8565 87068 -8499
rect 87228 -8507 87233 -8191
rect 87251 -8207 87258 -8199
rect 87262 -8207 87267 -8191
rect 87262 -8241 87303 -8207
rect 87307 -8241 87314 -8199
rect 87251 -8290 87258 -8279
rect 87262 -8290 87267 -8241
rect 87262 -8324 87303 -8290
rect 87307 -8324 87314 -8279
rect 87251 -8374 87258 -8363
rect 87262 -8374 87267 -8324
rect 87262 -8408 87303 -8374
rect 87307 -8408 87314 -8363
rect 87251 -8457 87258 -8446
rect 87262 -8457 87267 -8408
rect 87262 -8491 87303 -8457
rect 87307 -8491 87314 -8446
rect 87251 -8525 87258 -8499
rect 87262 -8541 87267 -8491
rect 86810 -8623 86851 -8589
rect 87171 -8605 87212 -8571
rect 86799 -8672 86806 -8661
rect 86810 -8672 86815 -8623
rect 86810 -8706 86851 -8672
rect 87293 -8673 87300 -8525
rect 87316 -8541 87319 -8191
rect 87350 -8507 87353 -8191
rect 87407 -8207 87414 -8199
rect 87356 -8241 87397 -8207
rect 87418 -8241 87469 -8207
rect 88333 -8231 88374 -8197
rect 88429 -8231 88470 -8197
rect 88525 -8231 88566 -8197
rect 90495 -8207 90502 -8199
rect 88126 -8250 88131 -8234
rect 88149 -8250 88156 -8242
rect 88160 -8250 88165 -8234
rect 87407 -8290 87414 -8279
rect 87586 -8284 87627 -8250
rect 87658 -8284 87699 -8250
rect 87730 -8284 87771 -8250
rect 87874 -8284 87915 -8250
rect 87946 -8284 88059 -8250
rect 88090 -8284 88131 -8250
rect 87418 -8324 87459 -8290
rect 87407 -8374 87414 -8363
rect 87983 -8367 88024 -8333
rect 87418 -8408 87459 -8374
rect 87407 -8457 87414 -8446
rect 87418 -8491 87459 -8457
rect 87648 -8517 87689 -8483
rect 87693 -8517 87700 -8472
rect 87770 -8534 87775 -8416
rect 87793 -8483 87800 -8472
rect 87804 -8483 87809 -8450
rect 87840 -8483 87845 -8450
rect 87804 -8517 87845 -8483
rect 87849 -8517 87856 -8472
rect 87804 -8568 87809 -8517
rect 87840 -8568 87845 -8517
rect 87874 -8534 87879 -8417
rect 87983 -8451 88024 -8417
rect 87983 -8534 88024 -8500
rect 88126 -8534 88131 -8284
rect 88160 -8284 88201 -8250
rect 88687 -8274 88728 -8240
rect 88783 -8274 88824 -8240
rect 88879 -8274 88920 -8240
rect 90386 -8241 90427 -8207
rect 90450 -8241 90502 -8207
rect 90530 -8241 90571 -8207
rect 88149 -8333 88156 -8322
rect 88160 -8333 88165 -8284
rect 88399 -8293 88406 -8285
rect 88499 -8293 88506 -8285
rect 88326 -8327 88395 -8293
rect 88398 -8327 88439 -8293
rect 88510 -8327 88551 -8293
rect 89041 -8317 89082 -8283
rect 89137 -8317 89178 -8283
rect 89233 -8317 89274 -8283
rect 89329 -8317 89370 -8283
rect 89425 -8317 89466 -8283
rect 90450 -8324 90491 -8290
rect 90495 -8324 90502 -8279
rect 88160 -8367 88201 -8333
rect 88753 -8336 88760 -8328
rect 88853 -8336 88860 -8328
rect 88149 -8417 88156 -8406
rect 88160 -8417 88165 -8367
rect 88354 -8410 88395 -8376
rect 88399 -8410 88406 -8365
rect 88499 -8376 88506 -8365
rect 88680 -8370 88749 -8336
rect 88752 -8370 88793 -8336
rect 88864 -8370 88905 -8336
rect 89589 -8360 89630 -8326
rect 89685 -8360 89726 -8326
rect 89781 -8360 89822 -8326
rect 89877 -8360 89918 -8326
rect 89973 -8360 90014 -8326
rect 90069 -8360 90110 -8326
rect 90165 -8360 90206 -8326
rect 88510 -8410 88551 -8376
rect 89143 -8379 89150 -8371
rect 88160 -8451 88201 -8417
rect 88149 -8500 88156 -8489
rect 88160 -8500 88165 -8451
rect 88354 -8494 88395 -8460
rect 88399 -8494 88406 -8449
rect 88499 -8460 88506 -8449
rect 88708 -8453 88749 -8419
rect 88753 -8453 88760 -8408
rect 88853 -8419 88860 -8408
rect 89034 -8413 89075 -8379
rect 89098 -8413 89150 -8379
rect 89178 -8413 89219 -8379
rect 88864 -8453 88905 -8419
rect 88510 -8494 88551 -8460
rect 88160 -8534 88201 -8500
rect 88160 -8568 88165 -8534
rect 86810 -8740 86815 -8706
rect 87106 -8723 87147 -8689
rect 87151 -8723 87158 -8681
rect 87293 -8741 87305 -8673
rect 87334 -8707 87339 -8639
rect 87379 -8671 87384 -8603
rect 87413 -8637 87418 -8571
rect 88354 -8577 88395 -8543
rect 88399 -8577 88406 -8532
rect 88499 -8543 88506 -8532
rect 88708 -8537 88749 -8503
rect 88753 -8537 88760 -8492
rect 88853 -8503 88860 -8492
rect 89098 -8496 89139 -8462
rect 89143 -8496 89150 -8451
rect 88864 -8537 88905 -8503
rect 88510 -8577 88551 -8543
rect 87423 -8621 87464 -8587
rect 87624 -8666 87665 -8632
rect 87393 -8689 87400 -8681
rect 87404 -8723 87445 -8689
rect 87624 -8734 87665 -8700
rect 84557 -8906 84598 -8872
rect 84629 -8906 84670 -8872
rect 84701 -8906 84742 -8872
rect 85014 -8913 85055 -8879
rect 85059 -8913 85066 -8868
rect 85159 -8879 85166 -8868
rect 85170 -8913 85211 -8879
rect 85754 -8895 85795 -8861
rect 85799 -8895 85806 -8853
rect 83648 -8959 84130 -8925
rect 84982 -8949 85023 -8915
rect 85054 -8949 85095 -8915
rect 85368 -8956 85409 -8922
rect 85413 -8956 85420 -8911
rect 85513 -8922 85520 -8911
rect 85941 -8913 85953 -8845
rect 85982 -8879 85987 -8811
rect 86027 -8843 86032 -8775
rect 86061 -8809 86066 -8743
rect 87293 -8753 87300 -8741
rect 87673 -8750 87678 -8616
rect 86071 -8793 86112 -8759
rect 86274 -8838 86315 -8804
rect 86041 -8861 86048 -8853
rect 86052 -8895 86093 -8861
rect 86274 -8906 86315 -8872
rect 85524 -8956 85565 -8922
rect 83648 -8985 84117 -8959
rect 83652 -8993 83859 -8985
rect 83668 -9003 83843 -8993
rect 83394 -9140 83575 -9114
rect 82901 -9174 82942 -9140
rect 82997 -9174 83038 -9140
rect 83093 -9174 83134 -9140
rect 83189 -9174 83230 -9140
rect 83285 -9174 83326 -9140
rect 83381 -9174 83575 -9140
rect 83394 -9200 83575 -9174
rect 83594 -9174 83701 -9050
rect 83853 -9062 83859 -9051
rect 83472 -9870 83513 -9200
rect 83594 -9228 83603 -9174
rect 83279 -9936 83430 -9924
rect 82947 -9970 83430 -9936
rect 83279 -9971 83430 -9970
rect 83460 -9971 83513 -9870
rect 83606 -9971 83647 -9174
rect 83652 -9971 83658 -9174
rect 83864 -9971 83905 -9062
rect 83998 -9971 84039 -8985
rect 84251 -9002 84292 -8968
rect 84347 -9002 84388 -8968
rect 84443 -9002 84484 -8968
rect 84539 -9002 84580 -8968
rect 84635 -9002 84676 -8968
rect 84731 -9002 84772 -8968
rect 84827 -9002 84868 -8968
rect 85336 -8992 85377 -8958
rect 85408 -8992 85449 -8958
rect 85754 -8995 85795 -8961
rect 85799 -8995 85806 -8950
rect 85941 -9001 85948 -8913
rect 86323 -8922 86328 -8788
rect 86041 -8961 86048 -8950
rect 86357 -8956 86362 -8762
rect 86397 -8778 86404 -8767
rect 86393 -8809 86404 -8778
rect 86719 -8796 86760 -8762
rect 86052 -8995 86093 -8961
rect 84989 -9045 85030 -9011
rect 85085 -9045 85126 -9011
rect 85181 -9045 85222 -9011
rect 85690 -9035 85731 -9001
rect 85762 -9035 85803 -9001
rect 85834 -9035 85875 -9001
rect 85906 -9029 85948 -9001
rect 86252 -9025 86293 -8991
rect 86297 -9025 86304 -8980
rect 86393 -8992 86398 -8809
rect 86427 -8995 86432 -8812
rect 85906 -9035 85947 -9029
rect 85343 -9088 85384 -9054
rect 85439 -9088 85480 -9054
rect 85535 -9088 85576 -9054
rect 86439 -9076 86446 -8809
rect 87068 -8819 87461 -8753
rect 87707 -8784 87712 -8590
rect 87747 -8606 87754 -8595
rect 87743 -8637 87754 -8606
rect 88069 -8624 88110 -8590
rect 86455 -8860 86496 -8826
rect 86804 -8830 86821 -8819
rect 86804 -8832 86810 -8830
rect 86455 -8928 86496 -8894
rect 86507 -8995 86512 -8860
rect 86738 -8874 86810 -8832
rect 86866 -8874 87461 -8819
rect 87602 -8853 87643 -8819
rect 87647 -8853 87654 -8808
rect 87743 -8820 87748 -8637
rect 87777 -8823 87782 -8640
rect 86738 -8877 87461 -8874
rect 86541 -8980 86546 -8892
rect 86658 -8942 86699 -8908
rect 86703 -8942 86710 -8900
rect 86539 -8991 86546 -8980
rect 86541 -9025 86546 -8991
rect 86550 -9025 86591 -8991
rect 86658 -9042 86699 -9008
rect 86703 -9042 86710 -8997
rect 86551 -9078 86592 -9044
rect 86623 -9078 86664 -9044
rect 86695 -9078 86736 -9044
rect 85697 -9131 85738 -9097
rect 85793 -9131 85834 -9097
rect 85889 -9131 85930 -9097
rect 85985 -9131 86026 -9097
rect 86081 -9131 86122 -9097
rect 86738 -9114 86889 -8877
rect 87068 -8899 87461 -8877
rect 86992 -8925 87461 -8899
rect 87789 -8904 87796 -8637
rect 87805 -8688 87846 -8654
rect 87805 -8756 87846 -8722
rect 87857 -8823 87862 -8688
rect 88419 -8691 88460 -8657
rect 88471 -8718 88476 -8641
rect 87891 -8808 87896 -8720
rect 88008 -8770 88049 -8736
rect 88053 -8770 88060 -8728
rect 88153 -8740 88160 -8729
rect 88164 -8774 88205 -8740
rect 88505 -8752 88510 -8607
rect 88708 -8620 88749 -8586
rect 88753 -8620 88760 -8575
rect 88853 -8586 88860 -8575
rect 89098 -8580 89139 -8546
rect 89143 -8580 89150 -8535
rect 88864 -8620 88905 -8586
rect 88773 -8734 88814 -8700
rect 88825 -8761 88830 -8684
rect 87889 -8819 87896 -8808
rect 88358 -8813 88399 -8779
rect 88403 -8813 88410 -8771
rect 88503 -8779 88510 -8771
rect 88514 -8813 88555 -8779
rect 88859 -8795 88864 -8650
rect 89098 -8663 89139 -8629
rect 89143 -8663 89150 -8618
rect 89220 -8679 89225 -8363
rect 89243 -8379 89250 -8371
rect 89254 -8379 89259 -8363
rect 89254 -8413 89295 -8379
rect 89299 -8413 89306 -8371
rect 89243 -8462 89250 -8451
rect 89254 -8462 89259 -8413
rect 89254 -8496 89295 -8462
rect 89299 -8496 89306 -8451
rect 89243 -8546 89250 -8535
rect 89254 -8546 89259 -8496
rect 89254 -8580 89295 -8546
rect 89299 -8580 89306 -8535
rect 89243 -8629 89250 -8618
rect 89254 -8629 89259 -8580
rect 89254 -8663 89295 -8629
rect 89299 -8663 89306 -8618
rect 89243 -8697 89250 -8671
rect 89254 -8713 89259 -8663
rect 89163 -8777 89204 -8743
rect 87891 -8853 87896 -8819
rect 87900 -8853 87941 -8819
rect 88008 -8870 88049 -8836
rect 88053 -8870 88060 -8825
rect 88153 -8832 88160 -8821
rect 88164 -8866 88205 -8832
rect 88712 -8856 88753 -8822
rect 88757 -8856 88764 -8814
rect 88857 -8822 88864 -8814
rect 88868 -8856 88909 -8822
rect 89285 -8845 89292 -8697
rect 89308 -8713 89311 -8363
rect 89342 -8679 89345 -8363
rect 89399 -8379 89406 -8371
rect 89348 -8413 89389 -8379
rect 89410 -8413 89461 -8379
rect 90120 -8422 90125 -8406
rect 90143 -8422 90150 -8414
rect 90154 -8422 90159 -8406
rect 90450 -8408 90491 -8374
rect 90495 -8408 90502 -8363
rect 89399 -8462 89406 -8451
rect 89580 -8456 89621 -8422
rect 89652 -8456 89693 -8422
rect 89724 -8456 89765 -8422
rect 89868 -8456 89909 -8422
rect 89940 -8456 90053 -8422
rect 90084 -8456 90125 -8422
rect 89410 -8496 89451 -8462
rect 89399 -8546 89406 -8535
rect 89977 -8539 90018 -8505
rect 89410 -8580 89451 -8546
rect 89399 -8629 89406 -8618
rect 89410 -8663 89451 -8629
rect 89642 -8689 89683 -8655
rect 89687 -8689 89694 -8644
rect 89764 -8706 89769 -8588
rect 89787 -8655 89794 -8644
rect 89798 -8655 89803 -8622
rect 89834 -8655 89839 -8622
rect 89798 -8689 89839 -8655
rect 89843 -8689 89850 -8644
rect 89798 -8740 89803 -8689
rect 89834 -8740 89839 -8689
rect 89868 -8706 89873 -8589
rect 89977 -8623 90018 -8589
rect 89977 -8706 90018 -8672
rect 90120 -8706 90125 -8456
rect 90154 -8456 90195 -8422
rect 90143 -8505 90150 -8494
rect 90154 -8505 90159 -8456
rect 90450 -8491 90491 -8457
rect 90495 -8491 90502 -8446
rect 90154 -8539 90195 -8505
rect 90143 -8589 90150 -8578
rect 90154 -8589 90159 -8539
rect 90303 -8565 90412 -8499
rect 90572 -8507 90577 -8191
rect 90595 -8207 90602 -8199
rect 90606 -8207 90611 -8191
rect 90606 -8241 90647 -8207
rect 90651 -8241 90658 -8199
rect 90595 -8290 90602 -8279
rect 90606 -8290 90611 -8241
rect 90606 -8324 90647 -8290
rect 90651 -8324 90658 -8279
rect 90595 -8374 90602 -8363
rect 90606 -8374 90611 -8324
rect 90606 -8408 90647 -8374
rect 90651 -8408 90658 -8363
rect 90595 -8457 90602 -8446
rect 90606 -8457 90611 -8408
rect 90606 -8491 90647 -8457
rect 90651 -8491 90658 -8446
rect 90595 -8525 90602 -8499
rect 90606 -8541 90611 -8491
rect 90154 -8623 90195 -8589
rect 90515 -8605 90556 -8571
rect 90143 -8672 90150 -8661
rect 90154 -8672 90159 -8623
rect 90154 -8706 90195 -8672
rect 90637 -8673 90644 -8525
rect 90660 -8541 90663 -8191
rect 90694 -8507 90697 -8191
rect 90751 -8207 90758 -8199
rect 90700 -8241 90741 -8207
rect 90762 -8241 90813 -8207
rect 91677 -8231 91718 -8197
rect 91773 -8231 91814 -8197
rect 91869 -8231 91910 -8197
rect 93839 -8207 93846 -8199
rect 91470 -8250 91475 -8234
rect 91493 -8250 91500 -8242
rect 91504 -8250 91509 -8234
rect 90751 -8290 90758 -8279
rect 90930 -8284 90971 -8250
rect 91002 -8284 91043 -8250
rect 91074 -8284 91115 -8250
rect 91218 -8284 91259 -8250
rect 91290 -8284 91403 -8250
rect 91434 -8284 91475 -8250
rect 90762 -8324 90803 -8290
rect 90751 -8374 90758 -8363
rect 91327 -8367 91368 -8333
rect 90762 -8408 90803 -8374
rect 90751 -8457 90758 -8446
rect 90762 -8491 90803 -8457
rect 90992 -8517 91033 -8483
rect 91037 -8517 91044 -8472
rect 91114 -8534 91119 -8416
rect 91137 -8483 91144 -8472
rect 91148 -8483 91153 -8450
rect 91184 -8483 91189 -8450
rect 91148 -8517 91189 -8483
rect 91193 -8517 91200 -8472
rect 91148 -8568 91153 -8517
rect 91184 -8568 91189 -8517
rect 91218 -8534 91223 -8417
rect 91327 -8451 91368 -8417
rect 91327 -8534 91368 -8500
rect 91470 -8534 91475 -8284
rect 91504 -8284 91545 -8250
rect 92031 -8274 92072 -8240
rect 92127 -8274 92168 -8240
rect 92223 -8274 92264 -8240
rect 93730 -8241 93771 -8207
rect 93794 -8241 93846 -8207
rect 93874 -8241 93915 -8207
rect 91493 -8333 91500 -8322
rect 91504 -8333 91509 -8284
rect 91743 -8293 91750 -8285
rect 91843 -8293 91850 -8285
rect 91670 -8327 91739 -8293
rect 91742 -8327 91783 -8293
rect 91854 -8327 91895 -8293
rect 92385 -8317 92426 -8283
rect 92481 -8317 92522 -8283
rect 92577 -8317 92618 -8283
rect 92673 -8317 92714 -8283
rect 92769 -8317 92810 -8283
rect 93794 -8324 93835 -8290
rect 93839 -8324 93846 -8279
rect 91504 -8367 91545 -8333
rect 92097 -8336 92104 -8328
rect 92197 -8336 92204 -8328
rect 91493 -8417 91500 -8406
rect 91504 -8417 91509 -8367
rect 91698 -8410 91739 -8376
rect 91743 -8410 91750 -8365
rect 91843 -8376 91850 -8365
rect 92024 -8370 92093 -8336
rect 92096 -8370 92137 -8336
rect 92208 -8370 92249 -8336
rect 92933 -8360 92974 -8326
rect 93029 -8360 93070 -8326
rect 93125 -8360 93166 -8326
rect 93221 -8360 93262 -8326
rect 93317 -8360 93358 -8326
rect 93413 -8360 93454 -8326
rect 93509 -8360 93550 -8326
rect 91854 -8410 91895 -8376
rect 92487 -8379 92494 -8371
rect 91504 -8451 91545 -8417
rect 91493 -8500 91500 -8489
rect 91504 -8500 91509 -8451
rect 91698 -8494 91739 -8460
rect 91743 -8494 91750 -8449
rect 91843 -8460 91850 -8449
rect 92052 -8453 92093 -8419
rect 92097 -8453 92104 -8408
rect 92197 -8419 92204 -8408
rect 92378 -8413 92419 -8379
rect 92442 -8413 92494 -8379
rect 92522 -8413 92563 -8379
rect 92208 -8453 92249 -8419
rect 91854 -8494 91895 -8460
rect 91504 -8534 91545 -8500
rect 91504 -8568 91509 -8534
rect 90154 -8740 90159 -8706
rect 90450 -8723 90491 -8689
rect 90495 -8723 90502 -8681
rect 90637 -8741 90649 -8673
rect 90678 -8707 90683 -8639
rect 90723 -8671 90728 -8603
rect 90757 -8637 90762 -8571
rect 91698 -8577 91739 -8543
rect 91743 -8577 91750 -8532
rect 91843 -8543 91850 -8532
rect 92052 -8537 92093 -8503
rect 92097 -8537 92104 -8492
rect 92197 -8503 92204 -8492
rect 92442 -8496 92483 -8462
rect 92487 -8496 92494 -8451
rect 92208 -8537 92249 -8503
rect 91854 -8577 91895 -8543
rect 90767 -8621 90808 -8587
rect 90968 -8666 91009 -8632
rect 90737 -8689 90744 -8681
rect 90748 -8723 90789 -8689
rect 90968 -8734 91009 -8700
rect 87901 -8906 87942 -8872
rect 87973 -8906 88014 -8872
rect 88045 -8906 88086 -8872
rect 88358 -8913 88399 -8879
rect 88403 -8913 88410 -8868
rect 88503 -8879 88510 -8868
rect 88514 -8913 88555 -8879
rect 89098 -8895 89139 -8861
rect 89143 -8895 89150 -8853
rect 86992 -8959 87474 -8925
rect 88326 -8949 88367 -8915
rect 88398 -8949 88439 -8915
rect 88712 -8956 88753 -8922
rect 88757 -8956 88764 -8911
rect 88857 -8922 88864 -8911
rect 89285 -8913 89297 -8845
rect 89326 -8879 89331 -8811
rect 89371 -8843 89376 -8775
rect 89405 -8809 89410 -8743
rect 90637 -8753 90644 -8741
rect 91017 -8750 91022 -8616
rect 89415 -8793 89456 -8759
rect 89618 -8838 89659 -8804
rect 89385 -8861 89392 -8853
rect 89396 -8895 89437 -8861
rect 89618 -8906 89659 -8872
rect 88868 -8956 88909 -8922
rect 86992 -8985 87461 -8959
rect 86996 -8993 87203 -8985
rect 87012 -9003 87187 -8993
rect 86738 -9140 86919 -9114
rect 86245 -9174 86286 -9140
rect 86341 -9174 86382 -9140
rect 86437 -9174 86478 -9140
rect 86533 -9174 86574 -9140
rect 86629 -9174 86670 -9140
rect 86725 -9174 86919 -9140
rect 86738 -9200 86919 -9174
rect 86938 -9174 87045 -9050
rect 87197 -9062 87203 -9051
rect 86816 -9870 86857 -9200
rect 86938 -9228 86947 -9174
rect 86623 -9936 86774 -9924
rect 86291 -9970 86774 -9936
rect 86623 -9971 86774 -9970
rect 86804 -9971 86857 -9870
rect 86950 -9971 86991 -9174
rect 86996 -9971 87002 -9174
rect 87208 -9971 87249 -9062
rect 87342 -9971 87383 -8985
rect 87595 -9002 87636 -8968
rect 87691 -9002 87732 -8968
rect 87787 -9002 87828 -8968
rect 87883 -9002 87924 -8968
rect 87979 -9002 88020 -8968
rect 88075 -9002 88116 -8968
rect 88171 -9002 88212 -8968
rect 88680 -8992 88721 -8958
rect 88752 -8992 88793 -8958
rect 89098 -8995 89139 -8961
rect 89143 -8995 89150 -8950
rect 89285 -9001 89292 -8913
rect 89667 -8922 89672 -8788
rect 89385 -8961 89392 -8950
rect 89701 -8956 89706 -8762
rect 89741 -8778 89748 -8767
rect 89737 -8809 89748 -8778
rect 90063 -8796 90104 -8762
rect 89396 -8995 89437 -8961
rect 88333 -9045 88374 -9011
rect 88429 -9045 88470 -9011
rect 88525 -9045 88566 -9011
rect 89034 -9035 89075 -9001
rect 89106 -9035 89147 -9001
rect 89178 -9035 89219 -9001
rect 89250 -9029 89292 -9001
rect 89596 -9025 89637 -8991
rect 89641 -9025 89648 -8980
rect 89737 -8992 89742 -8809
rect 89771 -8995 89776 -8812
rect 89250 -9035 89291 -9029
rect 88687 -9088 88728 -9054
rect 88783 -9088 88824 -9054
rect 88879 -9088 88920 -9054
rect 89783 -9076 89790 -8809
rect 90412 -8819 90805 -8753
rect 91051 -8784 91056 -8590
rect 91091 -8606 91098 -8595
rect 91087 -8637 91098 -8606
rect 91413 -8624 91454 -8590
rect 89799 -8860 89840 -8826
rect 90148 -8830 90165 -8819
rect 90148 -8832 90154 -8830
rect 89799 -8928 89840 -8894
rect 89851 -8995 89856 -8860
rect 90082 -8874 90154 -8832
rect 90210 -8874 90805 -8819
rect 90946 -8853 90987 -8819
rect 90991 -8853 90998 -8808
rect 91087 -8820 91092 -8637
rect 91121 -8823 91126 -8640
rect 90082 -8877 90805 -8874
rect 89885 -8980 89890 -8892
rect 90002 -8942 90043 -8908
rect 90047 -8942 90054 -8900
rect 89883 -8991 89890 -8980
rect 89885 -9025 89890 -8991
rect 89894 -9025 89935 -8991
rect 90002 -9042 90043 -9008
rect 90047 -9042 90054 -8997
rect 89895 -9078 89936 -9044
rect 89967 -9078 90008 -9044
rect 90039 -9078 90080 -9044
rect 89041 -9131 89082 -9097
rect 89137 -9131 89178 -9097
rect 89233 -9131 89274 -9097
rect 89329 -9131 89370 -9097
rect 89425 -9131 89466 -9097
rect 90082 -9114 90233 -8877
rect 90412 -8899 90805 -8877
rect 90336 -8925 90805 -8899
rect 91133 -8904 91140 -8637
rect 91149 -8688 91190 -8654
rect 91149 -8756 91190 -8722
rect 91201 -8823 91206 -8688
rect 91763 -8691 91804 -8657
rect 91815 -8718 91820 -8641
rect 91235 -8808 91240 -8720
rect 91352 -8770 91393 -8736
rect 91397 -8770 91404 -8728
rect 91497 -8740 91504 -8729
rect 91508 -8774 91549 -8740
rect 91849 -8752 91854 -8607
rect 92052 -8620 92093 -8586
rect 92097 -8620 92104 -8575
rect 92197 -8586 92204 -8575
rect 92442 -8580 92483 -8546
rect 92487 -8580 92494 -8535
rect 92208 -8620 92249 -8586
rect 92117 -8734 92158 -8700
rect 92169 -8761 92174 -8684
rect 91233 -8819 91240 -8808
rect 91702 -8813 91743 -8779
rect 91747 -8813 91754 -8771
rect 91847 -8779 91854 -8771
rect 91858 -8813 91899 -8779
rect 92203 -8795 92208 -8650
rect 92442 -8663 92483 -8629
rect 92487 -8663 92494 -8618
rect 92564 -8679 92569 -8363
rect 92587 -8379 92594 -8371
rect 92598 -8379 92603 -8363
rect 92598 -8413 92639 -8379
rect 92643 -8413 92650 -8371
rect 92587 -8462 92594 -8451
rect 92598 -8462 92603 -8413
rect 92598 -8496 92639 -8462
rect 92643 -8496 92650 -8451
rect 92587 -8546 92594 -8535
rect 92598 -8546 92603 -8496
rect 92598 -8580 92639 -8546
rect 92643 -8580 92650 -8535
rect 92587 -8629 92594 -8618
rect 92598 -8629 92603 -8580
rect 92598 -8663 92639 -8629
rect 92643 -8663 92650 -8618
rect 92587 -8697 92594 -8671
rect 92598 -8713 92603 -8663
rect 92507 -8777 92548 -8743
rect 91235 -8853 91240 -8819
rect 91244 -8853 91285 -8819
rect 91352 -8870 91393 -8836
rect 91397 -8870 91404 -8825
rect 91497 -8832 91504 -8821
rect 91508 -8866 91549 -8832
rect 92056 -8856 92097 -8822
rect 92101 -8856 92108 -8814
rect 92201 -8822 92208 -8814
rect 92212 -8856 92253 -8822
rect 92629 -8845 92636 -8697
rect 92652 -8713 92655 -8363
rect 92686 -8679 92689 -8363
rect 92743 -8379 92750 -8371
rect 92692 -8413 92733 -8379
rect 92754 -8413 92805 -8379
rect 93464 -8422 93469 -8406
rect 93487 -8422 93494 -8414
rect 93498 -8422 93503 -8406
rect 93794 -8408 93835 -8374
rect 93839 -8408 93846 -8363
rect 92743 -8462 92750 -8451
rect 92924 -8456 92965 -8422
rect 92996 -8456 93037 -8422
rect 93068 -8456 93109 -8422
rect 93212 -8456 93253 -8422
rect 93284 -8456 93397 -8422
rect 93428 -8456 93469 -8422
rect 92754 -8496 92795 -8462
rect 92743 -8546 92750 -8535
rect 93321 -8539 93362 -8505
rect 92754 -8580 92795 -8546
rect 92743 -8629 92750 -8618
rect 92754 -8663 92795 -8629
rect 92986 -8689 93027 -8655
rect 93031 -8689 93038 -8644
rect 93108 -8706 93113 -8588
rect 93131 -8655 93138 -8644
rect 93142 -8655 93147 -8622
rect 93178 -8655 93183 -8622
rect 93142 -8689 93183 -8655
rect 93187 -8689 93194 -8644
rect 93142 -8740 93147 -8689
rect 93178 -8740 93183 -8689
rect 93212 -8706 93217 -8589
rect 93321 -8623 93362 -8589
rect 93321 -8706 93362 -8672
rect 93464 -8706 93469 -8456
rect 93498 -8456 93539 -8422
rect 93487 -8505 93494 -8494
rect 93498 -8505 93503 -8456
rect 93794 -8491 93835 -8457
rect 93839 -8491 93846 -8446
rect 93498 -8539 93539 -8505
rect 93487 -8589 93494 -8578
rect 93498 -8589 93503 -8539
rect 93647 -8565 93756 -8499
rect 93916 -8507 93921 -8191
rect 93939 -8207 93946 -8199
rect 93950 -8207 93955 -8191
rect 93950 -8241 93991 -8207
rect 93995 -8241 94002 -8199
rect 93939 -8290 93946 -8279
rect 93950 -8290 93955 -8241
rect 93950 -8324 93991 -8290
rect 93995 -8324 94002 -8279
rect 93939 -8374 93946 -8363
rect 93950 -8374 93955 -8324
rect 93950 -8408 93991 -8374
rect 93995 -8408 94002 -8363
rect 93939 -8457 93946 -8446
rect 93950 -8457 93955 -8408
rect 93950 -8491 93991 -8457
rect 93995 -8491 94002 -8446
rect 93939 -8525 93946 -8499
rect 93950 -8541 93955 -8491
rect 93498 -8623 93539 -8589
rect 93859 -8605 93900 -8571
rect 93487 -8672 93494 -8661
rect 93498 -8672 93503 -8623
rect 93498 -8706 93539 -8672
rect 93981 -8673 93988 -8525
rect 94004 -8541 94007 -8191
rect 94038 -8507 94041 -8191
rect 94095 -8207 94102 -8199
rect 94044 -8241 94085 -8207
rect 94106 -8241 94157 -8207
rect 95021 -8231 95062 -8197
rect 95117 -8231 95158 -8197
rect 95213 -8231 95254 -8197
rect 97183 -8207 97190 -8199
rect 94814 -8250 94819 -8234
rect 94837 -8250 94844 -8242
rect 94848 -8250 94853 -8234
rect 94095 -8290 94102 -8279
rect 94274 -8284 94315 -8250
rect 94346 -8284 94387 -8250
rect 94418 -8284 94459 -8250
rect 94562 -8284 94603 -8250
rect 94634 -8284 94747 -8250
rect 94778 -8284 94819 -8250
rect 94106 -8324 94147 -8290
rect 94095 -8374 94102 -8363
rect 94671 -8367 94712 -8333
rect 94106 -8408 94147 -8374
rect 94095 -8457 94102 -8446
rect 94106 -8491 94147 -8457
rect 94336 -8517 94377 -8483
rect 94381 -8517 94388 -8472
rect 94458 -8534 94463 -8416
rect 94481 -8483 94488 -8472
rect 94492 -8483 94497 -8450
rect 94528 -8483 94533 -8450
rect 94492 -8517 94533 -8483
rect 94537 -8517 94544 -8472
rect 94492 -8568 94497 -8517
rect 94528 -8568 94533 -8517
rect 94562 -8534 94567 -8417
rect 94671 -8451 94712 -8417
rect 94671 -8534 94712 -8500
rect 94814 -8534 94819 -8284
rect 94848 -8284 94889 -8250
rect 95375 -8274 95416 -8240
rect 95471 -8274 95512 -8240
rect 95567 -8274 95608 -8240
rect 97074 -8241 97115 -8207
rect 97138 -8241 97190 -8207
rect 97218 -8241 97259 -8207
rect 94837 -8333 94844 -8322
rect 94848 -8333 94853 -8284
rect 95087 -8293 95094 -8285
rect 95187 -8293 95194 -8285
rect 95014 -8327 95083 -8293
rect 95086 -8327 95127 -8293
rect 95198 -8327 95239 -8293
rect 95729 -8317 95770 -8283
rect 95825 -8317 95866 -8283
rect 95921 -8317 95962 -8283
rect 96017 -8317 96058 -8283
rect 96113 -8317 96154 -8283
rect 97138 -8324 97179 -8290
rect 97183 -8324 97190 -8279
rect 94848 -8367 94889 -8333
rect 95441 -8336 95448 -8328
rect 95541 -8336 95548 -8328
rect 94837 -8417 94844 -8406
rect 94848 -8417 94853 -8367
rect 95042 -8410 95083 -8376
rect 95087 -8410 95094 -8365
rect 95187 -8376 95194 -8365
rect 95368 -8370 95437 -8336
rect 95440 -8370 95481 -8336
rect 95552 -8370 95593 -8336
rect 96277 -8360 96318 -8326
rect 96373 -8360 96414 -8326
rect 96469 -8360 96510 -8326
rect 96565 -8360 96606 -8326
rect 96661 -8360 96702 -8326
rect 96757 -8360 96798 -8326
rect 96853 -8360 96894 -8326
rect 95198 -8410 95239 -8376
rect 95831 -8379 95838 -8371
rect 94848 -8451 94889 -8417
rect 94837 -8500 94844 -8489
rect 94848 -8500 94853 -8451
rect 95042 -8494 95083 -8460
rect 95087 -8494 95094 -8449
rect 95187 -8460 95194 -8449
rect 95396 -8453 95437 -8419
rect 95441 -8453 95448 -8408
rect 95541 -8419 95548 -8408
rect 95722 -8413 95763 -8379
rect 95786 -8413 95838 -8379
rect 95866 -8413 95907 -8379
rect 95552 -8453 95593 -8419
rect 95198 -8494 95239 -8460
rect 94848 -8534 94889 -8500
rect 94848 -8568 94853 -8534
rect 93498 -8740 93503 -8706
rect 93794 -8723 93835 -8689
rect 93839 -8723 93846 -8681
rect 93981 -8741 93993 -8673
rect 94022 -8707 94027 -8639
rect 94067 -8671 94072 -8603
rect 94101 -8637 94106 -8571
rect 95042 -8577 95083 -8543
rect 95087 -8577 95094 -8532
rect 95187 -8543 95194 -8532
rect 95396 -8537 95437 -8503
rect 95441 -8537 95448 -8492
rect 95541 -8503 95548 -8492
rect 95786 -8496 95827 -8462
rect 95831 -8496 95838 -8451
rect 95552 -8537 95593 -8503
rect 95198 -8577 95239 -8543
rect 94111 -8621 94152 -8587
rect 94312 -8666 94353 -8632
rect 94081 -8689 94088 -8681
rect 94092 -8723 94133 -8689
rect 94312 -8734 94353 -8700
rect 91245 -8906 91286 -8872
rect 91317 -8906 91358 -8872
rect 91389 -8906 91430 -8872
rect 91702 -8913 91743 -8879
rect 91747 -8913 91754 -8868
rect 91847 -8879 91854 -8868
rect 91858 -8913 91899 -8879
rect 92442 -8895 92483 -8861
rect 92487 -8895 92494 -8853
rect 90336 -8959 90818 -8925
rect 91670 -8949 91711 -8915
rect 91742 -8949 91783 -8915
rect 92056 -8956 92097 -8922
rect 92101 -8956 92108 -8911
rect 92201 -8922 92208 -8911
rect 92629 -8913 92641 -8845
rect 92670 -8879 92675 -8811
rect 92715 -8843 92720 -8775
rect 92749 -8809 92754 -8743
rect 93981 -8753 93988 -8741
rect 94361 -8750 94366 -8616
rect 92759 -8793 92800 -8759
rect 92962 -8838 93003 -8804
rect 92729 -8861 92736 -8853
rect 92740 -8895 92781 -8861
rect 92962 -8906 93003 -8872
rect 92212 -8956 92253 -8922
rect 90336 -8985 90805 -8959
rect 90340 -8993 90547 -8985
rect 90356 -9003 90531 -8993
rect 90082 -9140 90263 -9114
rect 89589 -9174 89630 -9140
rect 89685 -9174 89726 -9140
rect 89781 -9174 89822 -9140
rect 89877 -9174 89918 -9140
rect 89973 -9174 90014 -9140
rect 90069 -9174 90263 -9140
rect 90082 -9200 90263 -9174
rect 90282 -9174 90389 -9050
rect 90541 -9062 90547 -9051
rect 90160 -9870 90201 -9200
rect 90282 -9228 90291 -9174
rect 89967 -9936 90118 -9924
rect 89635 -9970 90118 -9936
rect 89967 -9971 90118 -9970
rect 90148 -9971 90201 -9870
rect 90294 -9971 90335 -9174
rect 90340 -9971 90346 -9174
rect 90552 -9971 90593 -9062
rect 90686 -9971 90727 -8985
rect 90939 -9002 90980 -8968
rect 91035 -9002 91076 -8968
rect 91131 -9002 91172 -8968
rect 91227 -9002 91268 -8968
rect 91323 -9002 91364 -8968
rect 91419 -9002 91460 -8968
rect 91515 -9002 91556 -8968
rect 92024 -8992 92065 -8958
rect 92096 -8992 92137 -8958
rect 92442 -8995 92483 -8961
rect 92487 -8995 92494 -8950
rect 92629 -9001 92636 -8913
rect 93011 -8922 93016 -8788
rect 92729 -8961 92736 -8950
rect 93045 -8956 93050 -8762
rect 93085 -8778 93092 -8767
rect 93081 -8809 93092 -8778
rect 93407 -8796 93448 -8762
rect 92740 -8995 92781 -8961
rect 91677 -9045 91718 -9011
rect 91773 -9045 91814 -9011
rect 91869 -9045 91910 -9011
rect 92378 -9035 92419 -9001
rect 92450 -9035 92491 -9001
rect 92522 -9035 92563 -9001
rect 92594 -9029 92636 -9001
rect 92940 -9025 92981 -8991
rect 92985 -9025 92992 -8980
rect 93081 -8992 93086 -8809
rect 93115 -8995 93120 -8812
rect 92594 -9035 92635 -9029
rect 92031 -9088 92072 -9054
rect 92127 -9088 92168 -9054
rect 92223 -9088 92264 -9054
rect 93127 -9076 93134 -8809
rect 93756 -8819 94149 -8753
rect 94395 -8784 94400 -8590
rect 94435 -8606 94442 -8595
rect 94431 -8637 94442 -8606
rect 94757 -8624 94798 -8590
rect 93143 -8860 93184 -8826
rect 93492 -8830 93509 -8819
rect 93492 -8832 93498 -8830
rect 93143 -8928 93184 -8894
rect 93195 -8995 93200 -8860
rect 93426 -8874 93498 -8832
rect 93554 -8874 94149 -8819
rect 94290 -8853 94331 -8819
rect 94335 -8853 94342 -8808
rect 94431 -8820 94436 -8637
rect 94465 -8823 94470 -8640
rect 93426 -8877 94149 -8874
rect 93229 -8980 93234 -8892
rect 93346 -8942 93387 -8908
rect 93391 -8942 93398 -8900
rect 93227 -8991 93234 -8980
rect 93229 -9025 93234 -8991
rect 93238 -9025 93279 -8991
rect 93346 -9042 93387 -9008
rect 93391 -9042 93398 -8997
rect 93239 -9078 93280 -9044
rect 93311 -9078 93352 -9044
rect 93383 -9078 93424 -9044
rect 92385 -9131 92426 -9097
rect 92481 -9131 92522 -9097
rect 92577 -9131 92618 -9097
rect 92673 -9131 92714 -9097
rect 92769 -9131 92810 -9097
rect 93426 -9114 93577 -8877
rect 93756 -8899 94149 -8877
rect 93680 -8925 94149 -8899
rect 94477 -8904 94484 -8637
rect 94493 -8688 94534 -8654
rect 94493 -8756 94534 -8722
rect 94545 -8823 94550 -8688
rect 95107 -8691 95148 -8657
rect 95159 -8718 95164 -8641
rect 94579 -8808 94584 -8720
rect 94696 -8770 94737 -8736
rect 94741 -8770 94748 -8728
rect 94841 -8740 94848 -8729
rect 94852 -8774 94893 -8740
rect 95193 -8752 95198 -8607
rect 95396 -8620 95437 -8586
rect 95441 -8620 95448 -8575
rect 95541 -8586 95548 -8575
rect 95786 -8580 95827 -8546
rect 95831 -8580 95838 -8535
rect 95552 -8620 95593 -8586
rect 95461 -8734 95502 -8700
rect 95513 -8761 95518 -8684
rect 94577 -8819 94584 -8808
rect 95046 -8813 95087 -8779
rect 95091 -8813 95098 -8771
rect 95191 -8779 95198 -8771
rect 95202 -8813 95243 -8779
rect 95547 -8795 95552 -8650
rect 95786 -8663 95827 -8629
rect 95831 -8663 95838 -8618
rect 95908 -8679 95913 -8363
rect 95931 -8379 95938 -8371
rect 95942 -8379 95947 -8363
rect 95942 -8413 95983 -8379
rect 95987 -8413 95994 -8371
rect 95931 -8462 95938 -8451
rect 95942 -8462 95947 -8413
rect 95942 -8496 95983 -8462
rect 95987 -8496 95994 -8451
rect 95931 -8546 95938 -8535
rect 95942 -8546 95947 -8496
rect 95942 -8580 95983 -8546
rect 95987 -8580 95994 -8535
rect 95931 -8629 95938 -8618
rect 95942 -8629 95947 -8580
rect 95942 -8663 95983 -8629
rect 95987 -8663 95994 -8618
rect 95931 -8697 95938 -8671
rect 95942 -8713 95947 -8663
rect 95851 -8777 95892 -8743
rect 94579 -8853 94584 -8819
rect 94588 -8853 94629 -8819
rect 94696 -8870 94737 -8836
rect 94741 -8870 94748 -8825
rect 94841 -8832 94848 -8821
rect 94852 -8866 94893 -8832
rect 95400 -8856 95441 -8822
rect 95445 -8856 95452 -8814
rect 95545 -8822 95552 -8814
rect 95556 -8856 95597 -8822
rect 95973 -8845 95980 -8697
rect 95996 -8713 95999 -8363
rect 96030 -8679 96033 -8363
rect 96087 -8379 96094 -8371
rect 96036 -8413 96077 -8379
rect 96098 -8413 96149 -8379
rect 96808 -8422 96813 -8406
rect 96831 -8422 96838 -8414
rect 96842 -8422 96847 -8406
rect 97138 -8408 97179 -8374
rect 97183 -8408 97190 -8363
rect 96087 -8462 96094 -8451
rect 96268 -8456 96309 -8422
rect 96340 -8456 96381 -8422
rect 96412 -8456 96453 -8422
rect 96556 -8456 96597 -8422
rect 96628 -8456 96741 -8422
rect 96772 -8456 96813 -8422
rect 96098 -8496 96139 -8462
rect 96087 -8546 96094 -8535
rect 96665 -8539 96706 -8505
rect 96098 -8580 96139 -8546
rect 96087 -8629 96094 -8618
rect 96098 -8663 96139 -8629
rect 96330 -8689 96371 -8655
rect 96375 -8689 96382 -8644
rect 96452 -8706 96457 -8588
rect 96475 -8655 96482 -8644
rect 96486 -8655 96491 -8622
rect 96522 -8655 96527 -8622
rect 96486 -8689 96527 -8655
rect 96531 -8689 96538 -8644
rect 96486 -8740 96491 -8689
rect 96522 -8740 96527 -8689
rect 96556 -8706 96561 -8589
rect 96665 -8623 96706 -8589
rect 96665 -8706 96706 -8672
rect 96808 -8706 96813 -8456
rect 96842 -8456 96883 -8422
rect 96831 -8505 96838 -8494
rect 96842 -8505 96847 -8456
rect 97138 -8491 97179 -8457
rect 97183 -8491 97190 -8446
rect 96842 -8539 96883 -8505
rect 96831 -8589 96838 -8578
rect 96842 -8589 96847 -8539
rect 96991 -8565 97100 -8499
rect 97260 -8507 97265 -8191
rect 97283 -8207 97290 -8199
rect 97294 -8207 97299 -8191
rect 97294 -8241 97335 -8207
rect 97339 -8241 97346 -8199
rect 97283 -8290 97290 -8279
rect 97294 -8290 97299 -8241
rect 97294 -8324 97335 -8290
rect 97339 -8324 97346 -8279
rect 97283 -8374 97290 -8363
rect 97294 -8374 97299 -8324
rect 97294 -8408 97335 -8374
rect 97339 -8408 97346 -8363
rect 97283 -8457 97290 -8446
rect 97294 -8457 97299 -8408
rect 97294 -8491 97335 -8457
rect 97339 -8491 97346 -8446
rect 97283 -8525 97290 -8499
rect 97294 -8541 97299 -8491
rect 96842 -8623 96883 -8589
rect 97203 -8605 97244 -8571
rect 96831 -8672 96838 -8661
rect 96842 -8672 96847 -8623
rect 96842 -8706 96883 -8672
rect 97325 -8673 97332 -8525
rect 97348 -8541 97351 -8191
rect 97382 -8507 97385 -8191
rect 97439 -8207 97446 -8199
rect 97388 -8241 97429 -8207
rect 97450 -8241 97501 -8207
rect 98365 -8231 98406 -8197
rect 98461 -8231 98502 -8197
rect 98557 -8231 98598 -8197
rect 100527 -8207 100534 -8199
rect 98158 -8250 98163 -8234
rect 98181 -8250 98188 -8242
rect 98192 -8250 98197 -8234
rect 97439 -8290 97446 -8279
rect 97618 -8284 97659 -8250
rect 97690 -8284 97731 -8250
rect 97762 -8284 97803 -8250
rect 97906 -8284 97947 -8250
rect 97978 -8284 98091 -8250
rect 98122 -8284 98163 -8250
rect 97450 -8324 97491 -8290
rect 97439 -8374 97446 -8363
rect 98015 -8367 98056 -8333
rect 97450 -8408 97491 -8374
rect 97439 -8457 97446 -8446
rect 97450 -8491 97491 -8457
rect 97680 -8517 97721 -8483
rect 97725 -8517 97732 -8472
rect 97802 -8534 97807 -8416
rect 97825 -8483 97832 -8472
rect 97836 -8483 97841 -8450
rect 97872 -8483 97877 -8450
rect 97836 -8517 97877 -8483
rect 97881 -8517 97888 -8472
rect 97836 -8568 97841 -8517
rect 97872 -8568 97877 -8517
rect 97906 -8534 97911 -8417
rect 98015 -8451 98056 -8417
rect 98015 -8534 98056 -8500
rect 98158 -8534 98163 -8284
rect 98192 -8284 98233 -8250
rect 98719 -8274 98760 -8240
rect 98815 -8274 98856 -8240
rect 98911 -8274 98952 -8240
rect 100418 -8241 100459 -8207
rect 100482 -8241 100534 -8207
rect 100562 -8241 100603 -8207
rect 98181 -8333 98188 -8322
rect 98192 -8333 98197 -8284
rect 98431 -8293 98438 -8285
rect 98531 -8293 98538 -8285
rect 98358 -8327 98427 -8293
rect 98430 -8327 98471 -8293
rect 98542 -8327 98583 -8293
rect 99073 -8317 99114 -8283
rect 99169 -8317 99210 -8283
rect 99265 -8317 99306 -8283
rect 99361 -8317 99402 -8283
rect 99457 -8317 99498 -8283
rect 100482 -8324 100523 -8290
rect 100527 -8324 100534 -8279
rect 98192 -8367 98233 -8333
rect 98785 -8336 98792 -8328
rect 98885 -8336 98892 -8328
rect 98181 -8417 98188 -8406
rect 98192 -8417 98197 -8367
rect 98386 -8410 98427 -8376
rect 98431 -8410 98438 -8365
rect 98531 -8376 98538 -8365
rect 98712 -8370 98781 -8336
rect 98784 -8370 98825 -8336
rect 98896 -8370 98937 -8336
rect 99621 -8360 99662 -8326
rect 99717 -8360 99758 -8326
rect 99813 -8360 99854 -8326
rect 99909 -8360 99950 -8326
rect 100005 -8360 100046 -8326
rect 100101 -8360 100142 -8326
rect 100197 -8360 100238 -8326
rect 98542 -8410 98583 -8376
rect 99175 -8379 99182 -8371
rect 98192 -8451 98233 -8417
rect 98181 -8500 98188 -8489
rect 98192 -8500 98197 -8451
rect 98386 -8494 98427 -8460
rect 98431 -8494 98438 -8449
rect 98531 -8460 98538 -8449
rect 98740 -8453 98781 -8419
rect 98785 -8453 98792 -8408
rect 98885 -8419 98892 -8408
rect 99066 -8413 99107 -8379
rect 99130 -8413 99182 -8379
rect 99210 -8413 99251 -8379
rect 98896 -8453 98937 -8419
rect 98542 -8494 98583 -8460
rect 98192 -8534 98233 -8500
rect 98192 -8568 98197 -8534
rect 96842 -8740 96847 -8706
rect 97138 -8723 97179 -8689
rect 97183 -8723 97190 -8681
rect 97325 -8741 97337 -8673
rect 97366 -8707 97371 -8639
rect 97411 -8671 97416 -8603
rect 97445 -8637 97450 -8571
rect 98386 -8577 98427 -8543
rect 98431 -8577 98438 -8532
rect 98531 -8543 98538 -8532
rect 98740 -8537 98781 -8503
rect 98785 -8537 98792 -8492
rect 98885 -8503 98892 -8492
rect 99130 -8496 99171 -8462
rect 99175 -8496 99182 -8451
rect 98896 -8537 98937 -8503
rect 98542 -8577 98583 -8543
rect 97455 -8621 97496 -8587
rect 97656 -8666 97697 -8632
rect 97425 -8689 97432 -8681
rect 97436 -8723 97477 -8689
rect 97656 -8734 97697 -8700
rect 94589 -8906 94630 -8872
rect 94661 -8906 94702 -8872
rect 94733 -8906 94774 -8872
rect 95046 -8913 95087 -8879
rect 95091 -8913 95098 -8868
rect 95191 -8879 95198 -8868
rect 95202 -8913 95243 -8879
rect 95786 -8895 95827 -8861
rect 95831 -8895 95838 -8853
rect 93680 -8959 94162 -8925
rect 95014 -8949 95055 -8915
rect 95086 -8949 95127 -8915
rect 95400 -8956 95441 -8922
rect 95445 -8956 95452 -8911
rect 95545 -8922 95552 -8911
rect 95973 -8913 95985 -8845
rect 96014 -8879 96019 -8811
rect 96059 -8843 96064 -8775
rect 96093 -8809 96098 -8743
rect 97325 -8753 97332 -8741
rect 97705 -8750 97710 -8616
rect 96103 -8793 96144 -8759
rect 96306 -8838 96347 -8804
rect 96073 -8861 96080 -8853
rect 96084 -8895 96125 -8861
rect 96306 -8906 96347 -8872
rect 95556 -8956 95597 -8922
rect 93680 -8985 94149 -8959
rect 93684 -8993 93891 -8985
rect 93700 -9003 93875 -8993
rect 93426 -9140 93607 -9114
rect 92933 -9174 92974 -9140
rect 93029 -9174 93070 -9140
rect 93125 -9174 93166 -9140
rect 93221 -9174 93262 -9140
rect 93317 -9174 93358 -9140
rect 93413 -9174 93607 -9140
rect 93426 -9200 93607 -9174
rect 93626 -9174 93733 -9050
rect 93885 -9062 93891 -9051
rect 93504 -9870 93545 -9200
rect 93626 -9228 93635 -9174
rect 93311 -9936 93462 -9924
rect 92979 -9970 93462 -9936
rect 93311 -9971 93462 -9970
rect 93492 -9971 93545 -9870
rect 93638 -9971 93679 -9174
rect 93684 -9971 93690 -9174
rect 93896 -9971 93937 -9062
rect 94030 -9971 94071 -8985
rect 94283 -9002 94324 -8968
rect 94379 -9002 94420 -8968
rect 94475 -9002 94516 -8968
rect 94571 -9002 94612 -8968
rect 94667 -9002 94708 -8968
rect 94763 -9002 94804 -8968
rect 94859 -9002 94900 -8968
rect 95368 -8992 95409 -8958
rect 95440 -8992 95481 -8958
rect 95786 -8995 95827 -8961
rect 95831 -8995 95838 -8950
rect 95973 -9001 95980 -8913
rect 96355 -8922 96360 -8788
rect 96073 -8961 96080 -8950
rect 96389 -8956 96394 -8762
rect 96429 -8778 96436 -8767
rect 96425 -8809 96436 -8778
rect 96751 -8796 96792 -8762
rect 96084 -8995 96125 -8961
rect 95021 -9045 95062 -9011
rect 95117 -9045 95158 -9011
rect 95213 -9045 95254 -9011
rect 95722 -9035 95763 -9001
rect 95794 -9035 95835 -9001
rect 95866 -9035 95907 -9001
rect 95938 -9029 95980 -9001
rect 96284 -9025 96325 -8991
rect 96329 -9025 96336 -8980
rect 96425 -8992 96430 -8809
rect 96459 -8995 96464 -8812
rect 95938 -9035 95979 -9029
rect 95375 -9088 95416 -9054
rect 95471 -9088 95512 -9054
rect 95567 -9088 95608 -9054
rect 96471 -9076 96478 -8809
rect 97100 -8819 97493 -8753
rect 97739 -8784 97744 -8590
rect 97779 -8606 97786 -8595
rect 97775 -8637 97786 -8606
rect 98101 -8624 98142 -8590
rect 96487 -8860 96528 -8826
rect 96836 -8830 96853 -8819
rect 96836 -8832 96842 -8830
rect 96487 -8928 96528 -8894
rect 96539 -8995 96544 -8860
rect 96770 -8874 96842 -8832
rect 96898 -8874 97493 -8819
rect 97634 -8853 97675 -8819
rect 97679 -8853 97686 -8808
rect 97775 -8820 97780 -8637
rect 97809 -8823 97814 -8640
rect 96770 -8877 97493 -8874
rect 96573 -8980 96578 -8892
rect 96690 -8942 96731 -8908
rect 96735 -8942 96742 -8900
rect 96571 -8991 96578 -8980
rect 96573 -9025 96578 -8991
rect 96582 -9025 96623 -8991
rect 96690 -9042 96731 -9008
rect 96735 -9042 96742 -8997
rect 96583 -9078 96624 -9044
rect 96655 -9078 96696 -9044
rect 96727 -9078 96768 -9044
rect 95729 -9131 95770 -9097
rect 95825 -9131 95866 -9097
rect 95921 -9131 95962 -9097
rect 96017 -9131 96058 -9097
rect 96113 -9131 96154 -9097
rect 96770 -9114 96921 -8877
rect 97100 -8899 97493 -8877
rect 97024 -8925 97493 -8899
rect 97821 -8904 97828 -8637
rect 97837 -8688 97878 -8654
rect 97837 -8756 97878 -8722
rect 97889 -8823 97894 -8688
rect 98451 -8691 98492 -8657
rect 98503 -8718 98508 -8641
rect 97923 -8808 97928 -8720
rect 98040 -8770 98081 -8736
rect 98085 -8770 98092 -8728
rect 98185 -8740 98192 -8729
rect 98196 -8774 98237 -8740
rect 98537 -8752 98542 -8607
rect 98740 -8620 98781 -8586
rect 98785 -8620 98792 -8575
rect 98885 -8586 98892 -8575
rect 99130 -8580 99171 -8546
rect 99175 -8580 99182 -8535
rect 98896 -8620 98937 -8586
rect 98805 -8734 98846 -8700
rect 98857 -8761 98862 -8684
rect 97921 -8819 97928 -8808
rect 98390 -8813 98431 -8779
rect 98435 -8813 98442 -8771
rect 98535 -8779 98542 -8771
rect 98546 -8813 98587 -8779
rect 98891 -8795 98896 -8650
rect 99130 -8663 99171 -8629
rect 99175 -8663 99182 -8618
rect 99252 -8679 99257 -8363
rect 99275 -8379 99282 -8371
rect 99286 -8379 99291 -8363
rect 99286 -8413 99327 -8379
rect 99331 -8413 99338 -8371
rect 99275 -8462 99282 -8451
rect 99286 -8462 99291 -8413
rect 99286 -8496 99327 -8462
rect 99331 -8496 99338 -8451
rect 99275 -8546 99282 -8535
rect 99286 -8546 99291 -8496
rect 99286 -8580 99327 -8546
rect 99331 -8580 99338 -8535
rect 99275 -8629 99282 -8618
rect 99286 -8629 99291 -8580
rect 99286 -8663 99327 -8629
rect 99331 -8663 99338 -8618
rect 99275 -8697 99282 -8671
rect 99286 -8713 99291 -8663
rect 99195 -8777 99236 -8743
rect 97923 -8853 97928 -8819
rect 97932 -8853 97973 -8819
rect 98040 -8870 98081 -8836
rect 98085 -8870 98092 -8825
rect 98185 -8832 98192 -8821
rect 98196 -8866 98237 -8832
rect 98744 -8856 98785 -8822
rect 98789 -8856 98796 -8814
rect 98889 -8822 98896 -8814
rect 98900 -8856 98941 -8822
rect 99317 -8845 99324 -8697
rect 99340 -8713 99343 -8363
rect 99374 -8679 99377 -8363
rect 99431 -8379 99438 -8371
rect 99380 -8413 99421 -8379
rect 99442 -8413 99493 -8379
rect 100152 -8422 100157 -8406
rect 100175 -8422 100182 -8414
rect 100186 -8422 100191 -8406
rect 100482 -8408 100523 -8374
rect 100527 -8408 100534 -8363
rect 99431 -8462 99438 -8451
rect 99612 -8456 99653 -8422
rect 99684 -8456 99725 -8422
rect 99756 -8456 99797 -8422
rect 99900 -8456 99941 -8422
rect 99972 -8456 100085 -8422
rect 100116 -8456 100157 -8422
rect 99442 -8496 99483 -8462
rect 99431 -8546 99438 -8535
rect 100009 -8539 100050 -8505
rect 99442 -8580 99483 -8546
rect 99431 -8629 99438 -8618
rect 99442 -8663 99483 -8629
rect 99674 -8689 99715 -8655
rect 99719 -8689 99726 -8644
rect 99796 -8706 99801 -8588
rect 99819 -8655 99826 -8644
rect 99830 -8655 99835 -8622
rect 99866 -8655 99871 -8622
rect 99830 -8689 99871 -8655
rect 99875 -8689 99882 -8644
rect 99830 -8740 99835 -8689
rect 99866 -8740 99871 -8689
rect 99900 -8706 99905 -8589
rect 100009 -8623 100050 -8589
rect 100009 -8706 100050 -8672
rect 100152 -8706 100157 -8456
rect 100186 -8456 100227 -8422
rect 100175 -8505 100182 -8494
rect 100186 -8505 100191 -8456
rect 100482 -8491 100523 -8457
rect 100527 -8491 100534 -8446
rect 100186 -8539 100227 -8505
rect 100175 -8589 100182 -8578
rect 100186 -8589 100191 -8539
rect 100335 -8565 100444 -8499
rect 100604 -8507 100609 -8191
rect 100627 -8207 100634 -8199
rect 100638 -8207 100643 -8191
rect 100638 -8241 100679 -8207
rect 100683 -8241 100690 -8199
rect 100627 -8290 100634 -8279
rect 100638 -8290 100643 -8241
rect 100638 -8324 100679 -8290
rect 100683 -8324 100690 -8279
rect 100627 -8374 100634 -8363
rect 100638 -8374 100643 -8324
rect 100638 -8408 100679 -8374
rect 100683 -8408 100690 -8363
rect 100627 -8457 100634 -8446
rect 100638 -8457 100643 -8408
rect 100638 -8491 100679 -8457
rect 100683 -8491 100690 -8446
rect 100627 -8525 100634 -8499
rect 100638 -8541 100643 -8491
rect 100186 -8623 100227 -8589
rect 100547 -8605 100588 -8571
rect 100175 -8672 100182 -8661
rect 100186 -8672 100191 -8623
rect 100186 -8706 100227 -8672
rect 100669 -8673 100676 -8525
rect 100692 -8541 100695 -8191
rect 100726 -8507 100729 -8191
rect 100783 -8207 100790 -8199
rect 100732 -8241 100773 -8207
rect 100794 -8241 100845 -8207
rect 101709 -8231 101750 -8197
rect 101805 -8231 101846 -8197
rect 101901 -8231 101942 -8197
rect 103871 -8207 103878 -8199
rect 101502 -8250 101507 -8234
rect 101525 -8250 101532 -8242
rect 101536 -8250 101541 -8234
rect 100783 -8290 100790 -8279
rect 100962 -8284 101003 -8250
rect 101034 -8284 101075 -8250
rect 101106 -8284 101147 -8250
rect 101250 -8284 101291 -8250
rect 101322 -8284 101435 -8250
rect 101466 -8284 101507 -8250
rect 100794 -8324 100835 -8290
rect 100783 -8374 100790 -8363
rect 101359 -8367 101400 -8333
rect 100794 -8408 100835 -8374
rect 100783 -8457 100790 -8446
rect 100794 -8491 100835 -8457
rect 101024 -8517 101065 -8483
rect 101069 -8517 101076 -8472
rect 101146 -8534 101151 -8416
rect 101169 -8483 101176 -8472
rect 101180 -8483 101185 -8450
rect 101216 -8483 101221 -8450
rect 101180 -8517 101221 -8483
rect 101225 -8517 101232 -8472
rect 101180 -8568 101185 -8517
rect 101216 -8568 101221 -8517
rect 101250 -8534 101255 -8417
rect 101359 -8451 101400 -8417
rect 101359 -8534 101400 -8500
rect 101502 -8534 101507 -8284
rect 101536 -8284 101577 -8250
rect 102063 -8274 102104 -8240
rect 102159 -8274 102200 -8240
rect 102255 -8274 102296 -8240
rect 103762 -8241 103803 -8207
rect 103826 -8241 103878 -8207
rect 103906 -8241 103947 -8207
rect 101525 -8333 101532 -8322
rect 101536 -8333 101541 -8284
rect 101775 -8293 101782 -8285
rect 101875 -8293 101882 -8285
rect 101702 -8327 101771 -8293
rect 101774 -8327 101815 -8293
rect 101886 -8327 101927 -8293
rect 102417 -8317 102458 -8283
rect 102513 -8317 102554 -8283
rect 102609 -8317 102650 -8283
rect 102705 -8317 102746 -8283
rect 102801 -8317 102842 -8283
rect 103826 -8324 103867 -8290
rect 103871 -8324 103878 -8279
rect 101536 -8367 101577 -8333
rect 102129 -8336 102136 -8328
rect 102229 -8336 102236 -8328
rect 101525 -8417 101532 -8406
rect 101536 -8417 101541 -8367
rect 101730 -8410 101771 -8376
rect 101775 -8410 101782 -8365
rect 101875 -8376 101882 -8365
rect 102056 -8370 102125 -8336
rect 102128 -8370 102169 -8336
rect 102240 -8370 102281 -8336
rect 102965 -8360 103006 -8326
rect 103061 -8360 103102 -8326
rect 103157 -8360 103198 -8326
rect 103253 -8360 103294 -8326
rect 103349 -8360 103390 -8326
rect 103445 -8360 103486 -8326
rect 103541 -8360 103582 -8326
rect 101886 -8410 101927 -8376
rect 102519 -8379 102526 -8371
rect 101536 -8451 101577 -8417
rect 101525 -8500 101532 -8489
rect 101536 -8500 101541 -8451
rect 101730 -8494 101771 -8460
rect 101775 -8494 101782 -8449
rect 101875 -8460 101882 -8449
rect 102084 -8453 102125 -8419
rect 102129 -8453 102136 -8408
rect 102229 -8419 102236 -8408
rect 102410 -8413 102451 -8379
rect 102474 -8413 102526 -8379
rect 102554 -8413 102595 -8379
rect 102240 -8453 102281 -8419
rect 101886 -8494 101927 -8460
rect 101536 -8534 101577 -8500
rect 101536 -8568 101541 -8534
rect 100186 -8740 100191 -8706
rect 100482 -8723 100523 -8689
rect 100527 -8723 100534 -8681
rect 100669 -8741 100681 -8673
rect 100710 -8707 100715 -8639
rect 100755 -8671 100760 -8603
rect 100789 -8637 100794 -8571
rect 101730 -8577 101771 -8543
rect 101775 -8577 101782 -8532
rect 101875 -8543 101882 -8532
rect 102084 -8537 102125 -8503
rect 102129 -8537 102136 -8492
rect 102229 -8503 102236 -8492
rect 102474 -8496 102515 -8462
rect 102519 -8496 102526 -8451
rect 102240 -8537 102281 -8503
rect 101886 -8577 101927 -8543
rect 100800 -8621 100840 -8587
rect 101000 -8666 101041 -8632
rect 100769 -8689 100776 -8681
rect 100780 -8723 100821 -8689
rect 101000 -8734 101041 -8700
rect 97933 -8906 97974 -8872
rect 98005 -8906 98046 -8872
rect 98077 -8906 98118 -8872
rect 98390 -8913 98431 -8879
rect 98435 -8913 98442 -8868
rect 98535 -8879 98542 -8868
rect 98546 -8913 98587 -8879
rect 99130 -8895 99171 -8861
rect 99175 -8895 99182 -8853
rect 97024 -8959 97506 -8925
rect 98358 -8949 98399 -8915
rect 98430 -8949 98471 -8915
rect 98744 -8956 98785 -8922
rect 98789 -8956 98796 -8911
rect 98889 -8922 98896 -8911
rect 99317 -8913 99329 -8845
rect 99358 -8879 99363 -8811
rect 99403 -8843 99408 -8775
rect 99437 -8809 99442 -8743
rect 100669 -8753 100676 -8741
rect 101049 -8750 101054 -8616
rect 99447 -8793 99488 -8759
rect 99650 -8838 99691 -8804
rect 99417 -8861 99424 -8853
rect 99428 -8895 99469 -8861
rect 99650 -8906 99691 -8872
rect 98900 -8956 98941 -8922
rect 97024 -8985 97493 -8959
rect 97028 -8993 97235 -8985
rect 97044 -9003 97219 -8993
rect 96770 -9140 96951 -9114
rect 96277 -9174 96318 -9140
rect 96373 -9174 96414 -9140
rect 96469 -9174 96510 -9140
rect 96565 -9174 96606 -9140
rect 96661 -9174 96702 -9140
rect 96757 -9174 96951 -9140
rect 96770 -9200 96951 -9174
rect 96970 -9174 97077 -9050
rect 97229 -9062 97235 -9051
rect 96848 -9870 96889 -9200
rect 96970 -9228 96979 -9174
rect 96655 -9936 96806 -9924
rect 96323 -9970 96806 -9936
rect 96655 -9971 96806 -9970
rect 96836 -9971 96889 -9870
rect 96982 -9971 97023 -9174
rect 97028 -9971 97034 -9174
rect 97240 -9971 97281 -9062
rect 97374 -9971 97415 -8985
rect 97627 -9002 97668 -8968
rect 97723 -9002 97764 -8968
rect 97819 -9002 97860 -8968
rect 97915 -9002 97956 -8968
rect 98011 -9002 98052 -8968
rect 98107 -9002 98148 -8968
rect 98203 -9002 98244 -8968
rect 98712 -8992 98753 -8958
rect 98784 -8992 98825 -8958
rect 99130 -8995 99171 -8961
rect 99175 -8995 99182 -8950
rect 99317 -9001 99324 -8913
rect 99699 -8922 99704 -8788
rect 99417 -8961 99424 -8950
rect 99733 -8956 99738 -8762
rect 99773 -8778 99780 -8767
rect 99769 -8809 99780 -8778
rect 100095 -8796 100136 -8762
rect 99428 -8995 99469 -8961
rect 98365 -9045 98406 -9011
rect 98461 -9045 98502 -9011
rect 98557 -9045 98598 -9011
rect 99066 -9035 99107 -9001
rect 99138 -9035 99179 -9001
rect 99210 -9035 99251 -9001
rect 99282 -9029 99324 -9001
rect 99628 -9025 99669 -8991
rect 99673 -9025 99680 -8980
rect 99769 -8992 99774 -8809
rect 99803 -8995 99808 -8812
rect 99282 -9035 99323 -9029
rect 98719 -9088 98760 -9054
rect 98815 -9088 98856 -9054
rect 98911 -9088 98952 -9054
rect 99815 -9076 99822 -8809
rect 100444 -8819 100837 -8753
rect 101083 -8784 101088 -8590
rect 101123 -8606 101130 -8595
rect 101119 -8637 101130 -8606
rect 101445 -8624 101486 -8590
rect 99831 -8860 99872 -8826
rect 100180 -8830 100197 -8819
rect 100180 -8832 100186 -8830
rect 99831 -8928 99872 -8894
rect 99883 -8995 99888 -8860
rect 100114 -8874 100186 -8832
rect 100242 -8874 100837 -8819
rect 100978 -8853 101019 -8819
rect 101023 -8853 101030 -8808
rect 101119 -8820 101124 -8637
rect 101153 -8823 101158 -8640
rect 100114 -8877 100837 -8874
rect 99917 -8980 99922 -8892
rect 100034 -8942 100075 -8908
rect 100079 -8942 100086 -8900
rect 99915 -8991 99922 -8980
rect 99917 -9025 99922 -8991
rect 99926 -9025 99967 -8991
rect 100034 -9042 100075 -9008
rect 100079 -9042 100086 -8997
rect 99927 -9078 99968 -9044
rect 99999 -9078 100040 -9044
rect 100071 -9078 100112 -9044
rect 99073 -9131 99114 -9097
rect 99169 -9131 99210 -9097
rect 99265 -9131 99306 -9097
rect 99361 -9131 99402 -9097
rect 99457 -9131 99498 -9097
rect 100114 -9114 100265 -8877
rect 100444 -8899 100837 -8877
rect 100368 -8925 100837 -8899
rect 101165 -8904 101172 -8637
rect 101181 -8688 101222 -8654
rect 101181 -8756 101222 -8722
rect 101233 -8823 101238 -8688
rect 101795 -8691 101836 -8657
rect 101847 -8718 101852 -8641
rect 101267 -8808 101272 -8720
rect 101384 -8770 101425 -8736
rect 101429 -8770 101436 -8728
rect 101529 -8740 101536 -8729
rect 101540 -8774 101581 -8740
rect 101881 -8752 101886 -8607
rect 102084 -8620 102125 -8586
rect 102129 -8620 102136 -8575
rect 102229 -8586 102236 -8575
rect 102474 -8580 102515 -8546
rect 102519 -8580 102526 -8535
rect 102240 -8620 102281 -8586
rect 102149 -8734 102190 -8700
rect 102201 -8761 102206 -8684
rect 101265 -8819 101272 -8808
rect 101734 -8813 101775 -8779
rect 101779 -8813 101786 -8771
rect 101879 -8779 101886 -8771
rect 101890 -8813 101931 -8779
rect 102235 -8795 102240 -8650
rect 102474 -8663 102515 -8629
rect 102519 -8663 102526 -8618
rect 102596 -8679 102601 -8363
rect 102619 -8379 102626 -8371
rect 102630 -8379 102635 -8363
rect 102630 -8413 102671 -8379
rect 102675 -8413 102682 -8371
rect 102619 -8462 102626 -8451
rect 102630 -8462 102635 -8413
rect 102630 -8496 102671 -8462
rect 102675 -8496 102682 -8451
rect 102619 -8546 102626 -8535
rect 102630 -8546 102635 -8496
rect 102630 -8580 102671 -8546
rect 102675 -8580 102682 -8535
rect 102619 -8629 102626 -8618
rect 102630 -8629 102635 -8580
rect 102630 -8663 102671 -8629
rect 102675 -8663 102682 -8618
rect 102619 -8697 102626 -8671
rect 102630 -8713 102635 -8663
rect 102539 -8777 102580 -8743
rect 101267 -8853 101272 -8819
rect 101276 -8853 101317 -8819
rect 101384 -8870 101425 -8836
rect 101429 -8870 101436 -8825
rect 101529 -8832 101536 -8821
rect 101540 -8866 101581 -8832
rect 102088 -8856 102129 -8822
rect 102133 -8856 102140 -8814
rect 102233 -8822 102240 -8814
rect 102244 -8856 102285 -8822
rect 102661 -8845 102668 -8697
rect 102684 -8713 102687 -8363
rect 102718 -8679 102721 -8363
rect 102775 -8379 102782 -8371
rect 102724 -8413 102765 -8379
rect 102786 -8413 102837 -8379
rect 103496 -8422 103501 -8406
rect 103519 -8422 103526 -8414
rect 103530 -8422 103535 -8406
rect 103826 -8408 103867 -8374
rect 103871 -8408 103878 -8363
rect 102775 -8462 102782 -8451
rect 102956 -8456 102997 -8422
rect 103028 -8456 103069 -8422
rect 103100 -8456 103141 -8422
rect 103244 -8456 103285 -8422
rect 103316 -8456 103429 -8422
rect 103460 -8456 103501 -8422
rect 102786 -8496 102827 -8462
rect 102775 -8546 102782 -8535
rect 103353 -8539 103394 -8505
rect 102786 -8580 102827 -8546
rect 102775 -8629 102782 -8618
rect 102786 -8663 102827 -8629
rect 103018 -8689 103059 -8655
rect 103063 -8689 103070 -8644
rect 103140 -8706 103145 -8588
rect 103163 -8655 103170 -8644
rect 103174 -8655 103179 -8622
rect 103210 -8655 103215 -8622
rect 103174 -8689 103215 -8655
rect 103219 -8689 103226 -8644
rect 103174 -8740 103179 -8689
rect 103210 -8740 103215 -8689
rect 103244 -8706 103249 -8589
rect 103353 -8623 103394 -8589
rect 103353 -8706 103394 -8672
rect 103496 -8706 103501 -8456
rect 103530 -8456 103571 -8422
rect 103519 -8505 103526 -8494
rect 103530 -8505 103535 -8456
rect 103826 -8491 103867 -8457
rect 103871 -8491 103878 -8446
rect 103530 -8539 103571 -8505
rect 103519 -8589 103526 -8578
rect 103530 -8589 103535 -8539
rect 103679 -8565 103788 -8499
rect 103948 -8507 103953 -8191
rect 103971 -8207 103978 -8199
rect 103982 -8207 103987 -8191
rect 103982 -8241 104023 -8207
rect 104027 -8241 104034 -8199
rect 103971 -8290 103978 -8279
rect 103982 -8290 103987 -8241
rect 103982 -8324 104023 -8290
rect 104027 -8324 104034 -8279
rect 103971 -8374 103978 -8363
rect 103982 -8374 103987 -8324
rect 103982 -8408 104023 -8374
rect 104027 -8408 104034 -8363
rect 103971 -8457 103978 -8446
rect 103982 -8457 103987 -8408
rect 103982 -8491 104023 -8457
rect 104027 -8491 104034 -8446
rect 103971 -8525 103978 -8499
rect 103982 -8541 103987 -8491
rect 103530 -8623 103571 -8589
rect 103891 -8605 103932 -8571
rect 103519 -8672 103526 -8661
rect 103530 -8672 103535 -8623
rect 103530 -8706 103571 -8672
rect 104013 -8673 104020 -8525
rect 104036 -8541 104039 -8191
rect 104070 -8507 104073 -8191
rect 104127 -8207 104134 -8199
rect 104076 -8241 104117 -8207
rect 104138 -8241 104189 -8207
rect 105053 -8231 105094 -8197
rect 105149 -8231 105190 -8197
rect 105245 -8231 105286 -8197
rect 104846 -8250 104851 -8234
rect 104869 -8250 104876 -8242
rect 104880 -8250 104885 -8234
rect 104127 -8290 104134 -8279
rect 104306 -8284 104347 -8250
rect 104378 -8284 104419 -8250
rect 104450 -8284 104491 -8250
rect 104594 -8284 104635 -8250
rect 104666 -8284 104779 -8250
rect 104810 -8284 104851 -8250
rect 104138 -8324 104179 -8290
rect 104127 -8374 104134 -8363
rect 104703 -8367 104744 -8333
rect 104138 -8408 104179 -8374
rect 104127 -8457 104134 -8446
rect 104138 -8491 104179 -8457
rect 104368 -8517 104409 -8483
rect 104413 -8517 104420 -8472
rect 104490 -8534 104495 -8416
rect 104513 -8483 104520 -8472
rect 104524 -8483 104529 -8450
rect 104560 -8483 104565 -8450
rect 104524 -8517 104565 -8483
rect 104569 -8517 104576 -8472
rect 104524 -8568 104529 -8517
rect 104560 -8568 104565 -8517
rect 104594 -8534 104599 -8417
rect 104703 -8451 104744 -8417
rect 104703 -8534 104744 -8500
rect 104846 -8534 104851 -8284
rect 104880 -8284 104921 -8250
rect 105407 -8274 105448 -8240
rect 105503 -8274 105544 -8240
rect 105599 -8274 105640 -8240
rect 107112 -8241 107147 -8207
rect 107176 -8241 107219 -8207
rect 107221 -8241 107222 -8199
rect 107321 -8207 107322 -8199
rect 107256 -8241 107291 -8207
rect 107332 -8241 107367 -8207
rect 107377 -8241 107378 -8199
rect 107477 -8207 107478 -8199
rect 107426 -8241 107461 -8207
rect 107488 -8241 107533 -8207
rect 108403 -8231 108438 -8197
rect 108499 -8231 108534 -8197
rect 108595 -8231 108630 -8197
rect 108219 -8250 108220 -8242
rect 104869 -8333 104876 -8322
rect 104880 -8333 104885 -8284
rect 105119 -8293 105126 -8285
rect 105219 -8293 105226 -8285
rect 105046 -8327 105115 -8293
rect 105118 -8327 105159 -8293
rect 105230 -8327 105271 -8293
rect 105761 -8317 105802 -8283
rect 105857 -8317 105898 -8283
rect 105953 -8317 105994 -8283
rect 106049 -8317 106090 -8283
rect 106145 -8317 106186 -8283
rect 107176 -8324 107211 -8290
rect 107221 -8324 107222 -8279
rect 107321 -8290 107322 -8279
rect 107332 -8324 107367 -8290
rect 107377 -8324 107378 -8279
rect 107477 -8290 107478 -8279
rect 107656 -8284 107691 -8250
rect 107728 -8284 107763 -8250
rect 107800 -8284 107835 -8250
rect 107944 -8284 107979 -8250
rect 108016 -8284 108051 -8250
rect 108053 -8284 108123 -8250
rect 108160 -8284 108195 -8250
rect 108230 -8284 108265 -8250
rect 108757 -8274 108792 -8240
rect 108853 -8274 108888 -8240
rect 108949 -8274 108984 -8240
rect 110456 -8241 110491 -8207
rect 110520 -8241 110563 -8207
rect 110565 -8241 110566 -8199
rect 110665 -8207 110666 -8199
rect 110600 -8241 110635 -8207
rect 110676 -8241 110711 -8207
rect 110721 -8241 110722 -8199
rect 110821 -8207 110822 -8199
rect 110770 -8241 110805 -8207
rect 110832 -8241 110877 -8207
rect 111747 -8231 111782 -8197
rect 111843 -8231 111878 -8197
rect 111939 -8231 111974 -8197
rect 111563 -8250 111564 -8242
rect 107488 -8324 107523 -8290
rect 108469 -8293 108470 -8285
rect 108569 -8293 108570 -8285
rect 104880 -8367 104921 -8333
rect 105473 -8336 105480 -8328
rect 105573 -8336 105580 -8328
rect 104869 -8417 104876 -8406
rect 104880 -8417 104885 -8367
rect 105074 -8410 105115 -8376
rect 105119 -8410 105126 -8365
rect 105219 -8376 105226 -8365
rect 105400 -8370 105469 -8336
rect 105472 -8370 105513 -8336
rect 105584 -8370 105625 -8336
rect 106309 -8360 106350 -8326
rect 106405 -8360 106446 -8326
rect 106501 -8360 106542 -8326
rect 106597 -8360 106638 -8326
rect 106693 -8360 106734 -8326
rect 106789 -8360 106830 -8326
rect 106885 -8360 106926 -8326
rect 108219 -8333 108220 -8322
rect 108396 -8327 108459 -8293
rect 108468 -8327 108503 -8293
rect 108580 -8327 108615 -8293
rect 109111 -8317 109146 -8283
rect 109207 -8317 109242 -8283
rect 109303 -8317 109338 -8283
rect 109399 -8317 109434 -8283
rect 109495 -8317 109530 -8283
rect 110520 -8324 110555 -8290
rect 110565 -8324 110566 -8279
rect 110665 -8290 110666 -8279
rect 110676 -8324 110711 -8290
rect 110721 -8324 110722 -8279
rect 110821 -8290 110822 -8279
rect 111000 -8284 111035 -8250
rect 111072 -8284 111107 -8250
rect 111144 -8284 111179 -8250
rect 111288 -8284 111323 -8250
rect 111360 -8284 111395 -8250
rect 111397 -8284 111467 -8250
rect 111504 -8284 111539 -8250
rect 111574 -8284 111609 -8250
rect 112101 -8274 112136 -8240
rect 112197 -8274 112232 -8240
rect 112293 -8274 112328 -8240
rect 113800 -8241 113835 -8207
rect 113864 -8241 113907 -8207
rect 113909 -8241 113910 -8199
rect 114009 -8207 114010 -8199
rect 113944 -8241 113979 -8207
rect 114020 -8241 114055 -8207
rect 114065 -8241 114066 -8199
rect 114165 -8207 114166 -8199
rect 114114 -8241 114149 -8207
rect 114176 -8241 114221 -8207
rect 115091 -8231 115126 -8197
rect 115187 -8231 115222 -8197
rect 115283 -8231 115318 -8197
rect 114907 -8250 114908 -8242
rect 110832 -8324 110867 -8290
rect 111813 -8293 111814 -8285
rect 111913 -8293 111914 -8285
rect 105230 -8410 105271 -8376
rect 105863 -8379 105870 -8371
rect 104880 -8451 104921 -8417
rect 104869 -8500 104876 -8489
rect 104880 -8500 104885 -8451
rect 105074 -8494 105115 -8460
rect 105119 -8494 105126 -8449
rect 105219 -8460 105226 -8449
rect 105428 -8453 105469 -8419
rect 105473 -8453 105480 -8408
rect 105573 -8419 105580 -8408
rect 105754 -8413 105795 -8379
rect 105818 -8413 105870 -8379
rect 105898 -8413 105939 -8379
rect 105584 -8453 105625 -8419
rect 105230 -8494 105271 -8460
rect 104880 -8534 104921 -8500
rect 104880 -8568 104885 -8534
rect 103530 -8740 103535 -8706
rect 103826 -8723 103867 -8689
rect 103871 -8723 103878 -8681
rect 104013 -8741 104025 -8673
rect 104054 -8707 104059 -8639
rect 104099 -8671 104104 -8603
rect 104133 -8637 104138 -8571
rect 105074 -8577 105115 -8543
rect 105119 -8577 105126 -8532
rect 105219 -8543 105226 -8532
rect 105428 -8537 105469 -8503
rect 105473 -8537 105480 -8492
rect 105573 -8503 105580 -8492
rect 105818 -8496 105859 -8462
rect 105863 -8496 105870 -8451
rect 105584 -8537 105625 -8503
rect 105230 -8577 105271 -8543
rect 104143 -8621 104184 -8587
rect 104344 -8666 104385 -8632
rect 104113 -8689 104120 -8681
rect 104124 -8723 104165 -8689
rect 104344 -8734 104385 -8700
rect 101277 -8906 101318 -8872
rect 101349 -8906 101390 -8872
rect 101421 -8906 101462 -8872
rect 101734 -8913 101775 -8879
rect 101779 -8913 101786 -8868
rect 101879 -8879 101886 -8868
rect 101890 -8913 101931 -8879
rect 102474 -8895 102515 -8861
rect 102519 -8895 102526 -8853
rect 100368 -8959 100850 -8925
rect 101702 -8949 101743 -8915
rect 101774 -8949 101815 -8915
rect 102088 -8956 102129 -8922
rect 102133 -8956 102140 -8911
rect 102233 -8922 102240 -8911
rect 102661 -8913 102673 -8845
rect 102702 -8879 102707 -8811
rect 102747 -8843 102752 -8775
rect 102781 -8809 102786 -8743
rect 104013 -8753 104020 -8741
rect 104393 -8750 104398 -8616
rect 102791 -8793 102832 -8759
rect 102994 -8838 103035 -8804
rect 102761 -8861 102768 -8853
rect 102772 -8895 102813 -8861
rect 102994 -8906 103035 -8872
rect 102244 -8956 102285 -8922
rect 100368 -8985 100837 -8959
rect 100372 -8993 100579 -8985
rect 100388 -9003 100563 -8993
rect 100114 -9140 100295 -9114
rect 99621 -9174 99662 -9140
rect 99717 -9174 99758 -9140
rect 99813 -9174 99854 -9140
rect 99909 -9174 99950 -9140
rect 100005 -9174 100046 -9140
rect 100101 -9174 100295 -9140
rect 100114 -9200 100295 -9174
rect 100314 -9174 100421 -9050
rect 100573 -9062 100579 -9051
rect 100192 -9870 100233 -9200
rect 100314 -9228 100323 -9174
rect 99999 -9936 100150 -9924
rect 99667 -9970 100150 -9936
rect 99999 -9971 100150 -9970
rect 100180 -9971 100233 -9870
rect 100326 -9971 100367 -9174
rect 100372 -9971 100378 -9174
rect 100584 -9971 100625 -9062
rect 100718 -9971 100759 -8985
rect 100971 -9002 101012 -8968
rect 101067 -9002 101108 -8968
rect 101163 -9002 101204 -8968
rect 101259 -9002 101300 -8968
rect 101355 -9002 101396 -8968
rect 101451 -9002 101492 -8968
rect 101547 -9002 101588 -8968
rect 102056 -8992 102097 -8958
rect 102128 -8992 102169 -8958
rect 102474 -8995 102515 -8961
rect 102519 -8995 102526 -8950
rect 102661 -9001 102668 -8913
rect 103043 -8922 103048 -8788
rect 102761 -8961 102768 -8950
rect 103077 -8956 103082 -8762
rect 103117 -8778 103124 -8767
rect 103113 -8809 103124 -8778
rect 103439 -8796 103480 -8762
rect 102772 -8995 102813 -8961
rect 101709 -9045 101750 -9011
rect 101805 -9045 101846 -9011
rect 101901 -9045 101942 -9011
rect 102410 -9035 102451 -9001
rect 102482 -9035 102523 -9001
rect 102554 -9035 102595 -9001
rect 102626 -9029 102668 -9001
rect 102972 -9025 103013 -8991
rect 103017 -9025 103024 -8980
rect 103113 -8992 103118 -8809
rect 103147 -8995 103152 -8812
rect 102626 -9035 102667 -9029
rect 102063 -9088 102104 -9054
rect 102159 -9088 102200 -9054
rect 102255 -9088 102296 -9054
rect 103159 -9076 103166 -8809
rect 103788 -8819 104181 -8753
rect 104427 -8784 104432 -8590
rect 104467 -8606 104474 -8595
rect 104463 -8637 104474 -8606
rect 104789 -8624 104830 -8590
rect 103175 -8860 103216 -8826
rect 103524 -8830 103541 -8819
rect 103524 -8832 103530 -8830
rect 103175 -8928 103216 -8894
rect 103227 -8995 103232 -8860
rect 103458 -8874 103530 -8832
rect 103586 -8874 104181 -8819
rect 104322 -8853 104363 -8819
rect 104367 -8853 104374 -8808
rect 104463 -8820 104468 -8637
rect 104497 -8823 104502 -8640
rect 103458 -8877 104181 -8874
rect 103261 -8980 103266 -8892
rect 103378 -8942 103419 -8908
rect 103423 -8942 103430 -8900
rect 103259 -8991 103266 -8980
rect 103261 -9025 103266 -8991
rect 103270 -9025 103311 -8991
rect 103378 -9042 103419 -9008
rect 103423 -9042 103430 -8997
rect 103271 -9078 103312 -9044
rect 103343 -9078 103384 -9044
rect 103415 -9078 103456 -9044
rect 102417 -9131 102458 -9097
rect 102513 -9131 102554 -9097
rect 102609 -9131 102650 -9097
rect 102705 -9131 102746 -9097
rect 102801 -9131 102842 -9097
rect 103458 -9114 103609 -8877
rect 103788 -8899 104181 -8877
rect 103712 -8925 104181 -8899
rect 104509 -8904 104516 -8637
rect 104525 -8688 104566 -8654
rect 104525 -8756 104566 -8722
rect 104577 -8823 104582 -8688
rect 105139 -8691 105180 -8657
rect 105191 -8718 105196 -8641
rect 104611 -8808 104616 -8720
rect 104728 -8770 104769 -8736
rect 104773 -8770 104780 -8728
rect 104873 -8740 104880 -8729
rect 104884 -8774 104925 -8740
rect 105225 -8752 105230 -8607
rect 105428 -8620 105469 -8586
rect 105473 -8620 105480 -8575
rect 105573 -8586 105580 -8575
rect 105818 -8580 105859 -8546
rect 105863 -8580 105870 -8535
rect 105584 -8620 105625 -8586
rect 105493 -8734 105534 -8700
rect 105545 -8761 105550 -8684
rect 104609 -8819 104616 -8808
rect 105078 -8813 105119 -8779
rect 105123 -8813 105130 -8771
rect 105223 -8779 105230 -8771
rect 105234 -8813 105275 -8779
rect 105579 -8795 105584 -8650
rect 105818 -8663 105859 -8629
rect 105863 -8663 105870 -8618
rect 105940 -8679 105945 -8363
rect 105963 -8379 105970 -8371
rect 105974 -8379 105979 -8363
rect 105974 -8413 106015 -8379
rect 106019 -8413 106026 -8371
rect 105963 -8462 105970 -8451
rect 105974 -8462 105979 -8413
rect 105974 -8496 106015 -8462
rect 106019 -8496 106026 -8451
rect 105963 -8546 105970 -8535
rect 105974 -8546 105979 -8496
rect 105974 -8580 106015 -8546
rect 106019 -8580 106026 -8535
rect 105963 -8629 105970 -8618
rect 105974 -8629 105979 -8580
rect 105974 -8663 106015 -8629
rect 106019 -8663 106026 -8618
rect 105963 -8697 105970 -8671
rect 105974 -8713 105979 -8663
rect 105883 -8777 105924 -8743
rect 104611 -8853 104616 -8819
rect 104620 -8853 104661 -8819
rect 104728 -8870 104769 -8836
rect 104773 -8870 104780 -8825
rect 104873 -8832 104880 -8821
rect 104884 -8866 104925 -8832
rect 105432 -8856 105473 -8822
rect 105477 -8856 105484 -8814
rect 105577 -8822 105584 -8814
rect 105588 -8856 105629 -8822
rect 106005 -8845 106012 -8697
rect 106028 -8713 106031 -8363
rect 106062 -8679 106065 -8363
rect 106119 -8379 106126 -8371
rect 106068 -8413 106109 -8379
rect 106130 -8413 106181 -8379
rect 106840 -8422 106845 -8406
rect 106863 -8422 106870 -8414
rect 106874 -8422 106879 -8406
rect 107176 -8408 107211 -8374
rect 107221 -8408 107222 -8363
rect 107321 -8374 107322 -8363
rect 107332 -8408 107367 -8374
rect 107377 -8408 107378 -8363
rect 107477 -8374 107478 -8363
rect 108053 -8367 108088 -8333
rect 108230 -8367 108265 -8333
rect 108823 -8336 108824 -8328
rect 108923 -8336 108924 -8328
rect 107488 -8408 107523 -8374
rect 108219 -8417 108220 -8406
rect 108424 -8410 108459 -8376
rect 108469 -8410 108470 -8365
rect 108569 -8376 108570 -8365
rect 108750 -8370 108813 -8336
rect 108822 -8370 108857 -8336
rect 108934 -8370 108969 -8336
rect 109659 -8360 109694 -8326
rect 109755 -8360 109790 -8326
rect 109851 -8360 109886 -8326
rect 109947 -8360 109982 -8326
rect 110043 -8360 110078 -8326
rect 110139 -8360 110174 -8326
rect 110235 -8360 110270 -8326
rect 111563 -8333 111564 -8322
rect 111740 -8327 111803 -8293
rect 111812 -8327 111847 -8293
rect 111924 -8327 111959 -8293
rect 112455 -8317 112490 -8283
rect 112551 -8317 112586 -8283
rect 112647 -8317 112682 -8283
rect 112743 -8317 112778 -8283
rect 112839 -8317 112874 -8283
rect 113864 -8324 113899 -8290
rect 113909 -8324 113910 -8279
rect 114009 -8290 114010 -8279
rect 114020 -8324 114055 -8290
rect 114065 -8324 114066 -8279
rect 114165 -8290 114166 -8279
rect 114344 -8284 114379 -8250
rect 114416 -8284 114451 -8250
rect 114488 -8284 114523 -8250
rect 114632 -8284 114667 -8250
rect 114704 -8284 114739 -8250
rect 114741 -8284 114811 -8250
rect 114848 -8284 114883 -8250
rect 114918 -8284 114953 -8250
rect 115445 -8274 115480 -8240
rect 115541 -8274 115576 -8240
rect 115637 -8274 115672 -8240
rect 117144 -8241 117179 -8207
rect 117208 -8241 117251 -8207
rect 117253 -8241 117254 -8199
rect 117353 -8207 117354 -8199
rect 117288 -8241 117323 -8207
rect 117364 -8241 117399 -8207
rect 117409 -8241 117410 -8199
rect 117509 -8207 117510 -8199
rect 117458 -8241 117493 -8207
rect 117520 -8241 117565 -8207
rect 118435 -8231 118470 -8197
rect 118531 -8231 118566 -8197
rect 118627 -8231 118662 -8197
rect 118251 -8250 118252 -8242
rect 114176 -8324 114211 -8290
rect 115157 -8293 115158 -8285
rect 115257 -8293 115258 -8285
rect 108580 -8410 108615 -8376
rect 106119 -8462 106126 -8451
rect 106300 -8456 106341 -8422
rect 106372 -8456 106413 -8422
rect 106444 -8456 106485 -8422
rect 106588 -8456 106629 -8422
rect 106660 -8456 106773 -8422
rect 106804 -8456 106845 -8422
rect 106130 -8496 106171 -8462
rect 106119 -8546 106126 -8535
rect 106697 -8539 106738 -8505
rect 106130 -8580 106171 -8546
rect 106119 -8629 106126 -8618
rect 106130 -8663 106171 -8629
rect 106362 -8689 106403 -8655
rect 106407 -8689 106414 -8644
rect 106484 -8706 106489 -8588
rect 106507 -8655 106514 -8644
rect 106518 -8655 106523 -8622
rect 106554 -8655 106559 -8622
rect 106518 -8689 106559 -8655
rect 106563 -8689 106570 -8644
rect 106518 -8740 106523 -8689
rect 106554 -8740 106559 -8689
rect 106588 -8706 106593 -8589
rect 106697 -8623 106738 -8589
rect 106697 -8706 106738 -8672
rect 106840 -8706 106845 -8456
rect 106874 -8456 106915 -8422
rect 106863 -8505 106870 -8494
rect 106874 -8505 106879 -8456
rect 107176 -8491 107211 -8457
rect 107221 -8491 107222 -8446
rect 107321 -8457 107322 -8446
rect 107332 -8491 107367 -8457
rect 107377 -8491 107378 -8446
rect 107477 -8457 107478 -8446
rect 108053 -8451 108088 -8417
rect 108230 -8451 108265 -8417
rect 107488 -8491 107523 -8457
rect 106874 -8539 106915 -8505
rect 106863 -8589 106870 -8578
rect 106874 -8589 106879 -8539
rect 107023 -8565 107138 -8499
rect 107321 -8525 107322 -8499
rect 107718 -8517 107753 -8483
rect 107763 -8517 107764 -8472
rect 107863 -8483 107864 -8472
rect 107874 -8517 107909 -8483
rect 107919 -8517 107920 -8472
rect 108219 -8500 108220 -8489
rect 108424 -8494 108459 -8460
rect 108469 -8494 108470 -8449
rect 108569 -8460 108570 -8449
rect 108778 -8453 108813 -8419
rect 108823 -8453 108824 -8408
rect 108923 -8419 108924 -8408
rect 109104 -8413 109139 -8379
rect 109168 -8413 109211 -8379
rect 109213 -8413 109214 -8371
rect 109313 -8379 109314 -8371
rect 109248 -8413 109283 -8379
rect 109324 -8413 109359 -8379
rect 109369 -8413 109370 -8371
rect 109469 -8379 109470 -8371
rect 109418 -8413 109453 -8379
rect 109480 -8413 109525 -8379
rect 110520 -8408 110555 -8374
rect 110565 -8408 110566 -8363
rect 110665 -8374 110666 -8363
rect 110676 -8408 110711 -8374
rect 110721 -8408 110722 -8363
rect 110821 -8374 110822 -8363
rect 111397 -8367 111432 -8333
rect 111574 -8367 111609 -8333
rect 112167 -8336 112168 -8328
rect 112267 -8336 112268 -8328
rect 110832 -8408 110867 -8374
rect 108934 -8453 108969 -8419
rect 110213 -8422 110214 -8414
rect 111563 -8417 111564 -8406
rect 111768 -8410 111803 -8376
rect 111813 -8410 111814 -8365
rect 111913 -8376 111914 -8365
rect 112094 -8370 112157 -8336
rect 112166 -8370 112201 -8336
rect 112278 -8370 112313 -8336
rect 113003 -8360 113038 -8326
rect 113099 -8360 113134 -8326
rect 113195 -8360 113230 -8326
rect 113291 -8360 113326 -8326
rect 113387 -8360 113422 -8326
rect 113483 -8360 113518 -8326
rect 113579 -8360 113614 -8326
rect 114907 -8333 114908 -8322
rect 115084 -8327 115147 -8293
rect 115156 -8327 115191 -8293
rect 115268 -8327 115303 -8293
rect 115799 -8317 115834 -8283
rect 115895 -8317 115930 -8283
rect 115991 -8317 116026 -8283
rect 116087 -8317 116122 -8283
rect 116183 -8317 116218 -8283
rect 117208 -8324 117243 -8290
rect 117253 -8324 117254 -8279
rect 117353 -8290 117354 -8279
rect 117364 -8324 117399 -8290
rect 117409 -8324 117410 -8279
rect 117509 -8290 117510 -8279
rect 117688 -8284 117723 -8250
rect 117760 -8284 117795 -8250
rect 117832 -8284 117867 -8250
rect 117976 -8284 118011 -8250
rect 118048 -8284 118083 -8250
rect 118085 -8284 118155 -8250
rect 118192 -8284 118227 -8250
rect 118262 -8284 118297 -8250
rect 118789 -8274 118824 -8240
rect 118885 -8274 118920 -8240
rect 118981 -8274 119016 -8240
rect 120488 -8241 120523 -8207
rect 120552 -8241 120595 -8207
rect 120597 -8241 120598 -8199
rect 120697 -8207 120698 -8199
rect 120632 -8241 120667 -8207
rect 120708 -8241 120743 -8207
rect 120753 -8241 120754 -8199
rect 120853 -8207 120854 -8199
rect 120802 -8241 120837 -8207
rect 120864 -8241 120909 -8207
rect 121779 -8231 121814 -8197
rect 121875 -8231 121910 -8197
rect 121971 -8231 122006 -8197
rect 121595 -8250 121596 -8242
rect 117520 -8324 117555 -8290
rect 118501 -8293 118502 -8285
rect 118601 -8293 118602 -8285
rect 111924 -8410 111959 -8376
rect 108580 -8494 108615 -8460
rect 106874 -8623 106915 -8589
rect 107241 -8605 107276 -8571
rect 106863 -8672 106870 -8661
rect 106874 -8672 106879 -8623
rect 106874 -8706 106915 -8672
rect 106874 -8740 106879 -8706
rect 107176 -8723 107211 -8689
rect 107221 -8723 107222 -8681
rect 104621 -8906 104662 -8872
rect 104693 -8906 104734 -8872
rect 104765 -8906 104806 -8872
rect 105078 -8913 105119 -8879
rect 105123 -8913 105130 -8868
rect 105223 -8879 105230 -8868
rect 105234 -8913 105275 -8879
rect 105818 -8895 105859 -8861
rect 105863 -8895 105870 -8853
rect 103712 -8959 104194 -8925
rect 105046 -8949 105087 -8915
rect 105118 -8949 105159 -8915
rect 105432 -8956 105473 -8922
rect 105477 -8956 105484 -8911
rect 105577 -8922 105584 -8911
rect 106005 -8913 106017 -8845
rect 106046 -8879 106051 -8811
rect 106091 -8843 106096 -8775
rect 106125 -8809 106130 -8743
rect 107363 -8753 107364 -8525
rect 108053 -8534 108088 -8500
rect 108230 -8534 108265 -8500
rect 108424 -8577 108459 -8543
rect 108469 -8577 108470 -8532
rect 108569 -8543 108570 -8532
rect 108778 -8537 108813 -8503
rect 108823 -8537 108824 -8492
rect 108923 -8503 108924 -8492
rect 109168 -8496 109203 -8462
rect 109213 -8496 109214 -8451
rect 109313 -8462 109314 -8451
rect 109324 -8496 109359 -8462
rect 109369 -8496 109370 -8451
rect 109469 -8462 109470 -8451
rect 109650 -8456 109685 -8422
rect 109722 -8456 109757 -8422
rect 109794 -8456 109829 -8422
rect 109938 -8456 109973 -8422
rect 110010 -8456 110045 -8422
rect 110047 -8456 110117 -8422
rect 110154 -8456 110189 -8422
rect 110224 -8456 110259 -8422
rect 109480 -8496 109515 -8462
rect 110520 -8491 110555 -8457
rect 110565 -8491 110566 -8446
rect 110665 -8457 110666 -8446
rect 110676 -8491 110711 -8457
rect 110721 -8491 110722 -8446
rect 110821 -8457 110822 -8446
rect 111397 -8451 111432 -8417
rect 111574 -8451 111609 -8417
rect 110832 -8491 110867 -8457
rect 108934 -8537 108969 -8503
rect 110213 -8505 110214 -8494
rect 108580 -8577 108615 -8543
rect 107493 -8621 107528 -8587
rect 107694 -8666 107729 -8632
rect 107817 -8637 107818 -8595
rect 108139 -8624 108174 -8590
rect 108778 -8620 108813 -8586
rect 108823 -8620 108824 -8575
rect 108923 -8586 108924 -8575
rect 109168 -8580 109203 -8546
rect 109213 -8580 109214 -8535
rect 109313 -8546 109314 -8535
rect 109324 -8580 109359 -8546
rect 109369 -8580 109370 -8535
rect 109469 -8546 109470 -8535
rect 110047 -8539 110082 -8505
rect 110224 -8539 110259 -8505
rect 109480 -8580 109515 -8546
rect 110367 -8565 110482 -8499
rect 110665 -8525 110666 -8499
rect 111062 -8517 111097 -8483
rect 111107 -8517 111108 -8472
rect 111207 -8483 111208 -8472
rect 111218 -8517 111253 -8483
rect 111263 -8517 111264 -8472
rect 111563 -8500 111564 -8489
rect 111768 -8494 111803 -8460
rect 111813 -8494 111814 -8449
rect 111913 -8460 111914 -8449
rect 112122 -8453 112157 -8419
rect 112167 -8453 112168 -8408
rect 112267 -8419 112268 -8408
rect 112448 -8413 112483 -8379
rect 112512 -8413 112555 -8379
rect 112557 -8413 112558 -8371
rect 112657 -8379 112658 -8371
rect 112592 -8413 112627 -8379
rect 112668 -8413 112703 -8379
rect 112713 -8413 112714 -8371
rect 112813 -8379 112814 -8371
rect 112762 -8413 112797 -8379
rect 112824 -8413 112869 -8379
rect 113864 -8408 113899 -8374
rect 113909 -8408 113910 -8363
rect 114009 -8374 114010 -8363
rect 114020 -8408 114055 -8374
rect 114065 -8408 114066 -8363
rect 114165 -8374 114166 -8363
rect 114741 -8367 114776 -8333
rect 114918 -8367 114953 -8333
rect 115511 -8336 115512 -8328
rect 115611 -8336 115612 -8328
rect 114176 -8408 114211 -8374
rect 112278 -8453 112313 -8419
rect 113557 -8422 113558 -8414
rect 114907 -8417 114908 -8406
rect 115112 -8410 115147 -8376
rect 115157 -8410 115158 -8365
rect 115257 -8376 115258 -8365
rect 115438 -8370 115501 -8336
rect 115510 -8370 115545 -8336
rect 115622 -8370 115657 -8336
rect 116347 -8360 116382 -8326
rect 116443 -8360 116478 -8326
rect 116539 -8360 116574 -8326
rect 116635 -8360 116670 -8326
rect 116731 -8360 116766 -8326
rect 116827 -8360 116862 -8326
rect 116923 -8360 116958 -8326
rect 118251 -8333 118252 -8322
rect 118428 -8327 118491 -8293
rect 118500 -8327 118535 -8293
rect 118612 -8327 118647 -8293
rect 119143 -8317 119178 -8283
rect 119239 -8317 119274 -8283
rect 119335 -8317 119370 -8283
rect 119431 -8317 119466 -8283
rect 119527 -8317 119562 -8283
rect 120552 -8324 120587 -8290
rect 120597 -8324 120598 -8279
rect 120697 -8290 120698 -8279
rect 120708 -8324 120743 -8290
rect 120753 -8324 120754 -8279
rect 120853 -8290 120854 -8279
rect 121032 -8284 121067 -8250
rect 121104 -8284 121139 -8250
rect 121176 -8284 121211 -8250
rect 121320 -8284 121355 -8250
rect 121392 -8284 121427 -8250
rect 121429 -8284 121499 -8250
rect 121536 -8284 121571 -8250
rect 121606 -8284 121641 -8250
rect 122133 -8274 122168 -8240
rect 122229 -8274 122264 -8240
rect 122325 -8274 122360 -8240
rect 123832 -8241 123867 -8207
rect 123896 -8241 123939 -8207
rect 123941 -8241 123942 -8199
rect 124041 -8207 124042 -8199
rect 123976 -8241 124011 -8207
rect 124052 -8241 124087 -8207
rect 124097 -8241 124098 -8199
rect 124197 -8207 124198 -8199
rect 124146 -8241 124181 -8207
rect 124208 -8241 124253 -8207
rect 125123 -8231 125158 -8197
rect 125219 -8231 125254 -8197
rect 125315 -8231 125350 -8197
rect 124939 -8250 124940 -8242
rect 120864 -8324 120899 -8290
rect 121845 -8293 121846 -8285
rect 121945 -8293 121946 -8285
rect 115268 -8410 115303 -8376
rect 111924 -8494 111959 -8460
rect 108934 -8620 108969 -8586
rect 110213 -8589 110214 -8578
rect 107463 -8689 107464 -8681
rect 107474 -8723 107509 -8689
rect 107694 -8734 107729 -8700
rect 106135 -8793 106176 -8759
rect 106338 -8838 106379 -8804
rect 106105 -8861 106112 -8853
rect 106116 -8895 106157 -8861
rect 106338 -8906 106379 -8872
rect 105588 -8956 105629 -8922
rect 103712 -8985 104181 -8959
rect 103716 -8993 103923 -8985
rect 103732 -9003 103907 -8993
rect 103458 -9140 103639 -9114
rect 102965 -9174 103006 -9140
rect 103061 -9174 103102 -9140
rect 103157 -9174 103198 -9140
rect 103253 -9174 103294 -9140
rect 103349 -9174 103390 -9140
rect 103445 -9174 103639 -9140
rect 103458 -9200 103639 -9174
rect 103658 -9174 103765 -9050
rect 103917 -9062 103923 -9051
rect 103536 -9870 103577 -9200
rect 103658 -9228 103667 -9174
rect 103343 -9936 103494 -9924
rect 103011 -9970 103494 -9936
rect 103343 -9971 103494 -9970
rect 103524 -9971 103577 -9870
rect 103670 -9971 103711 -9174
rect 103716 -9971 103722 -9174
rect 103928 -9971 103969 -9062
rect 104062 -9971 104103 -8985
rect 104315 -9002 104356 -8968
rect 104411 -9002 104452 -8968
rect 104507 -9002 104548 -8968
rect 104603 -9002 104644 -8968
rect 104699 -9002 104740 -8968
rect 104795 -9002 104836 -8968
rect 104891 -9002 104932 -8968
rect 105400 -8992 105441 -8958
rect 105472 -8992 105513 -8958
rect 105818 -8995 105859 -8961
rect 105863 -8995 105870 -8950
rect 106005 -9001 106012 -8913
rect 106387 -8922 106392 -8788
rect 106105 -8961 106112 -8950
rect 106421 -8956 106426 -8762
rect 106461 -8778 106468 -8767
rect 106457 -8809 106468 -8778
rect 106783 -8796 106824 -8762
rect 106116 -8995 106157 -8961
rect 105053 -9045 105094 -9011
rect 105149 -9045 105190 -9011
rect 105245 -9045 105286 -9011
rect 105754 -9035 105795 -9001
rect 105826 -9035 105867 -9001
rect 105898 -9035 105939 -9001
rect 105970 -9029 106012 -9001
rect 106316 -9025 106357 -8991
rect 106361 -9025 106368 -8980
rect 106457 -8992 106462 -8809
rect 106491 -8995 106496 -8812
rect 105970 -9035 106011 -9029
rect 105407 -9088 105448 -9054
rect 105503 -9088 105544 -9054
rect 105599 -9088 105640 -9054
rect 106503 -9076 106510 -8809
rect 107138 -8819 107525 -8753
rect 106519 -8860 106560 -8826
rect 106868 -8830 106885 -8819
rect 106868 -8832 106874 -8830
rect 106519 -8928 106560 -8894
rect 106571 -8995 106576 -8860
rect 106802 -8874 106874 -8832
rect 106936 -8874 107525 -8819
rect 107672 -8853 107707 -8819
rect 107717 -8853 107718 -8808
rect 106802 -8877 107525 -8874
rect 106605 -8980 106610 -8892
rect 106722 -8942 106763 -8908
rect 106767 -8942 106774 -8900
rect 106603 -8991 106610 -8980
rect 106605 -9025 106610 -8991
rect 106614 -9025 106655 -8991
rect 106722 -9042 106763 -9008
rect 106767 -9042 106774 -8997
rect 106615 -9078 106656 -9044
rect 106687 -9078 106728 -9044
rect 106759 -9078 106800 -9044
rect 105761 -9131 105802 -9097
rect 105857 -9131 105898 -9097
rect 105953 -9131 105994 -9097
rect 106049 -9131 106090 -9097
rect 106145 -9131 106186 -9097
rect 106802 -9114 106953 -8877
rect 107138 -8899 107525 -8877
rect 107062 -8925 107525 -8899
rect 107859 -8904 107860 -8637
rect 107875 -8688 107910 -8654
rect 108489 -8691 108524 -8657
rect 109168 -8663 109203 -8629
rect 109213 -8663 109214 -8618
rect 109313 -8629 109314 -8618
rect 109324 -8663 109359 -8629
rect 109369 -8663 109370 -8618
rect 109469 -8629 109470 -8618
rect 110047 -8623 110082 -8589
rect 110224 -8623 110259 -8589
rect 110585 -8605 110620 -8571
rect 109480 -8663 109515 -8629
rect 109313 -8697 109314 -8671
rect 109712 -8689 109747 -8655
rect 109757 -8689 109758 -8644
rect 109857 -8655 109858 -8644
rect 109868 -8689 109903 -8655
rect 109913 -8689 109914 -8644
rect 110213 -8672 110214 -8661
rect 107875 -8756 107910 -8722
rect 108078 -8770 108113 -8736
rect 108123 -8770 108124 -8728
rect 108223 -8740 108224 -8729
rect 108843 -8734 108878 -8700
rect 108234 -8774 108269 -8740
rect 107959 -8819 107960 -8808
rect 108428 -8813 108463 -8779
rect 108473 -8813 108474 -8771
rect 108573 -8779 108574 -8771
rect 109233 -8777 109268 -8743
rect 108584 -8813 108619 -8779
rect 107970 -8853 108005 -8819
rect 108078 -8870 108113 -8836
rect 108123 -8870 108124 -8825
rect 108223 -8832 108224 -8821
rect 108234 -8866 108269 -8832
rect 108782 -8856 108817 -8822
rect 108827 -8856 108828 -8814
rect 108927 -8822 108928 -8814
rect 108938 -8856 108973 -8822
rect 107971 -8906 108006 -8872
rect 108043 -8906 108078 -8872
rect 108115 -8906 108150 -8872
rect 108428 -8913 108463 -8879
rect 108473 -8913 108474 -8868
rect 108573 -8879 108574 -8868
rect 108584 -8913 108619 -8879
rect 109168 -8895 109203 -8861
rect 109213 -8895 109214 -8853
rect 107062 -8959 107538 -8925
rect 108396 -8949 108431 -8915
rect 108468 -8949 108503 -8915
rect 108782 -8956 108817 -8922
rect 108827 -8956 108828 -8911
rect 108927 -8922 108928 -8911
rect 108938 -8956 108973 -8922
rect 107062 -8969 107525 -8959
rect 107060 -8985 107525 -8969
rect 107060 -8993 107267 -8985
rect 107076 -9003 107251 -8993
rect 106802 -9140 106983 -9114
rect 106309 -9174 106350 -9140
rect 106405 -9174 106446 -9140
rect 106501 -9174 106542 -9140
rect 106597 -9174 106638 -9140
rect 106693 -9174 106734 -9140
rect 106789 -9174 106983 -9140
rect 106802 -9200 106983 -9174
rect 107002 -9174 107109 -9050
rect 107261 -9062 107267 -9051
rect 106880 -9870 106921 -9200
rect 107002 -9228 107011 -9174
rect 106687 -9936 106838 -9924
rect 106355 -9970 106838 -9936
rect 106687 -9971 106838 -9970
rect 106868 -9971 106921 -9870
rect 107014 -9971 107055 -9174
rect 107060 -9971 107066 -9174
rect 107272 -9971 107313 -9062
rect 107406 -9971 107447 -8985
rect 107665 -9002 107700 -8968
rect 107761 -9002 107796 -8968
rect 107857 -9002 107892 -8968
rect 107953 -9002 107988 -8968
rect 108049 -9002 108084 -8968
rect 108145 -9002 108180 -8968
rect 108241 -9002 108276 -8968
rect 108750 -8992 108785 -8958
rect 108822 -8992 108857 -8958
rect 109168 -8995 109203 -8961
rect 109213 -8995 109214 -8950
rect 109355 -9001 109356 -8697
rect 110047 -8706 110082 -8672
rect 110224 -8706 110259 -8672
rect 110520 -8723 110555 -8689
rect 110565 -8723 110566 -8681
rect 110707 -8753 110708 -8525
rect 111397 -8534 111432 -8500
rect 111574 -8534 111609 -8500
rect 111768 -8577 111803 -8543
rect 111813 -8577 111814 -8532
rect 111913 -8543 111914 -8532
rect 112122 -8537 112157 -8503
rect 112167 -8537 112168 -8492
rect 112267 -8503 112268 -8492
rect 112512 -8496 112547 -8462
rect 112557 -8496 112558 -8451
rect 112657 -8462 112658 -8451
rect 112668 -8496 112703 -8462
rect 112713 -8496 112714 -8451
rect 112813 -8462 112814 -8451
rect 112994 -8456 113029 -8422
rect 113066 -8456 113101 -8422
rect 113138 -8456 113173 -8422
rect 113282 -8456 113317 -8422
rect 113354 -8456 113389 -8422
rect 113391 -8456 113461 -8422
rect 113498 -8456 113533 -8422
rect 113568 -8456 113603 -8422
rect 112824 -8496 112859 -8462
rect 113864 -8491 113899 -8457
rect 113909 -8491 113910 -8446
rect 114009 -8457 114010 -8446
rect 114020 -8491 114055 -8457
rect 114065 -8491 114066 -8446
rect 114165 -8457 114166 -8446
rect 114741 -8451 114776 -8417
rect 114918 -8451 114953 -8417
rect 114176 -8491 114211 -8457
rect 112278 -8537 112313 -8503
rect 113557 -8505 113558 -8494
rect 111924 -8577 111959 -8543
rect 110837 -8621 110872 -8587
rect 111038 -8666 111073 -8632
rect 111161 -8637 111162 -8595
rect 111483 -8624 111518 -8590
rect 112122 -8620 112157 -8586
rect 112167 -8620 112168 -8575
rect 112267 -8586 112268 -8575
rect 112512 -8580 112547 -8546
rect 112557 -8580 112558 -8535
rect 112657 -8546 112658 -8535
rect 112668 -8580 112703 -8546
rect 112713 -8580 112714 -8535
rect 112813 -8546 112814 -8535
rect 113391 -8539 113426 -8505
rect 113568 -8539 113603 -8505
rect 112824 -8580 112859 -8546
rect 113711 -8565 113826 -8499
rect 114009 -8525 114010 -8499
rect 114406 -8517 114441 -8483
rect 114451 -8517 114452 -8472
rect 114551 -8483 114552 -8472
rect 114562 -8517 114597 -8483
rect 114607 -8517 114608 -8472
rect 114907 -8500 114908 -8489
rect 115112 -8494 115147 -8460
rect 115157 -8494 115158 -8449
rect 115257 -8460 115258 -8449
rect 115466 -8453 115501 -8419
rect 115511 -8453 115512 -8408
rect 115611 -8419 115612 -8408
rect 115792 -8413 115827 -8379
rect 115856 -8413 115899 -8379
rect 115901 -8413 115902 -8371
rect 116001 -8379 116002 -8371
rect 115936 -8413 115971 -8379
rect 116012 -8413 116047 -8379
rect 116057 -8413 116058 -8371
rect 116157 -8379 116158 -8371
rect 116106 -8413 116141 -8379
rect 116168 -8413 116213 -8379
rect 117208 -8408 117243 -8374
rect 117253 -8408 117254 -8363
rect 117353 -8374 117354 -8363
rect 117364 -8408 117399 -8374
rect 117409 -8408 117410 -8363
rect 117509 -8374 117510 -8363
rect 118085 -8367 118120 -8333
rect 118262 -8367 118297 -8333
rect 118855 -8336 118856 -8328
rect 118955 -8336 118956 -8328
rect 117520 -8408 117555 -8374
rect 115622 -8453 115657 -8419
rect 116901 -8422 116902 -8414
rect 118251 -8417 118252 -8406
rect 118456 -8410 118491 -8376
rect 118501 -8410 118502 -8365
rect 118601 -8376 118602 -8365
rect 118782 -8370 118845 -8336
rect 118854 -8370 118889 -8336
rect 118966 -8370 119001 -8336
rect 119691 -8360 119726 -8326
rect 119787 -8360 119822 -8326
rect 119883 -8360 119918 -8326
rect 119979 -8360 120014 -8326
rect 120075 -8360 120110 -8326
rect 120171 -8360 120206 -8326
rect 120267 -8360 120302 -8326
rect 121595 -8333 121596 -8322
rect 121772 -8327 121835 -8293
rect 121844 -8327 121879 -8293
rect 121956 -8327 121991 -8293
rect 122487 -8317 122522 -8283
rect 122583 -8317 122618 -8283
rect 122679 -8317 122714 -8283
rect 122775 -8317 122810 -8283
rect 122871 -8317 122906 -8283
rect 123896 -8324 123931 -8290
rect 123941 -8324 123942 -8279
rect 124041 -8290 124042 -8279
rect 124052 -8324 124087 -8290
rect 124097 -8324 124098 -8279
rect 124197 -8290 124198 -8279
rect 124376 -8284 124411 -8250
rect 124448 -8284 124483 -8250
rect 124520 -8284 124555 -8250
rect 124664 -8284 124699 -8250
rect 124736 -8284 124771 -8250
rect 124773 -8284 124843 -8250
rect 124880 -8284 124915 -8250
rect 124950 -8284 124985 -8250
rect 125477 -8274 125512 -8240
rect 125573 -8274 125608 -8240
rect 125669 -8274 125704 -8240
rect 127176 -8241 127211 -8207
rect 127240 -8241 127283 -8207
rect 127285 -8241 127286 -8199
rect 127385 -8207 127386 -8199
rect 127320 -8241 127355 -8207
rect 127396 -8241 127431 -8207
rect 127441 -8241 127442 -8199
rect 127541 -8207 127542 -8199
rect 127490 -8241 127525 -8207
rect 127552 -8241 127597 -8207
rect 128467 -8231 128502 -8197
rect 128563 -8231 128598 -8197
rect 128659 -8231 128694 -8197
rect 128283 -8250 128284 -8242
rect 124208 -8324 124243 -8290
rect 125189 -8293 125190 -8285
rect 125289 -8293 125290 -8285
rect 118612 -8410 118647 -8376
rect 115268 -8494 115303 -8460
rect 112278 -8620 112313 -8586
rect 113557 -8589 113558 -8578
rect 110807 -8689 110808 -8681
rect 110818 -8723 110853 -8689
rect 111038 -8734 111073 -8700
rect 109485 -8793 109520 -8759
rect 109688 -8838 109723 -8804
rect 109811 -8809 109812 -8767
rect 110133 -8796 110168 -8762
rect 109455 -8861 109456 -8853
rect 109466 -8895 109501 -8861
rect 109688 -8906 109723 -8872
rect 109455 -8961 109456 -8950
rect 109466 -8995 109501 -8961
rect 108403 -9045 108438 -9011
rect 108499 -9045 108534 -9011
rect 108595 -9045 108630 -9011
rect 109104 -9035 109139 -9001
rect 109176 -9035 109211 -9001
rect 109248 -9035 109283 -9001
rect 109320 -9029 109356 -9001
rect 109666 -9025 109701 -8991
rect 109711 -9025 109712 -8980
rect 109320 -9035 109355 -9029
rect 108757 -9088 108792 -9054
rect 108853 -9088 108888 -9054
rect 108949 -9088 108984 -9054
rect 109853 -9076 109854 -8809
rect 110482 -8819 110869 -8753
rect 109869 -8860 109904 -8826
rect 110218 -8832 110229 -8819
rect 110152 -8874 110229 -8832
rect 110280 -8874 110869 -8819
rect 111016 -8853 111051 -8819
rect 111061 -8853 111062 -8808
rect 110152 -8877 110869 -8874
rect 109869 -8928 109904 -8894
rect 110072 -8942 110107 -8908
rect 110117 -8942 110118 -8900
rect 109953 -8991 109954 -8980
rect 109964 -9025 109999 -8991
rect 110072 -9042 110107 -9008
rect 110117 -9042 110118 -8997
rect 109965 -9078 110000 -9044
rect 110037 -9078 110072 -9044
rect 110109 -9078 110144 -9044
rect 109111 -9131 109146 -9097
rect 109207 -9131 109242 -9097
rect 109303 -9131 109338 -9097
rect 109399 -9131 109434 -9097
rect 109495 -9131 109530 -9097
rect 110152 -9114 110297 -8877
rect 110482 -8899 110869 -8877
rect 110406 -8925 110869 -8899
rect 111203 -8904 111204 -8637
rect 111219 -8688 111254 -8654
rect 111833 -8691 111868 -8657
rect 112512 -8663 112547 -8629
rect 112557 -8663 112558 -8618
rect 112657 -8629 112658 -8618
rect 112668 -8663 112703 -8629
rect 112713 -8663 112714 -8618
rect 112813 -8629 112814 -8618
rect 113391 -8623 113426 -8589
rect 113568 -8623 113603 -8589
rect 113929 -8605 113964 -8571
rect 112824 -8663 112859 -8629
rect 112657 -8697 112658 -8671
rect 113056 -8689 113091 -8655
rect 113101 -8689 113102 -8644
rect 113201 -8655 113202 -8644
rect 113212 -8689 113247 -8655
rect 113257 -8689 113258 -8644
rect 113557 -8672 113558 -8661
rect 111219 -8756 111254 -8722
rect 111422 -8770 111457 -8736
rect 111467 -8770 111468 -8728
rect 111567 -8740 111568 -8729
rect 112187 -8734 112222 -8700
rect 111578 -8774 111613 -8740
rect 111303 -8819 111304 -8808
rect 111772 -8813 111807 -8779
rect 111817 -8813 111818 -8771
rect 111917 -8779 111918 -8771
rect 112577 -8777 112612 -8743
rect 111928 -8813 111963 -8779
rect 111314 -8853 111349 -8819
rect 111422 -8870 111457 -8836
rect 111467 -8870 111468 -8825
rect 111567 -8832 111568 -8821
rect 111578 -8866 111613 -8832
rect 112126 -8856 112161 -8822
rect 112171 -8856 112172 -8814
rect 112271 -8822 112272 -8814
rect 112282 -8856 112317 -8822
rect 111315 -8906 111350 -8872
rect 111387 -8906 111422 -8872
rect 111459 -8906 111494 -8872
rect 111772 -8913 111807 -8879
rect 111817 -8913 111818 -8868
rect 111917 -8879 111918 -8868
rect 111928 -8913 111963 -8879
rect 112512 -8895 112547 -8861
rect 112557 -8895 112558 -8853
rect 110406 -8959 110882 -8925
rect 111740 -8949 111775 -8915
rect 111812 -8949 111847 -8915
rect 112126 -8956 112161 -8922
rect 112171 -8956 112172 -8911
rect 112271 -8922 112272 -8911
rect 112282 -8956 112317 -8922
rect 110406 -8985 110869 -8959
rect 110410 -8993 110611 -8985
rect 110426 -9003 110595 -8993
rect 110152 -9140 110327 -9114
rect 109659 -9174 109694 -9140
rect 109755 -9174 109790 -9140
rect 109851 -9174 109886 -9140
rect 109947 -9174 109982 -9140
rect 110043 -9174 110078 -9140
rect 110139 -9174 110327 -9140
rect 110152 -9200 110327 -9174
rect 110352 -9174 110453 -9050
rect 110230 -9870 110265 -9200
rect 110352 -9228 110355 -9174
rect 110037 -9936 110182 -9924
rect 109705 -9970 110182 -9936
rect 110037 -9971 110182 -9970
rect 110218 -9971 110265 -9870
rect 110364 -9971 110399 -9174
rect 110622 -9971 110657 -9062
rect 110756 -9971 110791 -8985
rect 111009 -9002 111044 -8968
rect 111105 -9002 111140 -8968
rect 111201 -9002 111236 -8968
rect 111297 -9002 111332 -8968
rect 111393 -9002 111428 -8968
rect 111489 -9002 111524 -8968
rect 111585 -9002 111620 -8968
rect 112094 -8992 112129 -8958
rect 112166 -8992 112201 -8958
rect 112512 -8995 112547 -8961
rect 112557 -8995 112558 -8950
rect 112699 -9001 112700 -8697
rect 113391 -8706 113426 -8672
rect 113568 -8706 113603 -8672
rect 113864 -8723 113899 -8689
rect 113909 -8723 113910 -8681
rect 114051 -8753 114052 -8525
rect 114741 -8534 114776 -8500
rect 114918 -8534 114953 -8500
rect 115112 -8577 115147 -8543
rect 115157 -8577 115158 -8532
rect 115257 -8543 115258 -8532
rect 115466 -8537 115501 -8503
rect 115511 -8537 115512 -8492
rect 115611 -8503 115612 -8492
rect 115856 -8496 115891 -8462
rect 115901 -8496 115902 -8451
rect 116001 -8462 116002 -8451
rect 116012 -8496 116047 -8462
rect 116057 -8496 116058 -8451
rect 116157 -8462 116158 -8451
rect 116338 -8456 116373 -8422
rect 116410 -8456 116445 -8422
rect 116482 -8456 116517 -8422
rect 116626 -8456 116661 -8422
rect 116698 -8456 116733 -8422
rect 116735 -8456 116805 -8422
rect 116842 -8456 116877 -8422
rect 116912 -8456 116947 -8422
rect 116168 -8496 116203 -8462
rect 117208 -8491 117243 -8457
rect 117253 -8491 117254 -8446
rect 117353 -8457 117354 -8446
rect 117364 -8491 117399 -8457
rect 117409 -8491 117410 -8446
rect 117509 -8457 117510 -8446
rect 118085 -8451 118120 -8417
rect 118262 -8451 118297 -8417
rect 117520 -8491 117555 -8457
rect 115622 -8537 115657 -8503
rect 116901 -8505 116902 -8494
rect 115268 -8577 115303 -8543
rect 114181 -8621 114216 -8587
rect 114382 -8666 114417 -8632
rect 114505 -8637 114506 -8595
rect 114827 -8624 114862 -8590
rect 115466 -8620 115501 -8586
rect 115511 -8620 115512 -8575
rect 115611 -8586 115612 -8575
rect 115856 -8580 115891 -8546
rect 115901 -8580 115902 -8535
rect 116001 -8546 116002 -8535
rect 116012 -8580 116047 -8546
rect 116057 -8580 116058 -8535
rect 116157 -8546 116158 -8535
rect 116735 -8539 116770 -8505
rect 116912 -8539 116947 -8505
rect 116168 -8580 116203 -8546
rect 117055 -8565 117170 -8499
rect 117353 -8525 117354 -8499
rect 117750 -8517 117785 -8483
rect 117795 -8517 117796 -8472
rect 117895 -8483 117896 -8472
rect 117906 -8517 117941 -8483
rect 117951 -8517 117952 -8472
rect 118251 -8500 118252 -8489
rect 118456 -8494 118491 -8460
rect 118501 -8494 118502 -8449
rect 118601 -8460 118602 -8449
rect 118810 -8453 118845 -8419
rect 118855 -8453 118856 -8408
rect 118955 -8419 118956 -8408
rect 119136 -8413 119171 -8379
rect 119200 -8413 119243 -8379
rect 119245 -8413 119246 -8371
rect 119345 -8379 119346 -8371
rect 119280 -8413 119315 -8379
rect 119356 -8413 119391 -8379
rect 119401 -8413 119402 -8371
rect 119501 -8379 119502 -8371
rect 119450 -8413 119485 -8379
rect 119512 -8413 119557 -8379
rect 120552 -8408 120587 -8374
rect 120597 -8408 120598 -8363
rect 120697 -8374 120698 -8363
rect 120708 -8408 120743 -8374
rect 120753 -8408 120754 -8363
rect 120853 -8374 120854 -8363
rect 121429 -8367 121464 -8333
rect 121606 -8367 121641 -8333
rect 122199 -8336 122200 -8328
rect 122299 -8336 122300 -8328
rect 120864 -8408 120899 -8374
rect 118966 -8453 119001 -8419
rect 120245 -8422 120246 -8414
rect 121595 -8417 121596 -8406
rect 121800 -8410 121835 -8376
rect 121845 -8410 121846 -8365
rect 121945 -8376 121946 -8365
rect 122126 -8370 122189 -8336
rect 122198 -8370 122233 -8336
rect 122310 -8370 122345 -8336
rect 123035 -8360 123070 -8326
rect 123131 -8360 123166 -8326
rect 123227 -8360 123262 -8326
rect 123323 -8360 123358 -8326
rect 123419 -8360 123454 -8326
rect 123515 -8360 123550 -8326
rect 123611 -8360 123646 -8326
rect 124939 -8333 124940 -8322
rect 125116 -8327 125179 -8293
rect 125188 -8327 125223 -8293
rect 125300 -8327 125335 -8293
rect 125831 -8317 125866 -8283
rect 125927 -8317 125962 -8283
rect 126023 -8317 126058 -8283
rect 126119 -8317 126154 -8283
rect 126215 -8317 126250 -8283
rect 127240 -8324 127275 -8290
rect 127285 -8324 127286 -8279
rect 127385 -8290 127386 -8279
rect 127396 -8324 127431 -8290
rect 127441 -8324 127442 -8279
rect 127541 -8290 127542 -8279
rect 127720 -8284 127755 -8250
rect 127792 -8284 127827 -8250
rect 127864 -8284 127899 -8250
rect 128008 -8284 128043 -8250
rect 128080 -8284 128115 -8250
rect 128117 -8284 128187 -8250
rect 128224 -8284 128259 -8250
rect 128294 -8284 128329 -8250
rect 128821 -8274 128856 -8240
rect 128917 -8274 128952 -8240
rect 129013 -8274 129048 -8240
rect 130520 -8241 130555 -8207
rect 130584 -8241 130627 -8207
rect 130629 -8241 130630 -8199
rect 130729 -8207 130730 -8199
rect 130664 -8241 130699 -8207
rect 130740 -8241 130775 -8207
rect 130785 -8241 130786 -8199
rect 130885 -8207 130886 -8199
rect 130834 -8241 130869 -8207
rect 130896 -8241 130941 -8207
rect 131811 -8231 131846 -8197
rect 131907 -8231 131942 -8197
rect 132003 -8231 132038 -8197
rect 131627 -8250 131628 -8242
rect 127552 -8324 127587 -8290
rect 128533 -8293 128534 -8285
rect 128633 -8293 128634 -8285
rect 121956 -8410 121991 -8376
rect 118612 -8494 118647 -8460
rect 115622 -8620 115657 -8586
rect 116901 -8589 116902 -8578
rect 114151 -8689 114152 -8681
rect 114162 -8723 114197 -8689
rect 114382 -8734 114417 -8700
rect 112829 -8793 112864 -8759
rect 113032 -8838 113067 -8804
rect 113155 -8809 113156 -8767
rect 113477 -8796 113512 -8762
rect 112799 -8861 112800 -8853
rect 112810 -8895 112845 -8861
rect 113032 -8906 113067 -8872
rect 112799 -8961 112800 -8950
rect 112810 -8995 112845 -8961
rect 111747 -9045 111782 -9011
rect 111843 -9045 111878 -9011
rect 111939 -9045 111974 -9011
rect 112448 -9035 112483 -9001
rect 112520 -9035 112555 -9001
rect 112592 -9035 112627 -9001
rect 112664 -9029 112700 -9001
rect 113010 -9025 113045 -8991
rect 113055 -9025 113056 -8980
rect 112664 -9035 112699 -9029
rect 112101 -9088 112136 -9054
rect 112197 -9088 112232 -9054
rect 112293 -9088 112328 -9054
rect 113197 -9076 113198 -8809
rect 113826 -8819 114213 -8753
rect 113213 -8860 113248 -8826
rect 113562 -8832 113573 -8819
rect 113496 -8874 113573 -8832
rect 113624 -8874 114213 -8819
rect 114360 -8853 114395 -8819
rect 114405 -8853 114406 -8808
rect 113496 -8877 114213 -8874
rect 113213 -8928 113248 -8894
rect 113416 -8942 113451 -8908
rect 113461 -8942 113462 -8900
rect 113297 -8991 113298 -8980
rect 113308 -9025 113343 -8991
rect 113416 -9042 113451 -9008
rect 113461 -9042 113462 -8997
rect 113309 -9078 113344 -9044
rect 113381 -9078 113416 -9044
rect 113453 -9078 113488 -9044
rect 112455 -9131 112490 -9097
rect 112551 -9131 112586 -9097
rect 112647 -9131 112682 -9097
rect 112743 -9131 112778 -9097
rect 112839 -9131 112874 -9097
rect 113496 -9114 113641 -8877
rect 113826 -8899 114213 -8877
rect 113750 -8925 114213 -8899
rect 114547 -8904 114548 -8637
rect 114563 -8688 114598 -8654
rect 115177 -8691 115212 -8657
rect 115856 -8663 115891 -8629
rect 115901 -8663 115902 -8618
rect 116001 -8629 116002 -8618
rect 116012 -8663 116047 -8629
rect 116057 -8663 116058 -8618
rect 116157 -8629 116158 -8618
rect 116735 -8623 116770 -8589
rect 116912 -8623 116947 -8589
rect 117273 -8605 117308 -8571
rect 116168 -8663 116203 -8629
rect 116001 -8697 116002 -8671
rect 116400 -8689 116435 -8655
rect 116445 -8689 116446 -8644
rect 116545 -8655 116546 -8644
rect 116556 -8689 116591 -8655
rect 116601 -8689 116602 -8644
rect 116901 -8672 116902 -8661
rect 114563 -8756 114598 -8722
rect 114766 -8770 114801 -8736
rect 114811 -8770 114812 -8728
rect 114911 -8740 114912 -8729
rect 115531 -8734 115566 -8700
rect 114922 -8774 114957 -8740
rect 114647 -8819 114648 -8808
rect 115116 -8813 115151 -8779
rect 115161 -8813 115162 -8771
rect 115261 -8779 115262 -8771
rect 115921 -8777 115956 -8743
rect 115272 -8813 115307 -8779
rect 114658 -8853 114693 -8819
rect 114766 -8870 114801 -8836
rect 114811 -8870 114812 -8825
rect 114911 -8832 114912 -8821
rect 114922 -8866 114957 -8832
rect 115470 -8856 115505 -8822
rect 115515 -8856 115516 -8814
rect 115615 -8822 115616 -8814
rect 115626 -8856 115661 -8822
rect 114659 -8906 114694 -8872
rect 114731 -8906 114766 -8872
rect 114803 -8906 114838 -8872
rect 115116 -8913 115151 -8879
rect 115161 -8913 115162 -8868
rect 115261 -8879 115262 -8868
rect 115272 -8913 115307 -8879
rect 115856 -8895 115891 -8861
rect 115901 -8895 115902 -8853
rect 113750 -8959 114226 -8925
rect 115084 -8949 115119 -8915
rect 115156 -8949 115191 -8915
rect 115470 -8956 115505 -8922
rect 115515 -8956 115516 -8911
rect 115615 -8922 115616 -8911
rect 115626 -8956 115661 -8922
rect 113750 -8985 114213 -8959
rect 113754 -8993 113955 -8985
rect 113770 -9003 113939 -8993
rect 113496 -9140 113671 -9114
rect 113003 -9174 113038 -9140
rect 113099 -9174 113134 -9140
rect 113195 -9174 113230 -9140
rect 113291 -9174 113326 -9140
rect 113387 -9174 113422 -9140
rect 113483 -9174 113671 -9140
rect 113496 -9200 113671 -9174
rect 113696 -9174 113797 -9050
rect 113574 -9870 113609 -9200
rect 113696 -9228 113699 -9174
rect 113381 -9936 113526 -9924
rect 113049 -9970 113526 -9936
rect 113381 -9971 113526 -9970
rect 113562 -9971 113609 -9870
rect 113708 -9971 113743 -9174
rect 113966 -9971 114001 -9062
rect 114100 -9971 114135 -8985
rect 114353 -9002 114388 -8968
rect 114449 -9002 114484 -8968
rect 114545 -9002 114580 -8968
rect 114641 -9002 114676 -8968
rect 114737 -9002 114772 -8968
rect 114833 -9002 114868 -8968
rect 114929 -9002 114964 -8968
rect 115438 -8992 115473 -8958
rect 115510 -8992 115545 -8958
rect 115856 -8995 115891 -8961
rect 115901 -8995 115902 -8950
rect 116043 -9001 116044 -8697
rect 116735 -8706 116770 -8672
rect 116912 -8706 116947 -8672
rect 117208 -8723 117243 -8689
rect 117253 -8723 117254 -8681
rect 117395 -8753 117396 -8525
rect 118085 -8534 118120 -8500
rect 118262 -8534 118297 -8500
rect 118456 -8577 118491 -8543
rect 118501 -8577 118502 -8532
rect 118601 -8543 118602 -8532
rect 118810 -8537 118845 -8503
rect 118855 -8537 118856 -8492
rect 118955 -8503 118956 -8492
rect 119200 -8496 119235 -8462
rect 119245 -8496 119246 -8451
rect 119345 -8462 119346 -8451
rect 119356 -8496 119391 -8462
rect 119401 -8496 119402 -8451
rect 119501 -8462 119502 -8451
rect 119682 -8456 119717 -8422
rect 119754 -8456 119789 -8422
rect 119826 -8456 119861 -8422
rect 119970 -8456 120005 -8422
rect 120042 -8456 120077 -8422
rect 120079 -8456 120149 -8422
rect 120186 -8456 120221 -8422
rect 120256 -8456 120291 -8422
rect 119512 -8496 119547 -8462
rect 120552 -8491 120587 -8457
rect 120597 -8491 120598 -8446
rect 120697 -8457 120698 -8446
rect 120708 -8491 120743 -8457
rect 120753 -8491 120754 -8446
rect 120853 -8457 120854 -8446
rect 121429 -8451 121464 -8417
rect 121606 -8451 121641 -8417
rect 120864 -8491 120899 -8457
rect 118966 -8537 119001 -8503
rect 120245 -8505 120246 -8494
rect 118612 -8577 118647 -8543
rect 117525 -8621 117560 -8587
rect 117726 -8666 117761 -8632
rect 117849 -8637 117850 -8595
rect 118171 -8624 118206 -8590
rect 118810 -8620 118845 -8586
rect 118855 -8620 118856 -8575
rect 118955 -8586 118956 -8575
rect 119200 -8580 119235 -8546
rect 119245 -8580 119246 -8535
rect 119345 -8546 119346 -8535
rect 119356 -8580 119391 -8546
rect 119401 -8580 119402 -8535
rect 119501 -8546 119502 -8535
rect 120079 -8539 120114 -8505
rect 120256 -8539 120291 -8505
rect 119512 -8580 119547 -8546
rect 120399 -8565 120514 -8499
rect 120697 -8525 120698 -8499
rect 121094 -8517 121129 -8483
rect 121139 -8517 121140 -8472
rect 121239 -8483 121240 -8472
rect 121250 -8517 121285 -8483
rect 121295 -8517 121296 -8472
rect 121595 -8500 121596 -8489
rect 121800 -8494 121835 -8460
rect 121845 -8494 121846 -8449
rect 121945 -8460 121946 -8449
rect 122154 -8453 122189 -8419
rect 122199 -8453 122200 -8408
rect 122299 -8419 122300 -8408
rect 122480 -8413 122515 -8379
rect 122544 -8413 122587 -8379
rect 122589 -8413 122590 -8371
rect 122689 -8379 122690 -8371
rect 122624 -8413 122659 -8379
rect 122700 -8413 122735 -8379
rect 122745 -8413 122746 -8371
rect 122845 -8379 122846 -8371
rect 122794 -8413 122829 -8379
rect 122856 -8413 122901 -8379
rect 123896 -8408 123931 -8374
rect 123941 -8408 123942 -8363
rect 124041 -8374 124042 -8363
rect 124052 -8408 124087 -8374
rect 124097 -8408 124098 -8363
rect 124197 -8374 124198 -8363
rect 124773 -8367 124808 -8333
rect 124950 -8367 124985 -8333
rect 125543 -8336 125544 -8328
rect 125643 -8336 125644 -8328
rect 124208 -8408 124243 -8374
rect 122310 -8453 122345 -8419
rect 123589 -8422 123590 -8414
rect 124939 -8417 124940 -8406
rect 125144 -8410 125179 -8376
rect 125189 -8410 125190 -8365
rect 125289 -8376 125290 -8365
rect 125470 -8370 125533 -8336
rect 125542 -8370 125577 -8336
rect 125654 -8370 125689 -8336
rect 126379 -8360 126414 -8326
rect 126475 -8360 126510 -8326
rect 126571 -8360 126606 -8326
rect 126667 -8360 126702 -8326
rect 126763 -8360 126798 -8326
rect 126859 -8360 126894 -8326
rect 126955 -8360 126990 -8326
rect 128283 -8333 128284 -8322
rect 128460 -8327 128523 -8293
rect 128532 -8327 128567 -8293
rect 128644 -8327 128679 -8293
rect 129175 -8317 129210 -8283
rect 129271 -8317 129306 -8283
rect 129367 -8317 129402 -8283
rect 129463 -8317 129498 -8283
rect 129559 -8317 129594 -8283
rect 130584 -8324 130619 -8290
rect 130629 -8324 130630 -8279
rect 130729 -8290 130730 -8279
rect 130740 -8324 130775 -8290
rect 130785 -8324 130786 -8279
rect 130885 -8290 130886 -8279
rect 131064 -8284 131099 -8250
rect 131136 -8284 131171 -8250
rect 131208 -8284 131243 -8250
rect 131352 -8284 131387 -8250
rect 131424 -8284 131459 -8250
rect 131461 -8284 131531 -8250
rect 131568 -8284 131603 -8250
rect 131638 -8284 131673 -8250
rect 132165 -8274 132200 -8240
rect 132261 -8274 132296 -8240
rect 132357 -8274 132392 -8240
rect 133864 -8241 133899 -8207
rect 133928 -8241 133971 -8207
rect 133973 -8241 133974 -8199
rect 134073 -8207 134074 -8199
rect 134008 -8241 134043 -8207
rect 134084 -8241 134119 -8207
rect 134129 -8241 134130 -8199
rect 134229 -8207 134230 -8199
rect 134178 -8241 134213 -8207
rect 134240 -8241 134285 -8207
rect 135155 -8231 135190 -8197
rect 135251 -8231 135286 -8197
rect 135347 -8231 135382 -8197
rect 134971 -8250 134972 -8242
rect 130896 -8324 130931 -8290
rect 131877 -8293 131878 -8285
rect 131977 -8293 131978 -8285
rect 125300 -8410 125335 -8376
rect 121956 -8494 121991 -8460
rect 118966 -8620 119001 -8586
rect 120245 -8589 120246 -8578
rect 117495 -8689 117496 -8681
rect 117506 -8723 117541 -8689
rect 117726 -8734 117761 -8700
rect 116173 -8793 116208 -8759
rect 116376 -8838 116411 -8804
rect 116499 -8809 116500 -8767
rect 116821 -8796 116856 -8762
rect 116143 -8861 116144 -8853
rect 116154 -8895 116189 -8861
rect 116376 -8906 116411 -8872
rect 116143 -8961 116144 -8950
rect 116154 -8995 116189 -8961
rect 115091 -9045 115126 -9011
rect 115187 -9045 115222 -9011
rect 115283 -9045 115318 -9011
rect 115792 -9035 115827 -9001
rect 115864 -9035 115899 -9001
rect 115936 -9035 115971 -9001
rect 116008 -9029 116044 -9001
rect 116354 -9025 116389 -8991
rect 116399 -9025 116400 -8980
rect 116008 -9035 116043 -9029
rect 115445 -9088 115480 -9054
rect 115541 -9088 115576 -9054
rect 115637 -9088 115672 -9054
rect 116541 -9076 116542 -8809
rect 117170 -8819 117557 -8753
rect 116557 -8860 116592 -8826
rect 116906 -8832 116917 -8819
rect 116840 -8874 116917 -8832
rect 116968 -8874 117557 -8819
rect 117704 -8853 117739 -8819
rect 117749 -8853 117750 -8808
rect 116840 -8877 117557 -8874
rect 116557 -8928 116592 -8894
rect 116760 -8942 116795 -8908
rect 116805 -8942 116806 -8900
rect 116641 -8991 116642 -8980
rect 116652 -9025 116687 -8991
rect 116760 -9042 116795 -9008
rect 116805 -9042 116806 -8997
rect 116653 -9078 116688 -9044
rect 116725 -9078 116760 -9044
rect 116797 -9078 116832 -9044
rect 115799 -9131 115834 -9097
rect 115895 -9131 115930 -9097
rect 115991 -9131 116026 -9097
rect 116087 -9131 116122 -9097
rect 116183 -9131 116218 -9097
rect 116840 -9114 116985 -8877
rect 117170 -8899 117557 -8877
rect 117094 -8925 117557 -8899
rect 117891 -8904 117892 -8637
rect 117907 -8688 117942 -8654
rect 118521 -8691 118556 -8657
rect 119200 -8663 119235 -8629
rect 119245 -8663 119246 -8618
rect 119345 -8629 119346 -8618
rect 119356 -8663 119391 -8629
rect 119401 -8663 119402 -8618
rect 119501 -8629 119502 -8618
rect 120079 -8623 120114 -8589
rect 120256 -8623 120291 -8589
rect 120617 -8605 120652 -8571
rect 119512 -8663 119547 -8629
rect 119345 -8697 119346 -8671
rect 119744 -8689 119779 -8655
rect 119789 -8689 119790 -8644
rect 119889 -8655 119890 -8644
rect 119900 -8689 119935 -8655
rect 119945 -8689 119946 -8644
rect 120245 -8672 120246 -8661
rect 117907 -8756 117942 -8722
rect 118110 -8770 118145 -8736
rect 118155 -8770 118156 -8728
rect 118255 -8740 118256 -8729
rect 118875 -8734 118910 -8700
rect 118266 -8774 118301 -8740
rect 117991 -8819 117992 -8808
rect 118460 -8813 118495 -8779
rect 118505 -8813 118506 -8771
rect 118605 -8779 118606 -8771
rect 119265 -8777 119300 -8743
rect 118616 -8813 118651 -8779
rect 118002 -8853 118037 -8819
rect 118110 -8870 118145 -8836
rect 118155 -8870 118156 -8825
rect 118255 -8832 118256 -8821
rect 118266 -8866 118301 -8832
rect 118814 -8856 118849 -8822
rect 118859 -8856 118860 -8814
rect 118959 -8822 118960 -8814
rect 118970 -8856 119005 -8822
rect 118003 -8906 118038 -8872
rect 118075 -8906 118110 -8872
rect 118147 -8906 118182 -8872
rect 118460 -8913 118495 -8879
rect 118505 -8913 118506 -8868
rect 118605 -8879 118606 -8868
rect 118616 -8913 118651 -8879
rect 119200 -8895 119235 -8861
rect 119245 -8895 119246 -8853
rect 117094 -8959 117570 -8925
rect 118428 -8949 118463 -8915
rect 118500 -8949 118535 -8915
rect 118814 -8956 118849 -8922
rect 118859 -8956 118860 -8911
rect 118959 -8922 118960 -8911
rect 118970 -8956 119005 -8922
rect 117094 -8985 117557 -8959
rect 117098 -8993 117299 -8985
rect 117114 -9003 117283 -8993
rect 116840 -9140 117015 -9114
rect 116347 -9174 116382 -9140
rect 116443 -9174 116478 -9140
rect 116539 -9174 116574 -9140
rect 116635 -9174 116670 -9140
rect 116731 -9174 116766 -9140
rect 116827 -9174 117015 -9140
rect 116840 -9200 117015 -9174
rect 117040 -9174 117141 -9050
rect 116918 -9870 116953 -9200
rect 117040 -9228 117043 -9174
rect 116725 -9936 116870 -9924
rect 116393 -9970 116870 -9936
rect 116725 -9971 116870 -9970
rect 116906 -9971 116953 -9870
rect 117052 -9971 117087 -9174
rect 117310 -9971 117345 -9062
rect 117444 -9971 117479 -8985
rect 117697 -9002 117732 -8968
rect 117793 -9002 117828 -8968
rect 117889 -9002 117924 -8968
rect 117985 -9002 118020 -8968
rect 118081 -9002 118116 -8968
rect 118177 -9002 118212 -8968
rect 118273 -9002 118308 -8968
rect 118782 -8992 118817 -8958
rect 118854 -8992 118889 -8958
rect 119200 -8995 119235 -8961
rect 119245 -8995 119246 -8950
rect 119387 -9001 119388 -8697
rect 120079 -8706 120114 -8672
rect 120256 -8706 120291 -8672
rect 120552 -8723 120587 -8689
rect 120597 -8723 120598 -8681
rect 120739 -8753 120740 -8525
rect 121429 -8534 121464 -8500
rect 121606 -8534 121641 -8500
rect 121800 -8577 121835 -8543
rect 121845 -8577 121846 -8532
rect 121945 -8543 121946 -8532
rect 122154 -8537 122189 -8503
rect 122199 -8537 122200 -8492
rect 122299 -8503 122300 -8492
rect 122544 -8496 122579 -8462
rect 122589 -8496 122590 -8451
rect 122689 -8462 122690 -8451
rect 122700 -8496 122735 -8462
rect 122745 -8496 122746 -8451
rect 122845 -8462 122846 -8451
rect 123026 -8456 123061 -8422
rect 123098 -8456 123133 -8422
rect 123170 -8456 123205 -8422
rect 123314 -8456 123349 -8422
rect 123386 -8456 123421 -8422
rect 123423 -8456 123493 -8422
rect 123530 -8456 123565 -8422
rect 123600 -8456 123635 -8422
rect 122856 -8496 122891 -8462
rect 123896 -8491 123931 -8457
rect 123941 -8491 123942 -8446
rect 124041 -8457 124042 -8446
rect 124052 -8491 124087 -8457
rect 124097 -8491 124098 -8446
rect 124197 -8457 124198 -8446
rect 124773 -8451 124808 -8417
rect 124950 -8451 124985 -8417
rect 124208 -8491 124243 -8457
rect 122310 -8537 122345 -8503
rect 123589 -8505 123590 -8494
rect 121956 -8577 121991 -8543
rect 120869 -8621 120904 -8587
rect 121070 -8666 121105 -8632
rect 121193 -8637 121194 -8595
rect 121515 -8624 121550 -8590
rect 122154 -8620 122189 -8586
rect 122199 -8620 122200 -8575
rect 122299 -8586 122300 -8575
rect 122544 -8580 122579 -8546
rect 122589 -8580 122590 -8535
rect 122689 -8546 122690 -8535
rect 122700 -8580 122735 -8546
rect 122745 -8580 122746 -8535
rect 122845 -8546 122846 -8535
rect 123423 -8539 123458 -8505
rect 123600 -8539 123635 -8505
rect 122856 -8580 122891 -8546
rect 123743 -8565 123858 -8499
rect 124041 -8525 124042 -8499
rect 124438 -8517 124473 -8483
rect 124483 -8517 124484 -8472
rect 124583 -8483 124584 -8472
rect 124594 -8517 124629 -8483
rect 124639 -8517 124640 -8472
rect 124939 -8500 124940 -8489
rect 125144 -8494 125179 -8460
rect 125189 -8494 125190 -8449
rect 125289 -8460 125290 -8449
rect 125498 -8453 125533 -8419
rect 125543 -8453 125544 -8408
rect 125643 -8419 125644 -8408
rect 125824 -8413 125859 -8379
rect 125888 -8413 125931 -8379
rect 125933 -8413 125934 -8371
rect 126033 -8379 126034 -8371
rect 125968 -8413 126003 -8379
rect 126044 -8413 126079 -8379
rect 126089 -8413 126090 -8371
rect 126189 -8379 126190 -8371
rect 126138 -8413 126173 -8379
rect 126200 -8413 126245 -8379
rect 127240 -8408 127275 -8374
rect 127285 -8408 127286 -8363
rect 127385 -8374 127386 -8363
rect 127396 -8408 127431 -8374
rect 127441 -8408 127442 -8363
rect 127541 -8374 127542 -8363
rect 128117 -8367 128152 -8333
rect 128294 -8367 128329 -8333
rect 128887 -8336 128888 -8328
rect 128987 -8336 128988 -8328
rect 127552 -8408 127587 -8374
rect 125654 -8453 125689 -8419
rect 126933 -8422 126934 -8414
rect 128283 -8417 128284 -8406
rect 128488 -8410 128523 -8376
rect 128533 -8410 128534 -8365
rect 128633 -8376 128634 -8365
rect 128814 -8370 128877 -8336
rect 128886 -8370 128921 -8336
rect 128998 -8370 129033 -8336
rect 129723 -8360 129758 -8326
rect 129819 -8360 129854 -8326
rect 129915 -8360 129950 -8326
rect 130011 -8360 130046 -8326
rect 130107 -8360 130142 -8326
rect 130203 -8360 130238 -8326
rect 130299 -8360 130334 -8326
rect 131627 -8333 131628 -8322
rect 131804 -8327 131867 -8293
rect 131876 -8327 131911 -8293
rect 131988 -8327 132023 -8293
rect 132519 -8317 132554 -8283
rect 132615 -8317 132650 -8283
rect 132711 -8317 132746 -8283
rect 132807 -8317 132842 -8283
rect 132903 -8317 132938 -8283
rect 133928 -8324 133963 -8290
rect 133973 -8324 133974 -8279
rect 134073 -8290 134074 -8279
rect 134084 -8324 134119 -8290
rect 134129 -8324 134130 -8279
rect 134229 -8290 134230 -8279
rect 134408 -8284 134443 -8250
rect 134480 -8284 134515 -8250
rect 134552 -8284 134587 -8250
rect 134696 -8284 134731 -8250
rect 134768 -8284 134803 -8250
rect 134805 -8284 134875 -8250
rect 134912 -8284 134947 -8250
rect 134982 -8284 135017 -8250
rect 135509 -8274 135544 -8240
rect 135605 -8274 135640 -8240
rect 135701 -8274 135736 -8240
rect 137208 -8241 137243 -8207
rect 137272 -8241 137315 -8207
rect 137317 -8241 137318 -8199
rect 137417 -8207 137418 -8199
rect 137352 -8241 137387 -8207
rect 137428 -8241 137463 -8207
rect 137473 -8241 137474 -8199
rect 137573 -8207 137574 -8199
rect 137522 -8241 137557 -8207
rect 137584 -8241 137629 -8207
rect 138499 -8231 138534 -8197
rect 138595 -8231 138630 -8197
rect 138691 -8231 138726 -8197
rect 138315 -8250 138316 -8242
rect 134240 -8324 134275 -8290
rect 135221 -8293 135222 -8285
rect 135321 -8293 135322 -8285
rect 128644 -8410 128679 -8376
rect 125300 -8494 125335 -8460
rect 122310 -8620 122345 -8586
rect 123589 -8589 123590 -8578
rect 120839 -8689 120840 -8681
rect 120850 -8723 120885 -8689
rect 121070 -8734 121105 -8700
rect 119517 -8793 119552 -8759
rect 119720 -8838 119755 -8804
rect 119843 -8809 119844 -8767
rect 120165 -8796 120200 -8762
rect 119487 -8861 119488 -8853
rect 119498 -8895 119533 -8861
rect 119720 -8906 119755 -8872
rect 119487 -8961 119488 -8950
rect 119498 -8995 119533 -8961
rect 118435 -9045 118470 -9011
rect 118531 -9045 118566 -9011
rect 118627 -9045 118662 -9011
rect 119136 -9035 119171 -9001
rect 119208 -9035 119243 -9001
rect 119280 -9035 119315 -9001
rect 119352 -9029 119388 -9001
rect 119698 -9025 119733 -8991
rect 119743 -9025 119744 -8980
rect 119352 -9035 119387 -9029
rect 118789 -9088 118824 -9054
rect 118885 -9088 118920 -9054
rect 118981 -9088 119016 -9054
rect 119885 -9076 119886 -8809
rect 120514 -8819 120901 -8753
rect 119901 -8860 119936 -8826
rect 120250 -8832 120261 -8819
rect 120184 -8874 120261 -8832
rect 120312 -8874 120901 -8819
rect 121048 -8853 121083 -8819
rect 121093 -8853 121094 -8808
rect 120184 -8877 120901 -8874
rect 119901 -8928 119936 -8894
rect 120104 -8942 120139 -8908
rect 120149 -8942 120150 -8900
rect 119985 -8991 119986 -8980
rect 119996 -9025 120031 -8991
rect 120104 -9042 120139 -9008
rect 120149 -9042 120150 -8997
rect 119997 -9078 120032 -9044
rect 120069 -9078 120104 -9044
rect 120141 -9078 120176 -9044
rect 119143 -9131 119178 -9097
rect 119239 -9131 119274 -9097
rect 119335 -9131 119370 -9097
rect 119431 -9131 119466 -9097
rect 119527 -9131 119562 -9097
rect 120184 -9114 120329 -8877
rect 120514 -8899 120901 -8877
rect 120438 -8925 120901 -8899
rect 121235 -8904 121236 -8637
rect 121251 -8688 121286 -8654
rect 121865 -8691 121900 -8657
rect 122544 -8663 122579 -8629
rect 122589 -8663 122590 -8618
rect 122689 -8629 122690 -8618
rect 122700 -8663 122735 -8629
rect 122745 -8663 122746 -8618
rect 122845 -8629 122846 -8618
rect 123423 -8623 123458 -8589
rect 123600 -8623 123635 -8589
rect 123961 -8605 123996 -8571
rect 122856 -8663 122891 -8629
rect 122689 -8697 122690 -8671
rect 123088 -8689 123123 -8655
rect 123133 -8689 123134 -8644
rect 123233 -8655 123234 -8644
rect 123244 -8689 123279 -8655
rect 123289 -8689 123290 -8644
rect 123589 -8672 123590 -8661
rect 121251 -8756 121286 -8722
rect 121454 -8770 121489 -8736
rect 121499 -8770 121500 -8728
rect 121599 -8740 121600 -8729
rect 122219 -8734 122254 -8700
rect 121610 -8774 121645 -8740
rect 121335 -8819 121336 -8808
rect 121804 -8813 121839 -8779
rect 121849 -8813 121850 -8771
rect 121949 -8779 121950 -8771
rect 122609 -8777 122644 -8743
rect 121960 -8813 121995 -8779
rect 121346 -8853 121381 -8819
rect 121454 -8870 121489 -8836
rect 121499 -8870 121500 -8825
rect 121599 -8832 121600 -8821
rect 121610 -8866 121645 -8832
rect 122158 -8856 122193 -8822
rect 122203 -8856 122204 -8814
rect 122303 -8822 122304 -8814
rect 122314 -8856 122349 -8822
rect 121347 -8906 121382 -8872
rect 121419 -8906 121454 -8872
rect 121491 -8906 121526 -8872
rect 121804 -8913 121839 -8879
rect 121849 -8913 121850 -8868
rect 121949 -8879 121950 -8868
rect 121960 -8913 121995 -8879
rect 122544 -8895 122579 -8861
rect 122589 -8895 122590 -8853
rect 120438 -8959 120914 -8925
rect 121772 -8949 121807 -8915
rect 121844 -8949 121879 -8915
rect 122158 -8956 122193 -8922
rect 122203 -8956 122204 -8911
rect 122303 -8922 122304 -8911
rect 122314 -8956 122349 -8922
rect 120438 -8985 120901 -8959
rect 120442 -8993 120643 -8985
rect 120458 -9003 120627 -8993
rect 120184 -9140 120359 -9114
rect 119691 -9174 119726 -9140
rect 119787 -9174 119822 -9140
rect 119883 -9174 119918 -9140
rect 119979 -9174 120014 -9140
rect 120075 -9174 120110 -9140
rect 120171 -9174 120359 -9140
rect 120184 -9200 120359 -9174
rect 120384 -9174 120485 -9050
rect 120262 -9870 120297 -9200
rect 120384 -9228 120387 -9174
rect 120069 -9936 120214 -9924
rect 119737 -9970 120214 -9936
rect 120069 -9971 120214 -9970
rect 120250 -9971 120297 -9870
rect 120396 -9971 120431 -9174
rect 120654 -9971 120689 -9062
rect 120788 -9971 120823 -8985
rect 121041 -9002 121076 -8968
rect 121137 -9002 121172 -8968
rect 121233 -9002 121268 -8968
rect 121329 -9002 121364 -8968
rect 121425 -9002 121460 -8968
rect 121521 -9002 121556 -8968
rect 121617 -9002 121652 -8968
rect 122126 -8992 122161 -8958
rect 122198 -8992 122233 -8958
rect 122544 -8995 122579 -8961
rect 122589 -8995 122590 -8950
rect 122731 -9001 122732 -8697
rect 123423 -8706 123458 -8672
rect 123600 -8706 123635 -8672
rect 123896 -8723 123931 -8689
rect 123941 -8723 123942 -8681
rect 124083 -8753 124084 -8525
rect 124773 -8534 124808 -8500
rect 124950 -8534 124985 -8500
rect 125144 -8577 125179 -8543
rect 125189 -8577 125190 -8532
rect 125289 -8543 125290 -8532
rect 125498 -8537 125533 -8503
rect 125543 -8537 125544 -8492
rect 125643 -8503 125644 -8492
rect 125888 -8496 125923 -8462
rect 125933 -8496 125934 -8451
rect 126033 -8462 126034 -8451
rect 126044 -8496 126079 -8462
rect 126089 -8496 126090 -8451
rect 126189 -8462 126190 -8451
rect 126370 -8456 126405 -8422
rect 126442 -8456 126477 -8422
rect 126514 -8456 126549 -8422
rect 126658 -8456 126693 -8422
rect 126730 -8456 126765 -8422
rect 126767 -8456 126837 -8422
rect 126874 -8456 126909 -8422
rect 126944 -8456 126979 -8422
rect 126200 -8496 126235 -8462
rect 127240 -8491 127275 -8457
rect 127285 -8491 127286 -8446
rect 127385 -8457 127386 -8446
rect 127396 -8491 127431 -8457
rect 127441 -8491 127442 -8446
rect 127541 -8457 127542 -8446
rect 128117 -8451 128152 -8417
rect 128294 -8451 128329 -8417
rect 127552 -8491 127587 -8457
rect 125654 -8537 125689 -8503
rect 126933 -8505 126934 -8494
rect 125300 -8577 125335 -8543
rect 124213 -8621 124248 -8587
rect 124414 -8666 124449 -8632
rect 124537 -8637 124538 -8595
rect 124859 -8624 124894 -8590
rect 125498 -8620 125533 -8586
rect 125543 -8620 125544 -8575
rect 125643 -8586 125644 -8575
rect 125888 -8580 125923 -8546
rect 125933 -8580 125934 -8535
rect 126033 -8546 126034 -8535
rect 126044 -8580 126079 -8546
rect 126089 -8580 126090 -8535
rect 126189 -8546 126190 -8535
rect 126767 -8539 126802 -8505
rect 126944 -8539 126979 -8505
rect 126200 -8580 126235 -8546
rect 127087 -8565 127202 -8499
rect 127385 -8525 127386 -8499
rect 127782 -8517 127817 -8483
rect 127827 -8517 127828 -8472
rect 127927 -8483 127928 -8472
rect 127938 -8517 127973 -8483
rect 127983 -8517 127984 -8472
rect 128283 -8500 128284 -8489
rect 128488 -8494 128523 -8460
rect 128533 -8494 128534 -8449
rect 128633 -8460 128634 -8449
rect 128842 -8453 128877 -8419
rect 128887 -8453 128888 -8408
rect 128987 -8419 128988 -8408
rect 129168 -8413 129203 -8379
rect 129232 -8413 129275 -8379
rect 129277 -8413 129278 -8371
rect 129377 -8379 129378 -8371
rect 129312 -8413 129347 -8379
rect 129388 -8413 129423 -8379
rect 129433 -8413 129434 -8371
rect 129533 -8379 129534 -8371
rect 129482 -8413 129517 -8379
rect 129544 -8413 129589 -8379
rect 130584 -8408 130619 -8374
rect 130629 -8408 130630 -8363
rect 130729 -8374 130730 -8363
rect 130740 -8408 130775 -8374
rect 130785 -8408 130786 -8363
rect 130885 -8374 130886 -8363
rect 131461 -8367 131496 -8333
rect 131638 -8367 131673 -8333
rect 132231 -8336 132232 -8328
rect 132331 -8336 132332 -8328
rect 130896 -8408 130931 -8374
rect 128998 -8453 129033 -8419
rect 130277 -8422 130278 -8414
rect 131627 -8417 131628 -8406
rect 131832 -8410 131867 -8376
rect 131877 -8410 131878 -8365
rect 131977 -8376 131978 -8365
rect 132158 -8370 132221 -8336
rect 132230 -8370 132265 -8336
rect 132342 -8370 132377 -8336
rect 133067 -8360 133102 -8326
rect 133163 -8360 133198 -8326
rect 133259 -8360 133294 -8326
rect 133355 -8360 133390 -8326
rect 133451 -8360 133486 -8326
rect 133547 -8360 133582 -8326
rect 133643 -8360 133678 -8326
rect 134971 -8333 134972 -8322
rect 135148 -8327 135211 -8293
rect 135220 -8327 135255 -8293
rect 135332 -8327 135367 -8293
rect 135863 -8317 135898 -8283
rect 135959 -8317 135994 -8283
rect 136055 -8317 136090 -8283
rect 136151 -8317 136186 -8283
rect 136247 -8317 136282 -8283
rect 137272 -8324 137307 -8290
rect 137317 -8324 137318 -8279
rect 137417 -8290 137418 -8279
rect 137428 -8324 137463 -8290
rect 137473 -8324 137474 -8279
rect 137573 -8290 137574 -8279
rect 137752 -8284 137787 -8250
rect 137824 -8284 137859 -8250
rect 137896 -8284 137931 -8250
rect 138040 -8284 138075 -8250
rect 138112 -8284 138147 -8250
rect 138149 -8284 138219 -8250
rect 138256 -8284 138291 -8250
rect 138326 -8284 138361 -8250
rect 138853 -8274 138888 -8240
rect 138949 -8274 138984 -8240
rect 139045 -8274 139080 -8240
rect 140552 -8241 140587 -8207
rect 140616 -8241 140659 -8207
rect 140661 -8241 140662 -8199
rect 140761 -8207 140762 -8199
rect 140696 -8241 140731 -8207
rect 140772 -8241 140807 -8207
rect 140817 -8241 140818 -8199
rect 140917 -8207 140918 -8199
rect 140866 -8241 140901 -8207
rect 140928 -8241 140973 -8207
rect 141843 -8231 141878 -8197
rect 141939 -8231 141974 -8197
rect 142035 -8231 142070 -8197
rect 141659 -8250 141660 -8242
rect 137584 -8324 137619 -8290
rect 138565 -8293 138566 -8285
rect 138665 -8293 138666 -8285
rect 131988 -8410 132023 -8376
rect 128644 -8494 128679 -8460
rect 125654 -8620 125689 -8586
rect 126933 -8589 126934 -8578
rect 124183 -8689 124184 -8681
rect 124194 -8723 124229 -8689
rect 124414 -8734 124449 -8700
rect 122861 -8793 122896 -8759
rect 123064 -8838 123099 -8804
rect 123187 -8809 123188 -8767
rect 123509 -8796 123544 -8762
rect 122831 -8861 122832 -8853
rect 122842 -8895 122877 -8861
rect 123064 -8906 123099 -8872
rect 122831 -8961 122832 -8950
rect 122842 -8995 122877 -8961
rect 121779 -9045 121814 -9011
rect 121875 -9045 121910 -9011
rect 121971 -9045 122006 -9011
rect 122480 -9035 122515 -9001
rect 122552 -9035 122587 -9001
rect 122624 -9035 122659 -9001
rect 122696 -9029 122732 -9001
rect 123042 -9025 123077 -8991
rect 123087 -9025 123088 -8980
rect 122696 -9035 122731 -9029
rect 122133 -9088 122168 -9054
rect 122229 -9088 122264 -9054
rect 122325 -9088 122360 -9054
rect 123229 -9076 123230 -8809
rect 123858 -8819 124245 -8753
rect 123245 -8860 123280 -8826
rect 123594 -8832 123605 -8819
rect 123528 -8874 123605 -8832
rect 123656 -8874 124245 -8819
rect 124392 -8853 124427 -8819
rect 124437 -8853 124438 -8808
rect 123528 -8877 124245 -8874
rect 123245 -8928 123280 -8894
rect 123448 -8942 123483 -8908
rect 123493 -8942 123494 -8900
rect 123329 -8991 123330 -8980
rect 123340 -9025 123375 -8991
rect 123448 -9042 123483 -9008
rect 123493 -9042 123494 -8997
rect 123341 -9078 123376 -9044
rect 123413 -9078 123448 -9044
rect 123485 -9078 123520 -9044
rect 122487 -9131 122522 -9097
rect 122583 -9131 122618 -9097
rect 122679 -9131 122714 -9097
rect 122775 -9131 122810 -9097
rect 122871 -9131 122906 -9097
rect 123528 -9114 123673 -8877
rect 123858 -8899 124245 -8877
rect 123782 -8925 124245 -8899
rect 124579 -8904 124580 -8637
rect 124595 -8688 124630 -8654
rect 125209 -8691 125244 -8657
rect 125888 -8663 125923 -8629
rect 125933 -8663 125934 -8618
rect 126033 -8629 126034 -8618
rect 126044 -8663 126079 -8629
rect 126089 -8663 126090 -8618
rect 126189 -8629 126190 -8618
rect 126767 -8623 126802 -8589
rect 126944 -8623 126979 -8589
rect 127305 -8605 127340 -8571
rect 126200 -8663 126235 -8629
rect 126033 -8697 126034 -8671
rect 126432 -8689 126467 -8655
rect 126477 -8689 126478 -8644
rect 126577 -8655 126578 -8644
rect 126588 -8689 126623 -8655
rect 126633 -8689 126634 -8644
rect 126933 -8672 126934 -8661
rect 124595 -8756 124630 -8722
rect 124798 -8770 124833 -8736
rect 124843 -8770 124844 -8728
rect 124943 -8740 124944 -8729
rect 125563 -8734 125598 -8700
rect 124954 -8774 124989 -8740
rect 124679 -8819 124680 -8808
rect 125148 -8813 125183 -8779
rect 125193 -8813 125194 -8771
rect 125293 -8779 125294 -8771
rect 125953 -8777 125988 -8743
rect 125304 -8813 125339 -8779
rect 124690 -8853 124725 -8819
rect 124798 -8870 124833 -8836
rect 124843 -8870 124844 -8825
rect 124943 -8832 124944 -8821
rect 124954 -8866 124989 -8832
rect 125502 -8856 125537 -8822
rect 125547 -8856 125548 -8814
rect 125647 -8822 125648 -8814
rect 125658 -8856 125693 -8822
rect 124691 -8906 124726 -8872
rect 124763 -8906 124798 -8872
rect 124835 -8906 124870 -8872
rect 125148 -8913 125183 -8879
rect 125193 -8913 125194 -8868
rect 125293 -8879 125294 -8868
rect 125304 -8913 125339 -8879
rect 125888 -8895 125923 -8861
rect 125933 -8895 125934 -8853
rect 123782 -8959 124258 -8925
rect 125116 -8949 125151 -8915
rect 125188 -8949 125223 -8915
rect 125502 -8956 125537 -8922
rect 125547 -8956 125548 -8911
rect 125647 -8922 125648 -8911
rect 125658 -8956 125693 -8922
rect 123782 -8985 124245 -8959
rect 123786 -8993 123987 -8985
rect 123802 -9003 123971 -8993
rect 123528 -9140 123703 -9114
rect 123035 -9174 123070 -9140
rect 123131 -9174 123166 -9140
rect 123227 -9174 123262 -9140
rect 123323 -9174 123358 -9140
rect 123419 -9174 123454 -9140
rect 123515 -9174 123703 -9140
rect 123528 -9200 123703 -9174
rect 123728 -9174 123829 -9050
rect 123606 -9870 123641 -9200
rect 123728 -9228 123731 -9174
rect 123413 -9936 123558 -9924
rect 123081 -9970 123558 -9936
rect 123413 -9971 123558 -9970
rect 123594 -9971 123641 -9870
rect 123740 -9971 123775 -9174
rect 123998 -9971 124033 -9062
rect 124132 -9971 124167 -8985
rect 124385 -9002 124420 -8968
rect 124481 -9002 124516 -8968
rect 124577 -9002 124612 -8968
rect 124673 -9002 124708 -8968
rect 124769 -9002 124804 -8968
rect 124865 -9002 124900 -8968
rect 124961 -9002 124996 -8968
rect 125470 -8992 125505 -8958
rect 125542 -8992 125577 -8958
rect 125888 -8995 125923 -8961
rect 125933 -8995 125934 -8950
rect 126075 -9001 126076 -8697
rect 126767 -8706 126802 -8672
rect 126944 -8706 126979 -8672
rect 127240 -8723 127275 -8689
rect 127285 -8723 127286 -8681
rect 127427 -8753 127428 -8525
rect 128117 -8534 128152 -8500
rect 128294 -8534 128329 -8500
rect 128488 -8577 128523 -8543
rect 128533 -8577 128534 -8532
rect 128633 -8543 128634 -8532
rect 128842 -8537 128877 -8503
rect 128887 -8537 128888 -8492
rect 128987 -8503 128988 -8492
rect 129232 -8496 129267 -8462
rect 129277 -8496 129278 -8451
rect 129377 -8462 129378 -8451
rect 129388 -8496 129423 -8462
rect 129433 -8496 129434 -8451
rect 129533 -8462 129534 -8451
rect 129714 -8456 129749 -8422
rect 129786 -8456 129821 -8422
rect 129858 -8456 129893 -8422
rect 130002 -8456 130037 -8422
rect 130074 -8456 130109 -8422
rect 130111 -8456 130181 -8422
rect 130218 -8456 130253 -8422
rect 130288 -8456 130323 -8422
rect 129544 -8496 129579 -8462
rect 130584 -8491 130619 -8457
rect 130629 -8491 130630 -8446
rect 130729 -8457 130730 -8446
rect 130740 -8491 130775 -8457
rect 130785 -8491 130786 -8446
rect 130885 -8457 130886 -8446
rect 131461 -8451 131496 -8417
rect 131638 -8451 131673 -8417
rect 130896 -8491 130931 -8457
rect 128998 -8537 129033 -8503
rect 130277 -8505 130278 -8494
rect 128644 -8577 128679 -8543
rect 127557 -8621 127592 -8587
rect 127758 -8666 127793 -8632
rect 127881 -8637 127882 -8595
rect 128203 -8624 128238 -8590
rect 128842 -8620 128877 -8586
rect 128887 -8620 128888 -8575
rect 128987 -8586 128988 -8575
rect 129232 -8580 129267 -8546
rect 129277 -8580 129278 -8535
rect 129377 -8546 129378 -8535
rect 129388 -8580 129423 -8546
rect 129433 -8580 129434 -8535
rect 129533 -8546 129534 -8535
rect 130111 -8539 130146 -8505
rect 130288 -8539 130323 -8505
rect 129544 -8580 129579 -8546
rect 130431 -8565 130546 -8499
rect 130729 -8525 130730 -8499
rect 131126 -8517 131161 -8483
rect 131171 -8517 131172 -8472
rect 131271 -8483 131272 -8472
rect 131282 -8517 131317 -8483
rect 131327 -8517 131328 -8472
rect 131627 -8500 131628 -8489
rect 131832 -8494 131867 -8460
rect 131877 -8494 131878 -8449
rect 131977 -8460 131978 -8449
rect 132186 -8453 132221 -8419
rect 132231 -8453 132232 -8408
rect 132331 -8419 132332 -8408
rect 132512 -8413 132547 -8379
rect 132576 -8413 132619 -8379
rect 132621 -8413 132622 -8371
rect 132721 -8379 132722 -8371
rect 132656 -8413 132691 -8379
rect 132732 -8413 132767 -8379
rect 132777 -8413 132778 -8371
rect 132877 -8379 132878 -8371
rect 132826 -8413 132861 -8379
rect 132888 -8413 132933 -8379
rect 133928 -8408 133963 -8374
rect 133973 -8408 133974 -8363
rect 134073 -8374 134074 -8363
rect 134084 -8408 134119 -8374
rect 134129 -8408 134130 -8363
rect 134229 -8374 134230 -8363
rect 134805 -8367 134840 -8333
rect 134982 -8367 135017 -8333
rect 135575 -8336 135576 -8328
rect 135675 -8336 135676 -8328
rect 134240 -8408 134275 -8374
rect 132342 -8453 132377 -8419
rect 133621 -8422 133622 -8414
rect 134971 -8417 134972 -8406
rect 135176 -8410 135211 -8376
rect 135221 -8410 135222 -8365
rect 135321 -8376 135322 -8365
rect 135502 -8370 135565 -8336
rect 135574 -8370 135609 -8336
rect 135686 -8370 135721 -8336
rect 136411 -8360 136446 -8326
rect 136507 -8360 136542 -8326
rect 136603 -8360 136638 -8326
rect 136699 -8360 136734 -8326
rect 136795 -8360 136830 -8326
rect 136891 -8360 136926 -8326
rect 136987 -8360 137022 -8326
rect 138315 -8333 138316 -8322
rect 138492 -8327 138555 -8293
rect 138564 -8327 138599 -8293
rect 138676 -8327 138711 -8293
rect 139207 -8317 139242 -8283
rect 139303 -8317 139338 -8283
rect 139399 -8317 139434 -8283
rect 139495 -8317 139530 -8283
rect 139591 -8317 139626 -8283
rect 140616 -8324 140651 -8290
rect 140661 -8324 140662 -8279
rect 140761 -8290 140762 -8279
rect 140772 -8324 140807 -8290
rect 140817 -8324 140818 -8279
rect 140917 -8290 140918 -8279
rect 141096 -8284 141131 -8250
rect 141168 -8284 141203 -8250
rect 141240 -8284 141275 -8250
rect 141384 -8284 141419 -8250
rect 141456 -8284 141491 -8250
rect 141493 -8284 141563 -8250
rect 141600 -8284 141635 -8250
rect 141670 -8284 141705 -8250
rect 142197 -8274 142232 -8240
rect 142293 -8274 142328 -8240
rect 142389 -8274 142424 -8240
rect 143896 -8241 143931 -8207
rect 143960 -8241 144003 -8207
rect 144005 -8241 144006 -8199
rect 144105 -8207 144106 -8199
rect 144040 -8241 144075 -8207
rect 144116 -8241 144151 -8207
rect 144161 -8241 144162 -8199
rect 144261 -8207 144262 -8199
rect 144210 -8241 144245 -8207
rect 144272 -8241 144317 -8207
rect 145187 -8231 145222 -8197
rect 145283 -8231 145318 -8197
rect 145379 -8231 145414 -8197
rect 145003 -8250 145004 -8242
rect 140928 -8324 140963 -8290
rect 141909 -8293 141910 -8285
rect 142009 -8293 142010 -8285
rect 135332 -8410 135367 -8376
rect 131988 -8494 132023 -8460
rect 128998 -8620 129033 -8586
rect 130277 -8589 130278 -8578
rect 127527 -8689 127528 -8681
rect 127538 -8723 127573 -8689
rect 127758 -8734 127793 -8700
rect 126205 -8793 126240 -8759
rect 126408 -8838 126443 -8804
rect 126531 -8809 126532 -8767
rect 126853 -8796 126888 -8762
rect 126175 -8861 126176 -8853
rect 126186 -8895 126221 -8861
rect 126408 -8906 126443 -8872
rect 126175 -8961 126176 -8950
rect 126186 -8995 126221 -8961
rect 125123 -9045 125158 -9011
rect 125219 -9045 125254 -9011
rect 125315 -9045 125350 -9011
rect 125824 -9035 125859 -9001
rect 125896 -9035 125931 -9001
rect 125968 -9035 126003 -9001
rect 126040 -9029 126076 -9001
rect 126386 -9025 126421 -8991
rect 126431 -9025 126432 -8980
rect 126040 -9035 126075 -9029
rect 125477 -9088 125512 -9054
rect 125573 -9088 125608 -9054
rect 125669 -9088 125704 -9054
rect 126573 -9076 126574 -8809
rect 127202 -8819 127589 -8753
rect 126589 -8860 126624 -8826
rect 126938 -8832 126949 -8819
rect 126872 -8874 126949 -8832
rect 127000 -8874 127589 -8819
rect 127736 -8853 127771 -8819
rect 127781 -8853 127782 -8808
rect 126872 -8877 127589 -8874
rect 126589 -8928 126624 -8894
rect 126792 -8942 126827 -8908
rect 126837 -8942 126838 -8900
rect 126673 -8991 126674 -8980
rect 126684 -9025 126719 -8991
rect 126792 -9042 126827 -9008
rect 126837 -9042 126838 -8997
rect 126685 -9078 126720 -9044
rect 126757 -9078 126792 -9044
rect 126829 -9078 126864 -9044
rect 125831 -9131 125866 -9097
rect 125927 -9131 125962 -9097
rect 126023 -9131 126058 -9097
rect 126119 -9131 126154 -9097
rect 126215 -9131 126250 -9097
rect 126872 -9114 127017 -8877
rect 127202 -8899 127589 -8877
rect 127126 -8925 127589 -8899
rect 127923 -8904 127924 -8637
rect 127939 -8688 127974 -8654
rect 128553 -8691 128588 -8657
rect 129232 -8663 129267 -8629
rect 129277 -8663 129278 -8618
rect 129377 -8629 129378 -8618
rect 129388 -8663 129423 -8629
rect 129433 -8663 129434 -8618
rect 129533 -8629 129534 -8618
rect 130111 -8623 130146 -8589
rect 130288 -8623 130323 -8589
rect 130649 -8605 130684 -8571
rect 129544 -8663 129579 -8629
rect 129377 -8697 129378 -8671
rect 129776 -8689 129811 -8655
rect 129821 -8689 129822 -8644
rect 129921 -8655 129922 -8644
rect 129932 -8689 129967 -8655
rect 129977 -8689 129978 -8644
rect 130277 -8672 130278 -8661
rect 127939 -8756 127974 -8722
rect 128142 -8770 128177 -8736
rect 128187 -8770 128188 -8728
rect 128287 -8740 128288 -8729
rect 128907 -8734 128942 -8700
rect 128298 -8774 128333 -8740
rect 128023 -8819 128024 -8808
rect 128492 -8813 128527 -8779
rect 128537 -8813 128538 -8771
rect 128637 -8779 128638 -8771
rect 129297 -8777 129332 -8743
rect 128648 -8813 128683 -8779
rect 128034 -8853 128069 -8819
rect 128142 -8870 128177 -8836
rect 128187 -8870 128188 -8825
rect 128287 -8832 128288 -8821
rect 128298 -8866 128333 -8832
rect 128846 -8856 128881 -8822
rect 128891 -8856 128892 -8814
rect 128991 -8822 128992 -8814
rect 129002 -8856 129037 -8822
rect 128035 -8906 128070 -8872
rect 128107 -8906 128142 -8872
rect 128179 -8906 128214 -8872
rect 128492 -8913 128527 -8879
rect 128537 -8913 128538 -8868
rect 128637 -8879 128638 -8868
rect 128648 -8913 128683 -8879
rect 129232 -8895 129267 -8861
rect 129277 -8895 129278 -8853
rect 127126 -8959 127602 -8925
rect 128460 -8949 128495 -8915
rect 128532 -8949 128567 -8915
rect 128846 -8956 128881 -8922
rect 128891 -8956 128892 -8911
rect 128991 -8922 128992 -8911
rect 129002 -8956 129037 -8922
rect 127126 -8985 127589 -8959
rect 127130 -8993 127331 -8985
rect 127146 -9003 127315 -8993
rect 126872 -9140 127047 -9114
rect 126379 -9174 126414 -9140
rect 126475 -9174 126510 -9140
rect 126571 -9174 126606 -9140
rect 126667 -9174 126702 -9140
rect 126763 -9174 126798 -9140
rect 126859 -9174 127047 -9140
rect 126872 -9200 127047 -9174
rect 127072 -9174 127173 -9050
rect 126950 -9870 126985 -9200
rect 127072 -9228 127075 -9174
rect 126757 -9936 126902 -9924
rect 126425 -9970 126902 -9936
rect 126757 -9971 126902 -9970
rect 126938 -9971 126985 -9870
rect 127084 -9971 127119 -9174
rect 127342 -9971 127377 -9062
rect 127476 -9971 127511 -8985
rect 127729 -9002 127764 -8968
rect 127825 -9002 127860 -8968
rect 127921 -9002 127956 -8968
rect 128017 -9002 128052 -8968
rect 128113 -9002 128148 -8968
rect 128209 -9002 128244 -8968
rect 128305 -9002 128340 -8968
rect 128814 -8992 128849 -8958
rect 128886 -8992 128921 -8958
rect 129232 -8995 129267 -8961
rect 129277 -8995 129278 -8950
rect 129419 -9001 129420 -8697
rect 130111 -8706 130146 -8672
rect 130288 -8706 130323 -8672
rect 130584 -8723 130619 -8689
rect 130629 -8723 130630 -8681
rect 130771 -8753 130772 -8525
rect 131461 -8534 131496 -8500
rect 131638 -8534 131673 -8500
rect 131832 -8577 131867 -8543
rect 131877 -8577 131878 -8532
rect 131977 -8543 131978 -8532
rect 132186 -8537 132221 -8503
rect 132231 -8537 132232 -8492
rect 132331 -8503 132332 -8492
rect 132576 -8496 132611 -8462
rect 132621 -8496 132622 -8451
rect 132721 -8462 132722 -8451
rect 132732 -8496 132767 -8462
rect 132777 -8496 132778 -8451
rect 132877 -8462 132878 -8451
rect 133058 -8456 133093 -8422
rect 133130 -8456 133165 -8422
rect 133202 -8456 133237 -8422
rect 133346 -8456 133381 -8422
rect 133418 -8456 133453 -8422
rect 133455 -8456 133525 -8422
rect 133562 -8456 133597 -8422
rect 133632 -8456 133667 -8422
rect 132888 -8496 132923 -8462
rect 133928 -8491 133963 -8457
rect 133973 -8491 133974 -8446
rect 134073 -8457 134074 -8446
rect 134084 -8491 134119 -8457
rect 134129 -8491 134130 -8446
rect 134229 -8457 134230 -8446
rect 134805 -8451 134840 -8417
rect 134982 -8451 135017 -8417
rect 134240 -8491 134275 -8457
rect 132342 -8537 132377 -8503
rect 133621 -8505 133622 -8494
rect 131988 -8577 132023 -8543
rect 130901 -8621 130936 -8587
rect 131102 -8666 131137 -8632
rect 131225 -8637 131226 -8595
rect 131547 -8624 131582 -8590
rect 132186 -8620 132221 -8586
rect 132231 -8620 132232 -8575
rect 132331 -8586 132332 -8575
rect 132576 -8580 132611 -8546
rect 132621 -8580 132622 -8535
rect 132721 -8546 132722 -8535
rect 132732 -8580 132767 -8546
rect 132777 -8580 132778 -8535
rect 132877 -8546 132878 -8535
rect 133455 -8539 133490 -8505
rect 133632 -8539 133667 -8505
rect 132888 -8580 132923 -8546
rect 133775 -8565 133890 -8499
rect 134073 -8525 134074 -8499
rect 134470 -8517 134505 -8483
rect 134515 -8517 134516 -8472
rect 134615 -8483 134616 -8472
rect 134626 -8517 134661 -8483
rect 134671 -8517 134672 -8472
rect 134971 -8500 134972 -8489
rect 135176 -8494 135211 -8460
rect 135221 -8494 135222 -8449
rect 135321 -8460 135322 -8449
rect 135530 -8453 135565 -8419
rect 135575 -8453 135576 -8408
rect 135675 -8419 135676 -8408
rect 135856 -8413 135891 -8379
rect 135920 -8413 135963 -8379
rect 135965 -8413 135966 -8371
rect 136065 -8379 136066 -8371
rect 136000 -8413 136035 -8379
rect 136076 -8413 136111 -8379
rect 136121 -8413 136122 -8371
rect 136221 -8379 136222 -8371
rect 136170 -8413 136205 -8379
rect 136232 -8413 136277 -8379
rect 137272 -8408 137307 -8374
rect 137317 -8408 137318 -8363
rect 137417 -8374 137418 -8363
rect 137428 -8408 137463 -8374
rect 137473 -8408 137474 -8363
rect 137573 -8374 137574 -8363
rect 138149 -8367 138184 -8333
rect 138326 -8367 138361 -8333
rect 138919 -8336 138920 -8328
rect 139019 -8336 139020 -8328
rect 137584 -8408 137619 -8374
rect 135686 -8453 135721 -8419
rect 136965 -8422 136966 -8414
rect 138315 -8417 138316 -8406
rect 138520 -8410 138555 -8376
rect 138565 -8410 138566 -8365
rect 138665 -8376 138666 -8365
rect 138846 -8370 138909 -8336
rect 138918 -8370 138953 -8336
rect 139030 -8370 139065 -8336
rect 139755 -8360 139790 -8326
rect 139851 -8360 139886 -8326
rect 139947 -8360 139982 -8326
rect 140043 -8360 140078 -8326
rect 140139 -8360 140174 -8326
rect 140235 -8360 140270 -8326
rect 140331 -8360 140366 -8326
rect 141659 -8333 141660 -8322
rect 141836 -8327 141899 -8293
rect 141908 -8327 141943 -8293
rect 142020 -8327 142055 -8293
rect 142551 -8317 142586 -8283
rect 142647 -8317 142682 -8283
rect 142743 -8317 142778 -8283
rect 142839 -8317 142874 -8283
rect 142935 -8317 142970 -8283
rect 143960 -8324 143995 -8290
rect 144005 -8324 144006 -8279
rect 144105 -8290 144106 -8279
rect 144116 -8324 144151 -8290
rect 144161 -8324 144162 -8279
rect 144261 -8290 144262 -8279
rect 144440 -8284 144475 -8250
rect 144512 -8284 144547 -8250
rect 144584 -8284 144619 -8250
rect 144728 -8284 144763 -8250
rect 144800 -8284 144835 -8250
rect 144837 -8284 144907 -8250
rect 144944 -8284 144979 -8250
rect 145014 -8284 145049 -8250
rect 145541 -8274 145576 -8240
rect 145637 -8274 145672 -8240
rect 145733 -8274 145768 -8240
rect 147240 -8241 147275 -8207
rect 147304 -8241 147347 -8207
rect 147349 -8241 147350 -8199
rect 147449 -8207 147450 -8199
rect 147384 -8241 147419 -8207
rect 147460 -8241 147495 -8207
rect 147505 -8241 147506 -8199
rect 147605 -8207 147606 -8199
rect 147554 -8241 147589 -8207
rect 147616 -8241 147661 -8207
rect 148531 -8231 148566 -8197
rect 148627 -8231 148662 -8197
rect 148723 -8231 148758 -8197
rect 148347 -8250 148348 -8242
rect 144272 -8324 144307 -8290
rect 145253 -8293 145254 -8285
rect 145353 -8293 145354 -8285
rect 138676 -8410 138711 -8376
rect 135332 -8494 135367 -8460
rect 132342 -8620 132377 -8586
rect 133621 -8589 133622 -8578
rect 130871 -8689 130872 -8681
rect 130882 -8723 130917 -8689
rect 131102 -8734 131137 -8700
rect 129549 -8793 129584 -8759
rect 129752 -8838 129787 -8804
rect 129875 -8809 129876 -8767
rect 130197 -8796 130232 -8762
rect 129519 -8861 129520 -8853
rect 129530 -8895 129565 -8861
rect 129752 -8906 129787 -8872
rect 129519 -8961 129520 -8950
rect 129530 -8995 129565 -8961
rect 128467 -9045 128502 -9011
rect 128563 -9045 128598 -9011
rect 128659 -9045 128694 -9011
rect 129168 -9035 129203 -9001
rect 129240 -9035 129275 -9001
rect 129312 -9035 129347 -9001
rect 129384 -9029 129420 -9001
rect 129730 -9025 129765 -8991
rect 129775 -9025 129776 -8980
rect 129384 -9035 129419 -9029
rect 128821 -9088 128856 -9054
rect 128917 -9088 128952 -9054
rect 129013 -9088 129048 -9054
rect 129917 -9076 129918 -8809
rect 130546 -8819 130933 -8753
rect 129933 -8860 129968 -8826
rect 130282 -8832 130293 -8819
rect 130216 -8874 130293 -8832
rect 130344 -8874 130933 -8819
rect 131080 -8853 131115 -8819
rect 131125 -8853 131126 -8808
rect 130216 -8877 130933 -8874
rect 129933 -8928 129968 -8894
rect 130136 -8942 130171 -8908
rect 130181 -8942 130182 -8900
rect 130017 -8991 130018 -8980
rect 130028 -9025 130063 -8991
rect 130136 -9042 130171 -9008
rect 130181 -9042 130182 -8997
rect 130029 -9078 130064 -9044
rect 130101 -9078 130136 -9044
rect 130173 -9078 130208 -9044
rect 129175 -9131 129210 -9097
rect 129271 -9131 129306 -9097
rect 129367 -9131 129402 -9097
rect 129463 -9131 129498 -9097
rect 129559 -9131 129594 -9097
rect 130216 -9114 130361 -8877
rect 130546 -8899 130933 -8877
rect 130470 -8925 130933 -8899
rect 131267 -8904 131268 -8637
rect 131283 -8688 131318 -8654
rect 131897 -8691 131932 -8657
rect 132576 -8663 132611 -8629
rect 132621 -8663 132622 -8618
rect 132721 -8629 132722 -8618
rect 132732 -8663 132767 -8629
rect 132777 -8663 132778 -8618
rect 132877 -8629 132878 -8618
rect 133455 -8623 133490 -8589
rect 133632 -8623 133667 -8589
rect 133993 -8605 134028 -8571
rect 132888 -8663 132923 -8629
rect 132721 -8697 132722 -8671
rect 133120 -8689 133155 -8655
rect 133165 -8689 133166 -8644
rect 133265 -8655 133266 -8644
rect 133276 -8689 133311 -8655
rect 133321 -8689 133322 -8644
rect 133621 -8672 133622 -8661
rect 131283 -8756 131318 -8722
rect 131486 -8770 131521 -8736
rect 131531 -8770 131532 -8728
rect 131631 -8740 131632 -8729
rect 132251 -8734 132286 -8700
rect 131642 -8774 131677 -8740
rect 131367 -8819 131368 -8808
rect 131836 -8813 131871 -8779
rect 131881 -8813 131882 -8771
rect 131981 -8779 131982 -8771
rect 132641 -8777 132676 -8743
rect 131992 -8813 132027 -8779
rect 131378 -8853 131413 -8819
rect 131486 -8870 131521 -8836
rect 131531 -8870 131532 -8825
rect 131631 -8832 131632 -8821
rect 131642 -8866 131677 -8832
rect 132190 -8856 132225 -8822
rect 132235 -8856 132236 -8814
rect 132335 -8822 132336 -8814
rect 132346 -8856 132381 -8822
rect 131379 -8906 131414 -8872
rect 131451 -8906 131486 -8872
rect 131523 -8906 131558 -8872
rect 131836 -8913 131871 -8879
rect 131881 -8913 131882 -8868
rect 131981 -8879 131982 -8868
rect 131992 -8913 132027 -8879
rect 132576 -8895 132611 -8861
rect 132621 -8895 132622 -8853
rect 130470 -8959 130946 -8925
rect 131804 -8949 131839 -8915
rect 131876 -8949 131911 -8915
rect 132190 -8956 132225 -8922
rect 132235 -8956 132236 -8911
rect 132335 -8922 132336 -8911
rect 132346 -8956 132381 -8922
rect 130470 -8985 130933 -8959
rect 130474 -8993 130675 -8985
rect 130490 -9003 130659 -8993
rect 130216 -9140 130391 -9114
rect 129723 -9174 129758 -9140
rect 129819 -9174 129854 -9140
rect 129915 -9174 129950 -9140
rect 130011 -9174 130046 -9140
rect 130107 -9174 130142 -9140
rect 130203 -9174 130391 -9140
rect 130216 -9200 130391 -9174
rect 130416 -9174 130517 -9050
rect 130294 -9870 130329 -9200
rect 130416 -9228 130419 -9174
rect 130101 -9936 130246 -9924
rect 129769 -9970 130246 -9936
rect 130101 -9971 130246 -9970
rect 130282 -9971 130329 -9870
rect 130428 -9971 130463 -9174
rect 130686 -9971 130721 -9062
rect 130820 -9971 130855 -8985
rect 131073 -9002 131108 -8968
rect 131169 -9002 131204 -8968
rect 131265 -9002 131300 -8968
rect 131361 -9002 131396 -8968
rect 131457 -9002 131492 -8968
rect 131553 -9002 131588 -8968
rect 131649 -9002 131684 -8968
rect 132158 -8992 132193 -8958
rect 132230 -8992 132265 -8958
rect 132576 -8995 132611 -8961
rect 132621 -8995 132622 -8950
rect 132763 -9001 132764 -8697
rect 133455 -8706 133490 -8672
rect 133632 -8706 133667 -8672
rect 133928 -8723 133963 -8689
rect 133973 -8723 133974 -8681
rect 134115 -8753 134116 -8525
rect 134805 -8534 134840 -8500
rect 134982 -8534 135017 -8500
rect 135176 -8577 135211 -8543
rect 135221 -8577 135222 -8532
rect 135321 -8543 135322 -8532
rect 135530 -8537 135565 -8503
rect 135575 -8537 135576 -8492
rect 135675 -8503 135676 -8492
rect 135920 -8496 135955 -8462
rect 135965 -8496 135966 -8451
rect 136065 -8462 136066 -8451
rect 136076 -8496 136111 -8462
rect 136121 -8496 136122 -8451
rect 136221 -8462 136222 -8451
rect 136402 -8456 136437 -8422
rect 136474 -8456 136509 -8422
rect 136546 -8456 136581 -8422
rect 136690 -8456 136725 -8422
rect 136762 -8456 136797 -8422
rect 136799 -8456 136869 -8422
rect 136906 -8456 136941 -8422
rect 136976 -8456 137011 -8422
rect 136232 -8496 136267 -8462
rect 137272 -8491 137307 -8457
rect 137317 -8491 137318 -8446
rect 137417 -8457 137418 -8446
rect 137428 -8491 137463 -8457
rect 137473 -8491 137474 -8446
rect 137573 -8457 137574 -8446
rect 138149 -8451 138184 -8417
rect 138326 -8451 138361 -8417
rect 137584 -8491 137619 -8457
rect 135686 -8537 135721 -8503
rect 136965 -8505 136966 -8494
rect 135332 -8577 135367 -8543
rect 134245 -8621 134280 -8587
rect 134446 -8666 134481 -8632
rect 134569 -8637 134570 -8595
rect 134891 -8624 134926 -8590
rect 135530 -8620 135565 -8586
rect 135575 -8620 135576 -8575
rect 135675 -8586 135676 -8575
rect 135920 -8580 135955 -8546
rect 135965 -8580 135966 -8535
rect 136065 -8546 136066 -8535
rect 136076 -8580 136111 -8546
rect 136121 -8580 136122 -8535
rect 136221 -8546 136222 -8535
rect 136799 -8539 136834 -8505
rect 136976 -8539 137011 -8505
rect 136232 -8580 136267 -8546
rect 137119 -8565 137234 -8499
rect 137417 -8525 137418 -8499
rect 137814 -8517 137849 -8483
rect 137859 -8517 137860 -8472
rect 137959 -8483 137960 -8472
rect 137970 -8517 138005 -8483
rect 138015 -8517 138016 -8472
rect 138315 -8500 138316 -8489
rect 138520 -8494 138555 -8460
rect 138565 -8494 138566 -8449
rect 138665 -8460 138666 -8449
rect 138874 -8453 138909 -8419
rect 138919 -8453 138920 -8408
rect 139019 -8419 139020 -8408
rect 139200 -8413 139235 -8379
rect 139264 -8413 139307 -8379
rect 139309 -8413 139310 -8371
rect 139409 -8379 139410 -8371
rect 139344 -8413 139379 -8379
rect 139420 -8413 139455 -8379
rect 139465 -8413 139466 -8371
rect 139565 -8379 139566 -8371
rect 139514 -8413 139549 -8379
rect 139576 -8413 139621 -8379
rect 140616 -8408 140651 -8374
rect 140661 -8408 140662 -8363
rect 140761 -8374 140762 -8363
rect 140772 -8408 140807 -8374
rect 140817 -8408 140818 -8363
rect 140917 -8374 140918 -8363
rect 141493 -8367 141528 -8333
rect 141670 -8367 141705 -8333
rect 142263 -8336 142264 -8328
rect 142363 -8336 142364 -8328
rect 140928 -8408 140963 -8374
rect 139030 -8453 139065 -8419
rect 140309 -8422 140310 -8414
rect 141659 -8417 141660 -8406
rect 141864 -8410 141899 -8376
rect 141909 -8410 141910 -8365
rect 142009 -8376 142010 -8365
rect 142190 -8370 142253 -8336
rect 142262 -8370 142297 -8336
rect 142374 -8370 142409 -8336
rect 143099 -8360 143134 -8326
rect 143195 -8360 143230 -8326
rect 143291 -8360 143326 -8326
rect 143387 -8360 143422 -8326
rect 143483 -8360 143518 -8326
rect 143579 -8360 143614 -8326
rect 143675 -8360 143710 -8326
rect 145003 -8333 145004 -8322
rect 145180 -8327 145243 -8293
rect 145252 -8327 145287 -8293
rect 145364 -8327 145399 -8293
rect 145895 -8317 145930 -8283
rect 145991 -8317 146026 -8283
rect 146087 -8317 146122 -8283
rect 146183 -8317 146218 -8283
rect 146279 -8317 146314 -8283
rect 147304 -8324 147339 -8290
rect 147349 -8324 147350 -8279
rect 147449 -8290 147450 -8279
rect 147460 -8324 147495 -8290
rect 147505 -8324 147506 -8279
rect 147605 -8290 147606 -8279
rect 147784 -8284 147819 -8250
rect 147856 -8284 147891 -8250
rect 147928 -8284 147963 -8250
rect 148072 -8284 148107 -8250
rect 148144 -8284 148179 -8250
rect 148181 -8284 148251 -8250
rect 148288 -8284 148323 -8250
rect 148358 -8284 148393 -8250
rect 148885 -8274 148920 -8240
rect 148981 -8274 149016 -8240
rect 149077 -8274 149112 -8240
rect 150584 -8241 150619 -8207
rect 150648 -8241 150691 -8207
rect 150693 -8241 150694 -8199
rect 150793 -8207 150794 -8199
rect 150728 -8241 150763 -8207
rect 150804 -8241 150839 -8207
rect 150849 -8241 150850 -8199
rect 150949 -8207 150950 -8199
rect 150898 -8241 150933 -8207
rect 150960 -8241 151005 -8207
rect 151875 -8231 151910 -8197
rect 151971 -8231 152006 -8197
rect 152067 -8231 152102 -8197
rect 151691 -8250 151692 -8242
rect 147616 -8324 147651 -8290
rect 148597 -8293 148598 -8285
rect 148697 -8293 148698 -8285
rect 142020 -8410 142055 -8376
rect 138676 -8494 138711 -8460
rect 135686 -8620 135721 -8586
rect 136965 -8589 136966 -8578
rect 134215 -8689 134216 -8681
rect 134226 -8723 134261 -8689
rect 134446 -8734 134481 -8700
rect 132893 -8793 132928 -8759
rect 133096 -8838 133131 -8804
rect 133219 -8809 133220 -8767
rect 133541 -8796 133576 -8762
rect 132863 -8861 132864 -8853
rect 132874 -8895 132909 -8861
rect 133096 -8906 133131 -8872
rect 132863 -8961 132864 -8950
rect 132874 -8995 132909 -8961
rect 131811 -9045 131846 -9011
rect 131907 -9045 131942 -9011
rect 132003 -9045 132038 -9011
rect 132512 -9035 132547 -9001
rect 132584 -9035 132619 -9001
rect 132656 -9035 132691 -9001
rect 132728 -9029 132764 -9001
rect 133074 -9025 133109 -8991
rect 133119 -9025 133120 -8980
rect 132728 -9035 132763 -9029
rect 132165 -9088 132200 -9054
rect 132261 -9088 132296 -9054
rect 132357 -9088 132392 -9054
rect 133261 -9076 133262 -8809
rect 133890 -8819 134277 -8753
rect 133277 -8860 133312 -8826
rect 133626 -8832 133637 -8819
rect 133560 -8874 133637 -8832
rect 133688 -8874 134277 -8819
rect 134424 -8853 134459 -8819
rect 134469 -8853 134470 -8808
rect 133560 -8877 134277 -8874
rect 133277 -8928 133312 -8894
rect 133480 -8942 133515 -8908
rect 133525 -8942 133526 -8900
rect 133361 -8991 133362 -8980
rect 133372 -9025 133407 -8991
rect 133480 -9042 133515 -9008
rect 133525 -9042 133526 -8997
rect 133373 -9078 133408 -9044
rect 133445 -9078 133480 -9044
rect 133517 -9078 133552 -9044
rect 132519 -9131 132554 -9097
rect 132615 -9131 132650 -9097
rect 132711 -9131 132746 -9097
rect 132807 -9131 132842 -9097
rect 132903 -9131 132938 -9097
rect 133560 -9114 133705 -8877
rect 133890 -8899 134277 -8877
rect 133814 -8925 134277 -8899
rect 134611 -8904 134612 -8637
rect 134627 -8688 134662 -8654
rect 135241 -8691 135276 -8657
rect 135920 -8663 135955 -8629
rect 135965 -8663 135966 -8618
rect 136065 -8629 136066 -8618
rect 136076 -8663 136111 -8629
rect 136121 -8663 136122 -8618
rect 136221 -8629 136222 -8618
rect 136799 -8623 136834 -8589
rect 136976 -8623 137011 -8589
rect 137337 -8605 137372 -8571
rect 136232 -8663 136267 -8629
rect 136065 -8697 136066 -8671
rect 136464 -8689 136499 -8655
rect 136509 -8689 136510 -8644
rect 136609 -8655 136610 -8644
rect 136620 -8689 136655 -8655
rect 136665 -8689 136666 -8644
rect 136965 -8672 136966 -8661
rect 134627 -8756 134662 -8722
rect 134830 -8770 134865 -8736
rect 134875 -8770 134876 -8728
rect 134975 -8740 134976 -8729
rect 135595 -8734 135630 -8700
rect 134986 -8774 135021 -8740
rect 134711 -8819 134712 -8808
rect 135180 -8813 135215 -8779
rect 135225 -8813 135226 -8771
rect 135325 -8779 135326 -8771
rect 135985 -8777 136020 -8743
rect 135336 -8813 135371 -8779
rect 134722 -8853 134757 -8819
rect 134830 -8870 134865 -8836
rect 134875 -8870 134876 -8825
rect 134975 -8832 134976 -8821
rect 134986 -8866 135021 -8832
rect 135534 -8856 135569 -8822
rect 135579 -8856 135580 -8814
rect 135679 -8822 135680 -8814
rect 135690 -8856 135725 -8822
rect 134723 -8906 134758 -8872
rect 134795 -8906 134830 -8872
rect 134867 -8906 134902 -8872
rect 135180 -8913 135215 -8879
rect 135225 -8913 135226 -8868
rect 135325 -8879 135326 -8868
rect 135336 -8913 135371 -8879
rect 135920 -8895 135955 -8861
rect 135965 -8895 135966 -8853
rect 133814 -8959 134290 -8925
rect 135148 -8949 135183 -8915
rect 135220 -8949 135255 -8915
rect 135534 -8956 135569 -8922
rect 135579 -8956 135580 -8911
rect 135679 -8922 135680 -8911
rect 135690 -8956 135725 -8922
rect 133814 -8985 134277 -8959
rect 133818 -8993 134019 -8985
rect 133834 -9003 134003 -8993
rect 133560 -9140 133735 -9114
rect 133067 -9174 133102 -9140
rect 133163 -9174 133198 -9140
rect 133259 -9174 133294 -9140
rect 133355 -9174 133390 -9140
rect 133451 -9174 133486 -9140
rect 133547 -9174 133735 -9140
rect 133560 -9200 133735 -9174
rect 133760 -9174 133861 -9050
rect 133638 -9870 133673 -9200
rect 133760 -9228 133763 -9174
rect 133445 -9936 133590 -9924
rect 133113 -9970 133590 -9936
rect 133445 -9971 133590 -9970
rect 133626 -9971 133673 -9870
rect 133772 -9971 133807 -9174
rect 134030 -9971 134065 -9062
rect 134164 -9971 134199 -8985
rect 134417 -9002 134452 -8968
rect 134513 -9002 134548 -8968
rect 134609 -9002 134644 -8968
rect 134705 -9002 134740 -8968
rect 134801 -9002 134836 -8968
rect 134897 -9002 134932 -8968
rect 134993 -9002 135028 -8968
rect 135502 -8992 135537 -8958
rect 135574 -8992 135609 -8958
rect 135920 -8995 135955 -8961
rect 135965 -8995 135966 -8950
rect 136107 -9001 136108 -8697
rect 136799 -8706 136834 -8672
rect 136976 -8706 137011 -8672
rect 137272 -8723 137307 -8689
rect 137317 -8723 137318 -8681
rect 137459 -8753 137460 -8525
rect 138149 -8534 138184 -8500
rect 138326 -8534 138361 -8500
rect 138520 -8577 138555 -8543
rect 138565 -8577 138566 -8532
rect 138665 -8543 138666 -8532
rect 138874 -8537 138909 -8503
rect 138919 -8537 138920 -8492
rect 139019 -8503 139020 -8492
rect 139264 -8496 139299 -8462
rect 139309 -8496 139310 -8451
rect 139409 -8462 139410 -8451
rect 139420 -8496 139455 -8462
rect 139465 -8496 139466 -8451
rect 139565 -8462 139566 -8451
rect 139746 -8456 139781 -8422
rect 139818 -8456 139853 -8422
rect 139890 -8456 139925 -8422
rect 140034 -8456 140069 -8422
rect 140106 -8456 140141 -8422
rect 140143 -8456 140213 -8422
rect 140250 -8456 140285 -8422
rect 140320 -8456 140355 -8422
rect 139576 -8496 139611 -8462
rect 140616 -8491 140651 -8457
rect 140661 -8491 140662 -8446
rect 140761 -8457 140762 -8446
rect 140772 -8491 140807 -8457
rect 140817 -8491 140818 -8446
rect 140917 -8457 140918 -8446
rect 141493 -8451 141528 -8417
rect 141670 -8451 141705 -8417
rect 140928 -8491 140963 -8457
rect 139030 -8537 139065 -8503
rect 140309 -8505 140310 -8494
rect 138676 -8577 138711 -8543
rect 137589 -8621 137624 -8587
rect 137790 -8666 137825 -8632
rect 137913 -8637 137914 -8595
rect 138235 -8624 138270 -8590
rect 138874 -8620 138909 -8586
rect 138919 -8620 138920 -8575
rect 139019 -8586 139020 -8575
rect 139264 -8580 139299 -8546
rect 139309 -8580 139310 -8535
rect 139409 -8546 139410 -8535
rect 139420 -8580 139455 -8546
rect 139465 -8580 139466 -8535
rect 139565 -8546 139566 -8535
rect 140143 -8539 140178 -8505
rect 140320 -8539 140355 -8505
rect 139576 -8580 139611 -8546
rect 140463 -8565 140578 -8499
rect 140761 -8525 140762 -8499
rect 141158 -8517 141193 -8483
rect 141203 -8517 141204 -8472
rect 141303 -8483 141304 -8472
rect 141314 -8517 141349 -8483
rect 141359 -8517 141360 -8472
rect 141659 -8500 141660 -8489
rect 141864 -8494 141899 -8460
rect 141909 -8494 141910 -8449
rect 142009 -8460 142010 -8449
rect 142218 -8453 142253 -8419
rect 142263 -8453 142264 -8408
rect 142363 -8419 142364 -8408
rect 142544 -8413 142579 -8379
rect 142608 -8413 142651 -8379
rect 142653 -8413 142654 -8371
rect 142753 -8379 142754 -8371
rect 142688 -8413 142723 -8379
rect 142764 -8413 142799 -8379
rect 142809 -8413 142810 -8371
rect 142909 -8379 142910 -8371
rect 142858 -8413 142893 -8379
rect 142920 -8413 142965 -8379
rect 143960 -8408 143995 -8374
rect 144005 -8408 144006 -8363
rect 144105 -8374 144106 -8363
rect 144116 -8408 144151 -8374
rect 144161 -8408 144162 -8363
rect 144261 -8374 144262 -8363
rect 144837 -8367 144872 -8333
rect 145014 -8367 145049 -8333
rect 145607 -8336 145608 -8328
rect 145707 -8336 145708 -8328
rect 144272 -8408 144307 -8374
rect 142374 -8453 142409 -8419
rect 143653 -8422 143654 -8414
rect 145003 -8417 145004 -8406
rect 145208 -8410 145243 -8376
rect 145253 -8410 145254 -8365
rect 145353 -8376 145354 -8365
rect 145534 -8370 145597 -8336
rect 145606 -8370 145641 -8336
rect 145718 -8370 145753 -8336
rect 146443 -8360 146478 -8326
rect 146539 -8360 146574 -8326
rect 146635 -8360 146670 -8326
rect 146731 -8360 146766 -8326
rect 146827 -8360 146862 -8326
rect 146923 -8360 146958 -8326
rect 147019 -8360 147054 -8326
rect 148347 -8333 148348 -8322
rect 148524 -8327 148587 -8293
rect 148596 -8327 148631 -8293
rect 148708 -8327 148743 -8293
rect 149239 -8317 149274 -8283
rect 149335 -8317 149370 -8283
rect 149431 -8317 149466 -8283
rect 149527 -8317 149562 -8283
rect 149623 -8317 149658 -8283
rect 150648 -8324 150683 -8290
rect 150693 -8324 150694 -8279
rect 150793 -8290 150794 -8279
rect 150804 -8324 150839 -8290
rect 150849 -8324 150850 -8279
rect 150949 -8290 150950 -8279
rect 151128 -8284 151163 -8250
rect 151200 -8284 151235 -8250
rect 151272 -8284 151307 -8250
rect 151416 -8284 151451 -8250
rect 151488 -8284 151523 -8250
rect 151525 -8284 151595 -8250
rect 151632 -8284 151667 -8250
rect 151702 -8284 151737 -8250
rect 152229 -8274 152264 -8240
rect 152325 -8274 152360 -8240
rect 152421 -8274 152456 -8240
rect 153928 -8241 153963 -8207
rect 153992 -8241 154035 -8207
rect 154037 -8241 154038 -8199
rect 154137 -8207 154138 -8199
rect 154072 -8241 154107 -8207
rect 154148 -8241 154183 -8207
rect 154193 -8241 154194 -8199
rect 154293 -8207 154294 -8199
rect 154242 -8241 154277 -8207
rect 154304 -8241 154349 -8207
rect 155219 -8231 155254 -8197
rect 155315 -8231 155350 -8197
rect 155411 -8231 155446 -8197
rect 155035 -8250 155036 -8242
rect 150960 -8324 150995 -8290
rect 151941 -8293 151942 -8285
rect 152041 -8293 152042 -8285
rect 145364 -8410 145399 -8376
rect 142020 -8494 142055 -8460
rect 139030 -8620 139065 -8586
rect 140309 -8589 140310 -8578
rect 137559 -8689 137560 -8681
rect 137570 -8723 137605 -8689
rect 137790 -8734 137825 -8700
rect 136237 -8793 136272 -8759
rect 136440 -8838 136475 -8804
rect 136563 -8809 136564 -8767
rect 136885 -8796 136920 -8762
rect 136207 -8861 136208 -8853
rect 136218 -8895 136253 -8861
rect 136440 -8906 136475 -8872
rect 136207 -8961 136208 -8950
rect 136218 -8995 136253 -8961
rect 135155 -9045 135190 -9011
rect 135251 -9045 135286 -9011
rect 135347 -9045 135382 -9011
rect 135856 -9035 135891 -9001
rect 135928 -9035 135963 -9001
rect 136000 -9035 136035 -9001
rect 136072 -9029 136108 -9001
rect 136418 -9025 136453 -8991
rect 136463 -9025 136464 -8980
rect 136072 -9035 136107 -9029
rect 135509 -9088 135544 -9054
rect 135605 -9088 135640 -9054
rect 135701 -9088 135736 -9054
rect 136605 -9076 136606 -8809
rect 137234 -8819 137621 -8753
rect 136621 -8860 136656 -8826
rect 136970 -8832 136981 -8819
rect 136904 -8874 136981 -8832
rect 137032 -8874 137621 -8819
rect 137768 -8853 137803 -8819
rect 137813 -8853 137814 -8808
rect 136904 -8877 137621 -8874
rect 136621 -8928 136656 -8894
rect 136824 -8942 136859 -8908
rect 136869 -8942 136870 -8900
rect 136705 -8991 136706 -8980
rect 136716 -9025 136751 -8991
rect 136824 -9042 136859 -9008
rect 136869 -9042 136870 -8997
rect 136717 -9078 136752 -9044
rect 136789 -9078 136824 -9044
rect 136861 -9078 136896 -9044
rect 135863 -9131 135898 -9097
rect 135959 -9131 135994 -9097
rect 136055 -9131 136090 -9097
rect 136151 -9131 136186 -9097
rect 136247 -9131 136282 -9097
rect 136904 -9114 137049 -8877
rect 137234 -8899 137621 -8877
rect 137158 -8925 137621 -8899
rect 137955 -8904 137956 -8637
rect 137971 -8688 138006 -8654
rect 138585 -8691 138620 -8657
rect 139264 -8663 139299 -8629
rect 139309 -8663 139310 -8618
rect 139409 -8629 139410 -8618
rect 139420 -8663 139455 -8629
rect 139465 -8663 139466 -8618
rect 139565 -8629 139566 -8618
rect 140143 -8623 140178 -8589
rect 140320 -8623 140355 -8589
rect 140681 -8605 140716 -8571
rect 139576 -8663 139611 -8629
rect 139409 -8697 139410 -8671
rect 139808 -8689 139843 -8655
rect 139853 -8689 139854 -8644
rect 139953 -8655 139954 -8644
rect 139964 -8689 139999 -8655
rect 140009 -8689 140010 -8644
rect 140309 -8672 140310 -8661
rect 137971 -8756 138006 -8722
rect 138174 -8770 138209 -8736
rect 138219 -8770 138220 -8728
rect 138319 -8740 138320 -8729
rect 138939 -8734 138974 -8700
rect 138330 -8774 138365 -8740
rect 138055 -8819 138056 -8808
rect 138524 -8813 138559 -8779
rect 138569 -8813 138570 -8771
rect 138669 -8779 138670 -8771
rect 139329 -8777 139364 -8743
rect 138680 -8813 138715 -8779
rect 138066 -8853 138101 -8819
rect 138174 -8870 138209 -8836
rect 138219 -8870 138220 -8825
rect 138319 -8832 138320 -8821
rect 138330 -8866 138365 -8832
rect 138878 -8856 138913 -8822
rect 138923 -8856 138924 -8814
rect 139023 -8822 139024 -8814
rect 139034 -8856 139069 -8822
rect 138067 -8906 138102 -8872
rect 138139 -8906 138174 -8872
rect 138211 -8906 138246 -8872
rect 138524 -8913 138559 -8879
rect 138569 -8913 138570 -8868
rect 138669 -8879 138670 -8868
rect 138680 -8913 138715 -8879
rect 139264 -8895 139299 -8861
rect 139309 -8895 139310 -8853
rect 137158 -8959 137634 -8925
rect 138492 -8949 138527 -8915
rect 138564 -8949 138599 -8915
rect 138878 -8956 138913 -8922
rect 138923 -8956 138924 -8911
rect 139023 -8922 139024 -8911
rect 139034 -8956 139069 -8922
rect 137158 -8985 137621 -8959
rect 137162 -8993 137363 -8985
rect 137178 -9003 137347 -8993
rect 136904 -9140 137079 -9114
rect 136411 -9174 136446 -9140
rect 136507 -9174 136542 -9140
rect 136603 -9174 136638 -9140
rect 136699 -9174 136734 -9140
rect 136795 -9174 136830 -9140
rect 136891 -9174 137079 -9140
rect 136904 -9200 137079 -9174
rect 137104 -9174 137205 -9050
rect 136982 -9870 137017 -9200
rect 137104 -9228 137107 -9174
rect 136789 -9936 136934 -9924
rect 136457 -9970 136934 -9936
rect 136789 -9971 136934 -9970
rect 136970 -9971 137017 -9870
rect 137116 -9971 137151 -9174
rect 137374 -9971 137409 -9062
rect 137508 -9971 137543 -8985
rect 137761 -9002 137796 -8968
rect 137857 -9002 137892 -8968
rect 137953 -9002 137988 -8968
rect 138049 -9002 138084 -8968
rect 138145 -9002 138180 -8968
rect 138241 -9002 138276 -8968
rect 138337 -9002 138372 -8968
rect 138846 -8992 138881 -8958
rect 138918 -8992 138953 -8958
rect 139264 -8995 139299 -8961
rect 139309 -8995 139310 -8950
rect 139451 -9001 139452 -8697
rect 140143 -8706 140178 -8672
rect 140320 -8706 140355 -8672
rect 140616 -8723 140651 -8689
rect 140661 -8723 140662 -8681
rect 140803 -8753 140804 -8525
rect 141493 -8534 141528 -8500
rect 141670 -8534 141705 -8500
rect 141864 -8577 141899 -8543
rect 141909 -8577 141910 -8532
rect 142009 -8543 142010 -8532
rect 142218 -8537 142253 -8503
rect 142263 -8537 142264 -8492
rect 142363 -8503 142364 -8492
rect 142608 -8496 142643 -8462
rect 142653 -8496 142654 -8451
rect 142753 -8462 142754 -8451
rect 142764 -8496 142799 -8462
rect 142809 -8496 142810 -8451
rect 142909 -8462 142910 -8451
rect 143090 -8456 143125 -8422
rect 143162 -8456 143197 -8422
rect 143234 -8456 143269 -8422
rect 143378 -8456 143413 -8422
rect 143450 -8456 143485 -8422
rect 143487 -8456 143557 -8422
rect 143594 -8456 143629 -8422
rect 143664 -8456 143699 -8422
rect 142920 -8496 142955 -8462
rect 143960 -8491 143995 -8457
rect 144005 -8491 144006 -8446
rect 144105 -8457 144106 -8446
rect 144116 -8491 144151 -8457
rect 144161 -8491 144162 -8446
rect 144261 -8457 144262 -8446
rect 144837 -8451 144872 -8417
rect 145014 -8451 145049 -8417
rect 144272 -8491 144307 -8457
rect 142374 -8537 142409 -8503
rect 143653 -8505 143654 -8494
rect 142020 -8577 142055 -8543
rect 140933 -8621 140968 -8587
rect 141134 -8666 141169 -8632
rect 141257 -8637 141258 -8595
rect 141579 -8624 141614 -8590
rect 142218 -8620 142253 -8586
rect 142263 -8620 142264 -8575
rect 142363 -8586 142364 -8575
rect 142608 -8580 142643 -8546
rect 142653 -8580 142654 -8535
rect 142753 -8546 142754 -8535
rect 142764 -8580 142799 -8546
rect 142809 -8580 142810 -8535
rect 142909 -8546 142910 -8535
rect 143487 -8539 143522 -8505
rect 143664 -8539 143699 -8505
rect 142920 -8580 142955 -8546
rect 143807 -8565 143922 -8499
rect 144105 -8525 144106 -8499
rect 144502 -8517 144537 -8483
rect 144547 -8517 144548 -8472
rect 144647 -8483 144648 -8472
rect 144658 -8517 144693 -8483
rect 144703 -8517 144704 -8472
rect 145003 -8500 145004 -8489
rect 145208 -8494 145243 -8460
rect 145253 -8494 145254 -8449
rect 145353 -8460 145354 -8449
rect 145562 -8453 145597 -8419
rect 145607 -8453 145608 -8408
rect 145707 -8419 145708 -8408
rect 145888 -8413 145923 -8379
rect 145952 -8413 145995 -8379
rect 145997 -8413 145998 -8371
rect 146097 -8379 146098 -8371
rect 146032 -8413 146067 -8379
rect 146108 -8413 146143 -8379
rect 146153 -8413 146154 -8371
rect 146253 -8379 146254 -8371
rect 146202 -8413 146237 -8379
rect 146264 -8413 146309 -8379
rect 147304 -8408 147339 -8374
rect 147349 -8408 147350 -8363
rect 147449 -8374 147450 -8363
rect 147460 -8408 147495 -8374
rect 147505 -8408 147506 -8363
rect 147605 -8374 147606 -8363
rect 148181 -8367 148216 -8333
rect 148358 -8367 148393 -8333
rect 148951 -8336 148952 -8328
rect 149051 -8336 149052 -8328
rect 147616 -8408 147651 -8374
rect 145718 -8453 145753 -8419
rect 146997 -8422 146998 -8414
rect 148347 -8417 148348 -8406
rect 148552 -8410 148587 -8376
rect 148597 -8410 148598 -8365
rect 148697 -8376 148698 -8365
rect 148878 -8370 148941 -8336
rect 148950 -8370 148985 -8336
rect 149062 -8370 149097 -8336
rect 149787 -8360 149822 -8326
rect 149883 -8360 149918 -8326
rect 149979 -8360 150014 -8326
rect 150075 -8360 150110 -8326
rect 150171 -8360 150206 -8326
rect 150267 -8360 150302 -8326
rect 150363 -8360 150398 -8326
rect 151691 -8333 151692 -8322
rect 151868 -8327 151931 -8293
rect 151940 -8327 151975 -8293
rect 152052 -8327 152087 -8293
rect 152583 -8317 152618 -8283
rect 152679 -8317 152714 -8283
rect 152775 -8317 152810 -8283
rect 152871 -8317 152906 -8283
rect 152967 -8317 153002 -8283
rect 153992 -8324 154027 -8290
rect 154037 -8324 154038 -8279
rect 154137 -8290 154138 -8279
rect 154148 -8324 154183 -8290
rect 154193 -8324 154194 -8279
rect 154293 -8290 154294 -8279
rect 154472 -8284 154507 -8250
rect 154544 -8284 154579 -8250
rect 154616 -8284 154651 -8250
rect 154760 -8284 154795 -8250
rect 154832 -8284 154867 -8250
rect 154869 -8284 154939 -8250
rect 154976 -8284 155011 -8250
rect 155046 -8284 155081 -8250
rect 155573 -8274 155608 -8240
rect 155669 -8274 155704 -8240
rect 155765 -8274 155800 -8240
rect 157272 -8241 157307 -8207
rect 157336 -8241 157379 -8207
rect 157381 -8241 157382 -8199
rect 157481 -8207 157482 -8199
rect 157416 -8241 157451 -8207
rect 157492 -8241 157527 -8207
rect 157537 -8241 157538 -8199
rect 157637 -8207 157638 -8199
rect 157586 -8241 157621 -8207
rect 157648 -8241 157693 -8207
rect 158563 -8231 158598 -8197
rect 158659 -8231 158694 -8197
rect 158755 -8231 158790 -8197
rect 158379 -8250 158380 -8242
rect 154304 -8324 154339 -8290
rect 155285 -8293 155286 -8285
rect 155385 -8293 155386 -8285
rect 148708 -8410 148743 -8376
rect 145364 -8494 145399 -8460
rect 142374 -8620 142409 -8586
rect 143653 -8589 143654 -8578
rect 140903 -8689 140904 -8681
rect 140914 -8723 140949 -8689
rect 141134 -8734 141169 -8700
rect 139581 -8793 139616 -8759
rect 139784 -8838 139819 -8804
rect 139907 -8809 139908 -8767
rect 140229 -8796 140264 -8762
rect 139551 -8861 139552 -8853
rect 139562 -8895 139597 -8861
rect 139784 -8906 139819 -8872
rect 139551 -8961 139552 -8950
rect 139562 -8995 139597 -8961
rect 138499 -9045 138534 -9011
rect 138595 -9045 138630 -9011
rect 138691 -9045 138726 -9011
rect 139200 -9035 139235 -9001
rect 139272 -9035 139307 -9001
rect 139344 -9035 139379 -9001
rect 139416 -9029 139452 -9001
rect 139762 -9025 139797 -8991
rect 139807 -9025 139808 -8980
rect 139416 -9035 139451 -9029
rect 138853 -9088 138888 -9054
rect 138949 -9088 138984 -9054
rect 139045 -9088 139080 -9054
rect 139949 -9076 139950 -8809
rect 140578 -8819 140965 -8753
rect 139965 -8860 140000 -8826
rect 140314 -8832 140325 -8819
rect 140248 -8874 140325 -8832
rect 140376 -8874 140965 -8819
rect 141112 -8853 141147 -8819
rect 141157 -8853 141158 -8808
rect 140248 -8877 140965 -8874
rect 139965 -8928 140000 -8894
rect 140168 -8942 140203 -8908
rect 140213 -8942 140214 -8900
rect 140049 -8991 140050 -8980
rect 140060 -9025 140095 -8991
rect 140168 -9042 140203 -9008
rect 140213 -9042 140214 -8997
rect 140061 -9078 140096 -9044
rect 140133 -9078 140168 -9044
rect 140205 -9078 140240 -9044
rect 139207 -9131 139242 -9097
rect 139303 -9131 139338 -9097
rect 139399 -9131 139434 -9097
rect 139495 -9131 139530 -9097
rect 139591 -9131 139626 -9097
rect 140248 -9114 140393 -8877
rect 140578 -8899 140965 -8877
rect 140502 -8925 140965 -8899
rect 141299 -8904 141300 -8637
rect 141315 -8688 141350 -8654
rect 141929 -8691 141964 -8657
rect 142608 -8663 142643 -8629
rect 142653 -8663 142654 -8618
rect 142753 -8629 142754 -8618
rect 142764 -8663 142799 -8629
rect 142809 -8663 142810 -8618
rect 142909 -8629 142910 -8618
rect 143487 -8623 143522 -8589
rect 143664 -8623 143699 -8589
rect 144025 -8605 144060 -8571
rect 142920 -8663 142955 -8629
rect 142753 -8697 142754 -8671
rect 143152 -8689 143187 -8655
rect 143197 -8689 143198 -8644
rect 143297 -8655 143298 -8644
rect 143308 -8689 143343 -8655
rect 143353 -8689 143354 -8644
rect 143653 -8672 143654 -8661
rect 141315 -8756 141350 -8722
rect 141518 -8770 141553 -8736
rect 141563 -8770 141564 -8728
rect 141663 -8740 141664 -8729
rect 142283 -8734 142318 -8700
rect 141674 -8774 141709 -8740
rect 141399 -8819 141400 -8808
rect 141868 -8813 141903 -8779
rect 141913 -8813 141914 -8771
rect 142013 -8779 142014 -8771
rect 142673 -8777 142708 -8743
rect 142024 -8813 142059 -8779
rect 141410 -8853 141445 -8819
rect 141518 -8870 141553 -8836
rect 141563 -8870 141564 -8825
rect 141663 -8832 141664 -8821
rect 141674 -8866 141709 -8832
rect 142222 -8856 142257 -8822
rect 142267 -8856 142268 -8814
rect 142367 -8822 142368 -8814
rect 142378 -8856 142413 -8822
rect 141411 -8906 141446 -8872
rect 141483 -8906 141518 -8872
rect 141555 -8906 141590 -8872
rect 141868 -8913 141903 -8879
rect 141913 -8913 141914 -8868
rect 142013 -8879 142014 -8868
rect 142024 -8913 142059 -8879
rect 142608 -8895 142643 -8861
rect 142653 -8895 142654 -8853
rect 140502 -8959 140978 -8925
rect 141836 -8949 141871 -8915
rect 141908 -8949 141943 -8915
rect 142222 -8956 142257 -8922
rect 142267 -8956 142268 -8911
rect 142367 -8922 142368 -8911
rect 142378 -8956 142413 -8922
rect 140502 -8985 140965 -8959
rect 140506 -8993 140707 -8985
rect 140522 -9003 140691 -8993
rect 140248 -9140 140423 -9114
rect 139755 -9174 139790 -9140
rect 139851 -9174 139886 -9140
rect 139947 -9174 139982 -9140
rect 140043 -9174 140078 -9140
rect 140139 -9174 140174 -9140
rect 140235 -9174 140423 -9140
rect 140248 -9200 140423 -9174
rect 140448 -9174 140549 -9050
rect 140326 -9870 140361 -9200
rect 140448 -9228 140451 -9174
rect 140133 -9936 140278 -9924
rect 139801 -9970 140278 -9936
rect 140133 -9971 140278 -9970
rect 140314 -9971 140361 -9870
rect 140460 -9971 140495 -9174
rect 140718 -9971 140753 -9062
rect 140852 -9971 140887 -8985
rect 141105 -9002 141140 -8968
rect 141201 -9002 141236 -8968
rect 141297 -9002 141332 -8968
rect 141393 -9002 141428 -8968
rect 141489 -9002 141524 -8968
rect 141585 -9002 141620 -8968
rect 141681 -9002 141716 -8968
rect 142190 -8992 142225 -8958
rect 142262 -8992 142297 -8958
rect 142608 -8995 142643 -8961
rect 142653 -8995 142654 -8950
rect 142795 -9001 142796 -8697
rect 143487 -8706 143522 -8672
rect 143664 -8706 143699 -8672
rect 143960 -8723 143995 -8689
rect 144005 -8723 144006 -8681
rect 144147 -8753 144148 -8525
rect 144837 -8534 144872 -8500
rect 145014 -8534 145049 -8500
rect 145208 -8577 145243 -8543
rect 145253 -8577 145254 -8532
rect 145353 -8543 145354 -8532
rect 145562 -8537 145597 -8503
rect 145607 -8537 145608 -8492
rect 145707 -8503 145708 -8492
rect 145952 -8496 145987 -8462
rect 145997 -8496 145998 -8451
rect 146097 -8462 146098 -8451
rect 146108 -8496 146143 -8462
rect 146153 -8496 146154 -8451
rect 146253 -8462 146254 -8451
rect 146434 -8456 146469 -8422
rect 146506 -8456 146541 -8422
rect 146578 -8456 146613 -8422
rect 146722 -8456 146757 -8422
rect 146794 -8456 146829 -8422
rect 146831 -8456 146901 -8422
rect 146938 -8456 146973 -8422
rect 147008 -8456 147043 -8422
rect 146264 -8496 146299 -8462
rect 147304 -8491 147339 -8457
rect 147349 -8491 147350 -8446
rect 147449 -8457 147450 -8446
rect 147460 -8491 147495 -8457
rect 147505 -8491 147506 -8446
rect 147605 -8457 147606 -8446
rect 148181 -8451 148216 -8417
rect 148358 -8451 148393 -8417
rect 147616 -8491 147651 -8457
rect 145718 -8537 145753 -8503
rect 146997 -8505 146998 -8494
rect 145364 -8577 145399 -8543
rect 144277 -8621 144312 -8587
rect 144478 -8666 144513 -8632
rect 144601 -8637 144602 -8595
rect 144923 -8624 144958 -8590
rect 145562 -8620 145597 -8586
rect 145607 -8620 145608 -8575
rect 145707 -8586 145708 -8575
rect 145952 -8580 145987 -8546
rect 145997 -8580 145998 -8535
rect 146097 -8546 146098 -8535
rect 146108 -8580 146143 -8546
rect 146153 -8580 146154 -8535
rect 146253 -8546 146254 -8535
rect 146831 -8539 146866 -8505
rect 147008 -8539 147043 -8505
rect 146264 -8580 146299 -8546
rect 147151 -8565 147266 -8499
rect 147449 -8525 147450 -8499
rect 147846 -8517 147881 -8483
rect 147891 -8517 147892 -8472
rect 147991 -8483 147992 -8472
rect 148002 -8517 148037 -8483
rect 148047 -8517 148048 -8472
rect 148347 -8500 148348 -8489
rect 148552 -8494 148587 -8460
rect 148597 -8494 148598 -8449
rect 148697 -8460 148698 -8449
rect 148906 -8453 148941 -8419
rect 148951 -8453 148952 -8408
rect 149051 -8419 149052 -8408
rect 149232 -8413 149267 -8379
rect 149296 -8413 149339 -8379
rect 149341 -8413 149342 -8371
rect 149441 -8379 149442 -8371
rect 149376 -8413 149411 -8379
rect 149452 -8413 149487 -8379
rect 149497 -8413 149498 -8371
rect 149597 -8379 149598 -8371
rect 149546 -8413 149581 -8379
rect 149608 -8413 149653 -8379
rect 150648 -8408 150683 -8374
rect 150693 -8408 150694 -8363
rect 150793 -8374 150794 -8363
rect 150804 -8408 150839 -8374
rect 150849 -8408 150850 -8363
rect 150949 -8374 150950 -8363
rect 151525 -8367 151560 -8333
rect 151702 -8367 151737 -8333
rect 152295 -8336 152296 -8328
rect 152395 -8336 152396 -8328
rect 150960 -8408 150995 -8374
rect 149062 -8453 149097 -8419
rect 150341 -8422 150342 -8414
rect 151691 -8417 151692 -8406
rect 151896 -8410 151931 -8376
rect 151941 -8410 151942 -8365
rect 152041 -8376 152042 -8365
rect 152222 -8370 152285 -8336
rect 152294 -8370 152329 -8336
rect 152406 -8370 152441 -8336
rect 153131 -8360 153166 -8326
rect 153227 -8360 153262 -8326
rect 153323 -8360 153358 -8326
rect 153419 -8360 153454 -8326
rect 153515 -8360 153550 -8326
rect 153611 -8360 153646 -8326
rect 153707 -8360 153742 -8326
rect 155035 -8333 155036 -8322
rect 155212 -8327 155275 -8293
rect 155284 -8327 155319 -8293
rect 155396 -8327 155431 -8293
rect 155927 -8317 155962 -8283
rect 156023 -8317 156058 -8283
rect 156119 -8317 156154 -8283
rect 156215 -8317 156250 -8283
rect 156311 -8317 156346 -8283
rect 157336 -8324 157371 -8290
rect 157381 -8324 157382 -8279
rect 157481 -8290 157482 -8279
rect 157492 -8324 157527 -8290
rect 157537 -8324 157538 -8279
rect 157637 -8290 157638 -8279
rect 157816 -8284 157851 -8250
rect 157888 -8284 157923 -8250
rect 157960 -8284 157995 -8250
rect 158104 -8284 158139 -8250
rect 158176 -8284 158211 -8250
rect 158213 -8284 158283 -8250
rect 158320 -8284 158355 -8250
rect 158390 -8284 158425 -8250
rect 158917 -8274 158952 -8240
rect 159013 -8274 159048 -8240
rect 159109 -8274 159144 -8240
rect 160616 -8241 160651 -8207
rect 160680 -8241 160723 -8207
rect 160725 -8241 160726 -8199
rect 160825 -8207 160826 -8199
rect 160760 -8241 160795 -8207
rect 160836 -8241 160871 -8207
rect 160881 -8241 160882 -8199
rect 160981 -8207 160982 -8199
rect 160930 -8241 160965 -8207
rect 160992 -8241 161037 -8207
rect 161907 -8231 161942 -8197
rect 162003 -8231 162038 -8197
rect 162099 -8231 162134 -8197
rect 161723 -8250 161724 -8242
rect 157648 -8324 157683 -8290
rect 158629 -8293 158630 -8285
rect 158729 -8293 158730 -8285
rect 152052 -8410 152087 -8376
rect 148708 -8494 148743 -8460
rect 145718 -8620 145753 -8586
rect 146997 -8589 146998 -8578
rect 144247 -8689 144248 -8681
rect 144258 -8723 144293 -8689
rect 144478 -8734 144513 -8700
rect 142925 -8793 142960 -8759
rect 143128 -8838 143163 -8804
rect 143251 -8809 143252 -8767
rect 143573 -8796 143608 -8762
rect 142895 -8861 142896 -8853
rect 142906 -8895 142941 -8861
rect 143128 -8906 143163 -8872
rect 142895 -8961 142896 -8950
rect 142906 -8995 142941 -8961
rect 141843 -9045 141878 -9011
rect 141939 -9045 141974 -9011
rect 142035 -9045 142070 -9011
rect 142544 -9035 142579 -9001
rect 142616 -9035 142651 -9001
rect 142688 -9035 142723 -9001
rect 142760 -9029 142796 -9001
rect 143106 -9025 143141 -8991
rect 143151 -9025 143152 -8980
rect 142760 -9035 142795 -9029
rect 142197 -9088 142232 -9054
rect 142293 -9088 142328 -9054
rect 142389 -9088 142424 -9054
rect 143293 -9076 143294 -8809
rect 143922 -8819 144309 -8753
rect 143309 -8860 143344 -8826
rect 143658 -8832 143669 -8819
rect 143592 -8874 143669 -8832
rect 143720 -8874 144309 -8819
rect 144456 -8853 144491 -8819
rect 144501 -8853 144502 -8808
rect 143592 -8877 144309 -8874
rect 143309 -8928 143344 -8894
rect 143512 -8942 143547 -8908
rect 143557 -8942 143558 -8900
rect 143393 -8991 143394 -8980
rect 143404 -9025 143439 -8991
rect 143512 -9042 143547 -9008
rect 143557 -9042 143558 -8997
rect 143405 -9078 143440 -9044
rect 143477 -9078 143512 -9044
rect 143549 -9078 143584 -9044
rect 142551 -9131 142586 -9097
rect 142647 -9131 142682 -9097
rect 142743 -9131 142778 -9097
rect 142839 -9131 142874 -9097
rect 142935 -9131 142970 -9097
rect 143592 -9114 143737 -8877
rect 143922 -8899 144309 -8877
rect 143846 -8925 144309 -8899
rect 144643 -8904 144644 -8637
rect 144659 -8688 144694 -8654
rect 145273 -8691 145308 -8657
rect 145952 -8663 145987 -8629
rect 145997 -8663 145998 -8618
rect 146097 -8629 146098 -8618
rect 146108 -8663 146143 -8629
rect 146153 -8663 146154 -8618
rect 146253 -8629 146254 -8618
rect 146831 -8623 146866 -8589
rect 147008 -8623 147043 -8589
rect 147369 -8605 147404 -8571
rect 146264 -8663 146299 -8629
rect 146097 -8697 146098 -8671
rect 146496 -8689 146531 -8655
rect 146541 -8689 146542 -8644
rect 146641 -8655 146642 -8644
rect 146652 -8689 146687 -8655
rect 146697 -8689 146698 -8644
rect 146997 -8672 146998 -8661
rect 144659 -8756 144694 -8722
rect 144862 -8770 144897 -8736
rect 144907 -8770 144908 -8728
rect 145007 -8740 145008 -8729
rect 145627 -8734 145662 -8700
rect 145018 -8774 145053 -8740
rect 144743 -8819 144744 -8808
rect 145212 -8813 145247 -8779
rect 145257 -8813 145258 -8771
rect 145357 -8779 145358 -8771
rect 146017 -8777 146052 -8743
rect 145368 -8813 145403 -8779
rect 144754 -8853 144789 -8819
rect 144862 -8870 144897 -8836
rect 144907 -8870 144908 -8825
rect 145007 -8832 145008 -8821
rect 145018 -8866 145053 -8832
rect 145566 -8856 145601 -8822
rect 145611 -8856 145612 -8814
rect 145711 -8822 145712 -8814
rect 145722 -8856 145757 -8822
rect 144755 -8906 144790 -8872
rect 144827 -8906 144862 -8872
rect 144899 -8906 144934 -8872
rect 145212 -8913 145247 -8879
rect 145257 -8913 145258 -8868
rect 145357 -8879 145358 -8868
rect 145368 -8913 145403 -8879
rect 145952 -8895 145987 -8861
rect 145997 -8895 145998 -8853
rect 143846 -8959 144322 -8925
rect 145180 -8949 145215 -8915
rect 145252 -8949 145287 -8915
rect 145566 -8956 145601 -8922
rect 145611 -8956 145612 -8911
rect 145711 -8922 145712 -8911
rect 145722 -8956 145757 -8922
rect 143846 -8985 144309 -8959
rect 143850 -8993 144051 -8985
rect 143866 -9003 144035 -8993
rect 143592 -9140 143767 -9114
rect 143099 -9174 143134 -9140
rect 143195 -9174 143230 -9140
rect 143291 -9174 143326 -9140
rect 143387 -9174 143422 -9140
rect 143483 -9174 143518 -9140
rect 143579 -9174 143767 -9140
rect 143592 -9200 143767 -9174
rect 143792 -9174 143893 -9050
rect 143670 -9870 143705 -9200
rect 143792 -9228 143795 -9174
rect 143477 -9936 143622 -9924
rect 143145 -9970 143622 -9936
rect 143477 -9971 143622 -9970
rect 143658 -9971 143705 -9870
rect 143804 -9971 143839 -9174
rect 144062 -9971 144097 -9062
rect 144196 -9971 144231 -8985
rect 144449 -9002 144484 -8968
rect 144545 -9002 144580 -8968
rect 144641 -9002 144676 -8968
rect 144737 -9002 144772 -8968
rect 144833 -9002 144868 -8968
rect 144929 -9002 144964 -8968
rect 145025 -9002 145060 -8968
rect 145534 -8992 145569 -8958
rect 145606 -8992 145641 -8958
rect 145952 -8995 145987 -8961
rect 145997 -8995 145998 -8950
rect 146139 -9001 146140 -8697
rect 146831 -8706 146866 -8672
rect 147008 -8706 147043 -8672
rect 147304 -8723 147339 -8689
rect 147349 -8723 147350 -8681
rect 147491 -8753 147492 -8525
rect 148181 -8534 148216 -8500
rect 148358 -8534 148393 -8500
rect 148552 -8577 148587 -8543
rect 148597 -8577 148598 -8532
rect 148697 -8543 148698 -8532
rect 148906 -8537 148941 -8503
rect 148951 -8537 148952 -8492
rect 149051 -8503 149052 -8492
rect 149296 -8496 149331 -8462
rect 149341 -8496 149342 -8451
rect 149441 -8462 149442 -8451
rect 149452 -8496 149487 -8462
rect 149497 -8496 149498 -8451
rect 149597 -8462 149598 -8451
rect 149778 -8456 149813 -8422
rect 149850 -8456 149885 -8422
rect 149922 -8456 149957 -8422
rect 150066 -8456 150101 -8422
rect 150138 -8456 150173 -8422
rect 150175 -8456 150245 -8422
rect 150282 -8456 150317 -8422
rect 150352 -8456 150387 -8422
rect 149608 -8496 149643 -8462
rect 150648 -8491 150683 -8457
rect 150693 -8491 150694 -8446
rect 150793 -8457 150794 -8446
rect 150804 -8491 150839 -8457
rect 150849 -8491 150850 -8446
rect 150949 -8457 150950 -8446
rect 151525 -8451 151560 -8417
rect 151702 -8451 151737 -8417
rect 150960 -8491 150995 -8457
rect 149062 -8537 149097 -8503
rect 150341 -8505 150342 -8494
rect 148708 -8577 148743 -8543
rect 147621 -8621 147656 -8587
rect 147822 -8666 147857 -8632
rect 147945 -8637 147946 -8595
rect 148267 -8624 148302 -8590
rect 148906 -8620 148941 -8586
rect 148951 -8620 148952 -8575
rect 149051 -8586 149052 -8575
rect 149296 -8580 149331 -8546
rect 149341 -8580 149342 -8535
rect 149441 -8546 149442 -8535
rect 149452 -8580 149487 -8546
rect 149497 -8580 149498 -8535
rect 149597 -8546 149598 -8535
rect 150175 -8539 150210 -8505
rect 150352 -8539 150387 -8505
rect 149608 -8580 149643 -8546
rect 150495 -8565 150610 -8499
rect 150793 -8525 150794 -8499
rect 151190 -8517 151225 -8483
rect 151235 -8517 151236 -8472
rect 151335 -8483 151336 -8472
rect 151346 -8517 151381 -8483
rect 151391 -8517 151392 -8472
rect 151691 -8500 151692 -8489
rect 151896 -8494 151931 -8460
rect 151941 -8494 151942 -8449
rect 152041 -8460 152042 -8449
rect 152250 -8453 152285 -8419
rect 152295 -8453 152296 -8408
rect 152395 -8419 152396 -8408
rect 152576 -8413 152611 -8379
rect 152640 -8413 152683 -8379
rect 152685 -8413 152686 -8371
rect 152785 -8379 152786 -8371
rect 152720 -8413 152755 -8379
rect 152796 -8413 152831 -8379
rect 152841 -8413 152842 -8371
rect 152941 -8379 152942 -8371
rect 152890 -8413 152925 -8379
rect 152952 -8413 152997 -8379
rect 153992 -8408 154027 -8374
rect 154037 -8408 154038 -8363
rect 154137 -8374 154138 -8363
rect 154148 -8408 154183 -8374
rect 154193 -8408 154194 -8363
rect 154293 -8374 154294 -8363
rect 154869 -8367 154904 -8333
rect 155046 -8367 155081 -8333
rect 155639 -8336 155640 -8328
rect 155739 -8336 155740 -8328
rect 154304 -8408 154339 -8374
rect 152406 -8453 152441 -8419
rect 153685 -8422 153686 -8414
rect 155035 -8417 155036 -8406
rect 155240 -8410 155275 -8376
rect 155285 -8410 155286 -8365
rect 155385 -8376 155386 -8365
rect 155566 -8370 155629 -8336
rect 155638 -8370 155673 -8336
rect 155750 -8370 155785 -8336
rect 156475 -8360 156510 -8326
rect 156571 -8360 156606 -8326
rect 156667 -8360 156702 -8326
rect 156763 -8360 156798 -8326
rect 156859 -8360 156894 -8326
rect 156955 -8360 156990 -8326
rect 157051 -8360 157086 -8326
rect 158379 -8333 158380 -8322
rect 158556 -8327 158619 -8293
rect 158628 -8327 158663 -8293
rect 158740 -8327 158775 -8293
rect 159271 -8317 159306 -8283
rect 159367 -8317 159402 -8283
rect 159463 -8317 159498 -8283
rect 159559 -8317 159594 -8283
rect 159655 -8317 159690 -8283
rect 160680 -8324 160715 -8290
rect 160725 -8324 160726 -8279
rect 160825 -8290 160826 -8279
rect 160836 -8324 160871 -8290
rect 160881 -8324 160882 -8279
rect 160981 -8290 160982 -8279
rect 161160 -8284 161195 -8250
rect 161232 -8284 161267 -8250
rect 161304 -8284 161339 -8250
rect 161448 -8284 161483 -8250
rect 161520 -8284 161555 -8250
rect 161557 -8284 161627 -8250
rect 161664 -8284 161699 -8250
rect 161734 -8284 161769 -8250
rect 162261 -8274 162296 -8240
rect 162357 -8274 162392 -8240
rect 162453 -8274 162488 -8240
rect 163960 -8241 163995 -8207
rect 164024 -8241 164067 -8207
rect 164069 -8241 164070 -8199
rect 164169 -8207 164170 -8199
rect 164104 -8241 164139 -8207
rect 164180 -8241 164215 -8207
rect 164225 -8241 164226 -8199
rect 164325 -8207 164326 -8199
rect 164274 -8241 164309 -8207
rect 164336 -8241 164381 -8207
rect 165251 -8231 165286 -8197
rect 165347 -8231 165382 -8197
rect 165443 -8231 165478 -8197
rect 165067 -8250 165068 -8242
rect 160992 -8324 161027 -8290
rect 161973 -8293 161974 -8285
rect 162073 -8293 162074 -8285
rect 155396 -8410 155431 -8376
rect 152052 -8494 152087 -8460
rect 149062 -8620 149097 -8586
rect 150341 -8589 150342 -8578
rect 147591 -8689 147592 -8681
rect 147602 -8723 147637 -8689
rect 147822 -8734 147857 -8700
rect 146269 -8793 146304 -8759
rect 146472 -8838 146507 -8804
rect 146595 -8809 146596 -8767
rect 146917 -8796 146952 -8762
rect 146239 -8861 146240 -8853
rect 146250 -8895 146285 -8861
rect 146472 -8906 146507 -8872
rect 146239 -8961 146240 -8950
rect 146250 -8995 146285 -8961
rect 145187 -9045 145222 -9011
rect 145283 -9045 145318 -9011
rect 145379 -9045 145414 -9011
rect 145888 -9035 145923 -9001
rect 145960 -9035 145995 -9001
rect 146032 -9035 146067 -9001
rect 146104 -9029 146140 -9001
rect 146450 -9025 146485 -8991
rect 146495 -9025 146496 -8980
rect 146104 -9035 146139 -9029
rect 145541 -9088 145576 -9054
rect 145637 -9088 145672 -9054
rect 145733 -9088 145768 -9054
rect 146637 -9076 146638 -8809
rect 147266 -8819 147653 -8753
rect 146653 -8860 146688 -8826
rect 147002 -8832 147013 -8819
rect 146936 -8874 147013 -8832
rect 147064 -8874 147653 -8819
rect 147800 -8853 147835 -8819
rect 147845 -8853 147846 -8808
rect 146936 -8877 147653 -8874
rect 146653 -8928 146688 -8894
rect 146856 -8942 146891 -8908
rect 146901 -8942 146902 -8900
rect 146737 -8991 146738 -8980
rect 146748 -9025 146783 -8991
rect 146856 -9042 146891 -9008
rect 146901 -9042 146902 -8997
rect 146749 -9078 146784 -9044
rect 146821 -9078 146856 -9044
rect 146893 -9078 146928 -9044
rect 145895 -9131 145930 -9097
rect 145991 -9131 146026 -9097
rect 146087 -9131 146122 -9097
rect 146183 -9131 146218 -9097
rect 146279 -9131 146314 -9097
rect 146936 -9114 147081 -8877
rect 147266 -8899 147653 -8877
rect 147190 -8925 147653 -8899
rect 147987 -8904 147988 -8637
rect 148003 -8688 148038 -8654
rect 148617 -8691 148652 -8657
rect 149296 -8663 149331 -8629
rect 149341 -8663 149342 -8618
rect 149441 -8629 149442 -8618
rect 149452 -8663 149487 -8629
rect 149497 -8663 149498 -8618
rect 149597 -8629 149598 -8618
rect 150175 -8623 150210 -8589
rect 150352 -8623 150387 -8589
rect 150713 -8605 150748 -8571
rect 149608 -8663 149643 -8629
rect 149441 -8697 149442 -8671
rect 149840 -8689 149875 -8655
rect 149885 -8689 149886 -8644
rect 149985 -8655 149986 -8644
rect 149996 -8689 150031 -8655
rect 150041 -8689 150042 -8644
rect 150341 -8672 150342 -8661
rect 148003 -8756 148038 -8722
rect 148206 -8770 148241 -8736
rect 148251 -8770 148252 -8728
rect 148351 -8740 148352 -8729
rect 148971 -8734 149006 -8700
rect 148362 -8774 148397 -8740
rect 148087 -8819 148088 -8808
rect 148556 -8813 148591 -8779
rect 148601 -8813 148602 -8771
rect 148701 -8779 148702 -8771
rect 149361 -8777 149396 -8743
rect 148712 -8813 148747 -8779
rect 148098 -8853 148133 -8819
rect 148206 -8870 148241 -8836
rect 148251 -8870 148252 -8825
rect 148351 -8832 148352 -8821
rect 148362 -8866 148397 -8832
rect 148910 -8856 148945 -8822
rect 148955 -8856 148956 -8814
rect 149055 -8822 149056 -8814
rect 149066 -8856 149101 -8822
rect 148099 -8906 148134 -8872
rect 148171 -8906 148206 -8872
rect 148243 -8906 148278 -8872
rect 148556 -8913 148591 -8879
rect 148601 -8913 148602 -8868
rect 148701 -8879 148702 -8868
rect 148712 -8913 148747 -8879
rect 149296 -8895 149331 -8861
rect 149341 -8895 149342 -8853
rect 147190 -8959 147666 -8925
rect 148524 -8949 148559 -8915
rect 148596 -8949 148631 -8915
rect 148910 -8956 148945 -8922
rect 148955 -8956 148956 -8911
rect 149055 -8922 149056 -8911
rect 149066 -8956 149101 -8922
rect 147190 -8985 147653 -8959
rect 147194 -8993 147395 -8985
rect 147210 -9003 147379 -8993
rect 146936 -9140 147111 -9114
rect 146443 -9174 146478 -9140
rect 146539 -9174 146574 -9140
rect 146635 -9174 146670 -9140
rect 146731 -9174 146766 -9140
rect 146827 -9174 146862 -9140
rect 146923 -9174 147111 -9140
rect 146936 -9200 147111 -9174
rect 147136 -9174 147237 -9050
rect 147014 -9870 147049 -9200
rect 147136 -9228 147139 -9174
rect 146821 -9936 146966 -9924
rect 146489 -9970 146966 -9936
rect 146821 -9971 146966 -9970
rect 147002 -9971 147049 -9870
rect 147148 -9971 147183 -9174
rect 147406 -9971 147441 -9062
rect 147540 -9971 147575 -8985
rect 147793 -9002 147828 -8968
rect 147889 -9002 147924 -8968
rect 147985 -9002 148020 -8968
rect 148081 -9002 148116 -8968
rect 148177 -9002 148212 -8968
rect 148273 -9002 148308 -8968
rect 148369 -9002 148404 -8968
rect 148878 -8992 148913 -8958
rect 148950 -8992 148985 -8958
rect 149296 -8995 149331 -8961
rect 149341 -8995 149342 -8950
rect 149483 -9001 149484 -8697
rect 150175 -8706 150210 -8672
rect 150352 -8706 150387 -8672
rect 150648 -8723 150683 -8689
rect 150693 -8723 150694 -8681
rect 150835 -8753 150836 -8525
rect 151525 -8534 151560 -8500
rect 151702 -8534 151737 -8500
rect 151896 -8577 151931 -8543
rect 151941 -8577 151942 -8532
rect 152041 -8543 152042 -8532
rect 152250 -8537 152285 -8503
rect 152295 -8537 152296 -8492
rect 152395 -8503 152396 -8492
rect 152640 -8496 152675 -8462
rect 152685 -8496 152686 -8451
rect 152785 -8462 152786 -8451
rect 152796 -8496 152831 -8462
rect 152841 -8496 152842 -8451
rect 152941 -8462 152942 -8451
rect 153122 -8456 153157 -8422
rect 153194 -8456 153229 -8422
rect 153266 -8456 153301 -8422
rect 153410 -8456 153445 -8422
rect 153482 -8456 153517 -8422
rect 153519 -8456 153589 -8422
rect 153626 -8456 153661 -8422
rect 153696 -8456 153731 -8422
rect 152952 -8496 152987 -8462
rect 153992 -8491 154027 -8457
rect 154037 -8491 154038 -8446
rect 154137 -8457 154138 -8446
rect 154148 -8491 154183 -8457
rect 154193 -8491 154194 -8446
rect 154293 -8457 154294 -8446
rect 154869 -8451 154904 -8417
rect 155046 -8451 155081 -8417
rect 154304 -8491 154339 -8457
rect 152406 -8537 152441 -8503
rect 153685 -8505 153686 -8494
rect 152052 -8577 152087 -8543
rect 150965 -8621 151000 -8587
rect 151166 -8666 151201 -8632
rect 151289 -8637 151290 -8595
rect 151611 -8624 151646 -8590
rect 152250 -8620 152285 -8586
rect 152295 -8620 152296 -8575
rect 152395 -8586 152396 -8575
rect 152640 -8580 152675 -8546
rect 152685 -8580 152686 -8535
rect 152785 -8546 152786 -8535
rect 152796 -8580 152831 -8546
rect 152841 -8580 152842 -8535
rect 152941 -8546 152942 -8535
rect 153519 -8539 153554 -8505
rect 153696 -8539 153731 -8505
rect 152952 -8580 152987 -8546
rect 153839 -8565 153954 -8499
rect 154137 -8525 154138 -8499
rect 154534 -8517 154569 -8483
rect 154579 -8517 154580 -8472
rect 154679 -8483 154680 -8472
rect 154690 -8517 154725 -8483
rect 154735 -8517 154736 -8472
rect 155035 -8500 155036 -8489
rect 155240 -8494 155275 -8460
rect 155285 -8494 155286 -8449
rect 155385 -8460 155386 -8449
rect 155594 -8453 155629 -8419
rect 155639 -8453 155640 -8408
rect 155739 -8419 155740 -8408
rect 155920 -8413 155955 -8379
rect 155984 -8413 156027 -8379
rect 156029 -8413 156030 -8371
rect 156129 -8379 156130 -8371
rect 156064 -8413 156099 -8379
rect 156140 -8413 156175 -8379
rect 156185 -8413 156186 -8371
rect 156285 -8379 156286 -8371
rect 156234 -8413 156269 -8379
rect 156296 -8413 156341 -8379
rect 157336 -8408 157371 -8374
rect 157381 -8408 157382 -8363
rect 157481 -8374 157482 -8363
rect 157492 -8408 157527 -8374
rect 157537 -8408 157538 -8363
rect 157637 -8374 157638 -8363
rect 158213 -8367 158248 -8333
rect 158390 -8367 158425 -8333
rect 158983 -8336 158984 -8328
rect 159083 -8336 159084 -8328
rect 157648 -8408 157683 -8374
rect 155750 -8453 155785 -8419
rect 157029 -8422 157030 -8414
rect 158379 -8417 158380 -8406
rect 158584 -8410 158619 -8376
rect 158629 -8410 158630 -8365
rect 158729 -8376 158730 -8365
rect 158910 -8370 158973 -8336
rect 158982 -8370 159017 -8336
rect 159094 -8370 159129 -8336
rect 159819 -8360 159854 -8326
rect 159915 -8360 159950 -8326
rect 160011 -8360 160046 -8326
rect 160107 -8360 160142 -8326
rect 160203 -8360 160238 -8326
rect 160299 -8360 160334 -8326
rect 160395 -8360 160430 -8326
rect 161723 -8333 161724 -8322
rect 161900 -8327 161963 -8293
rect 161972 -8327 162007 -8293
rect 162084 -8327 162119 -8293
rect 162615 -8317 162650 -8283
rect 162711 -8317 162746 -8283
rect 162807 -8317 162842 -8283
rect 162903 -8317 162938 -8283
rect 162999 -8317 163034 -8283
rect 164024 -8324 164059 -8290
rect 164069 -8324 164070 -8279
rect 164169 -8290 164170 -8279
rect 164180 -8324 164215 -8290
rect 164225 -8324 164226 -8279
rect 164325 -8290 164326 -8279
rect 164504 -8284 164539 -8250
rect 164576 -8284 164611 -8250
rect 164648 -8284 164683 -8250
rect 164792 -8284 164827 -8250
rect 164864 -8284 164899 -8250
rect 164901 -8284 164971 -8250
rect 165008 -8284 165043 -8250
rect 165078 -8284 165113 -8250
rect 165605 -8274 165640 -8240
rect 165701 -8274 165736 -8240
rect 165797 -8274 165832 -8240
rect 167304 -8241 167339 -8207
rect 167368 -8241 167411 -8207
rect 167413 -8241 167414 -8199
rect 167513 -8207 167514 -8199
rect 167448 -8241 167483 -8207
rect 167524 -8241 167559 -8207
rect 167569 -8241 167570 -8199
rect 167669 -8207 167670 -8199
rect 167618 -8241 167653 -8207
rect 167680 -8241 167725 -8207
rect 168595 -8231 168630 -8197
rect 168691 -8231 168726 -8197
rect 168787 -8231 168822 -8197
rect 168411 -8250 168412 -8242
rect 164336 -8324 164371 -8290
rect 165317 -8293 165318 -8285
rect 165417 -8293 165418 -8285
rect 158740 -8410 158775 -8376
rect 155396 -8494 155431 -8460
rect 152406 -8620 152441 -8586
rect 153685 -8589 153686 -8578
rect 150935 -8689 150936 -8681
rect 150946 -8723 150981 -8689
rect 151166 -8734 151201 -8700
rect 149613 -8793 149648 -8759
rect 149816 -8838 149851 -8804
rect 149939 -8809 149940 -8767
rect 150261 -8796 150296 -8762
rect 149583 -8861 149584 -8853
rect 149594 -8895 149629 -8861
rect 149816 -8906 149851 -8872
rect 149583 -8961 149584 -8950
rect 149594 -8995 149629 -8961
rect 148531 -9045 148566 -9011
rect 148627 -9045 148662 -9011
rect 148723 -9045 148758 -9011
rect 149232 -9035 149267 -9001
rect 149304 -9035 149339 -9001
rect 149376 -9035 149411 -9001
rect 149448 -9029 149484 -9001
rect 149794 -9025 149829 -8991
rect 149839 -9025 149840 -8980
rect 149448 -9035 149483 -9029
rect 148885 -9088 148920 -9054
rect 148981 -9088 149016 -9054
rect 149077 -9088 149112 -9054
rect 149981 -9076 149982 -8809
rect 150610 -8819 150997 -8753
rect 149997 -8860 150032 -8826
rect 150346 -8832 150357 -8819
rect 150280 -8874 150357 -8832
rect 150408 -8874 150997 -8819
rect 151144 -8853 151179 -8819
rect 151189 -8853 151190 -8808
rect 150280 -8877 150997 -8874
rect 149997 -8928 150032 -8894
rect 150200 -8942 150235 -8908
rect 150245 -8942 150246 -8900
rect 150081 -8991 150082 -8980
rect 150092 -9025 150127 -8991
rect 150200 -9042 150235 -9008
rect 150245 -9042 150246 -8997
rect 150093 -9078 150128 -9044
rect 150165 -9078 150200 -9044
rect 150237 -9078 150272 -9044
rect 149239 -9131 149274 -9097
rect 149335 -9131 149370 -9097
rect 149431 -9131 149466 -9097
rect 149527 -9131 149562 -9097
rect 149623 -9131 149658 -9097
rect 150280 -9114 150425 -8877
rect 150610 -8899 150997 -8877
rect 150534 -8925 150997 -8899
rect 151331 -8904 151332 -8637
rect 151347 -8688 151382 -8654
rect 151961 -8691 151996 -8657
rect 152640 -8663 152675 -8629
rect 152685 -8663 152686 -8618
rect 152785 -8629 152786 -8618
rect 152796 -8663 152831 -8629
rect 152841 -8663 152842 -8618
rect 152941 -8629 152942 -8618
rect 153519 -8623 153554 -8589
rect 153696 -8623 153731 -8589
rect 154057 -8605 154092 -8571
rect 152952 -8663 152987 -8629
rect 152785 -8697 152786 -8671
rect 153184 -8689 153219 -8655
rect 153229 -8689 153230 -8644
rect 153329 -8655 153330 -8644
rect 153340 -8689 153375 -8655
rect 153385 -8689 153386 -8644
rect 153685 -8672 153686 -8661
rect 151347 -8756 151382 -8722
rect 151550 -8770 151585 -8736
rect 151595 -8770 151596 -8728
rect 151695 -8740 151696 -8729
rect 152315 -8734 152350 -8700
rect 151706 -8774 151741 -8740
rect 151431 -8819 151432 -8808
rect 151900 -8813 151935 -8779
rect 151945 -8813 151946 -8771
rect 152045 -8779 152046 -8771
rect 152705 -8777 152740 -8743
rect 152056 -8813 152091 -8779
rect 151442 -8853 151477 -8819
rect 151550 -8870 151585 -8836
rect 151595 -8870 151596 -8825
rect 151695 -8832 151696 -8821
rect 151706 -8866 151741 -8832
rect 152254 -8856 152289 -8822
rect 152299 -8856 152300 -8814
rect 152399 -8822 152400 -8814
rect 152410 -8856 152445 -8822
rect 151443 -8906 151478 -8872
rect 151515 -8906 151550 -8872
rect 151587 -8906 151622 -8872
rect 151900 -8913 151935 -8879
rect 151945 -8913 151946 -8868
rect 152045 -8879 152046 -8868
rect 152056 -8913 152091 -8879
rect 152640 -8895 152675 -8861
rect 152685 -8895 152686 -8853
rect 150534 -8959 151010 -8925
rect 151868 -8949 151903 -8915
rect 151940 -8949 151975 -8915
rect 152254 -8956 152289 -8922
rect 152299 -8956 152300 -8911
rect 152399 -8922 152400 -8911
rect 152410 -8956 152445 -8922
rect 150534 -8985 150997 -8959
rect 150538 -8993 150739 -8985
rect 150554 -9003 150723 -8993
rect 150280 -9140 150455 -9114
rect 149787 -9174 149822 -9140
rect 149883 -9174 149918 -9140
rect 149979 -9174 150014 -9140
rect 150075 -9174 150110 -9140
rect 150171 -9174 150206 -9140
rect 150267 -9174 150455 -9140
rect 150280 -9200 150455 -9174
rect 150480 -9174 150581 -9050
rect 150358 -9870 150393 -9200
rect 150480 -9228 150483 -9174
rect 150165 -9936 150310 -9924
rect 149833 -9970 150310 -9936
rect 150165 -9971 150310 -9970
rect 150346 -9971 150393 -9870
rect 150492 -9971 150527 -9174
rect 150750 -9971 150785 -9062
rect 150884 -9971 150919 -8985
rect 151137 -9002 151172 -8968
rect 151233 -9002 151268 -8968
rect 151329 -9002 151364 -8968
rect 151425 -9002 151460 -8968
rect 151521 -9002 151556 -8968
rect 151617 -9002 151652 -8968
rect 151713 -9002 151748 -8968
rect 152222 -8992 152257 -8958
rect 152294 -8992 152329 -8958
rect 152640 -8995 152675 -8961
rect 152685 -8995 152686 -8950
rect 152827 -9001 152828 -8697
rect 153519 -8706 153554 -8672
rect 153696 -8706 153731 -8672
rect 153992 -8723 154027 -8689
rect 154037 -8723 154038 -8681
rect 154179 -8753 154180 -8525
rect 154869 -8534 154904 -8500
rect 155046 -8534 155081 -8500
rect 155240 -8577 155275 -8543
rect 155285 -8577 155286 -8532
rect 155385 -8543 155386 -8532
rect 155594 -8537 155629 -8503
rect 155639 -8537 155640 -8492
rect 155739 -8503 155740 -8492
rect 155984 -8496 156019 -8462
rect 156029 -8496 156030 -8451
rect 156129 -8462 156130 -8451
rect 156140 -8496 156175 -8462
rect 156185 -8496 156186 -8451
rect 156285 -8462 156286 -8451
rect 156466 -8456 156501 -8422
rect 156538 -8456 156573 -8422
rect 156610 -8456 156645 -8422
rect 156754 -8456 156789 -8422
rect 156826 -8456 156861 -8422
rect 156863 -8456 156933 -8422
rect 156970 -8456 157005 -8422
rect 157040 -8456 157075 -8422
rect 156296 -8496 156331 -8462
rect 157336 -8491 157371 -8457
rect 157381 -8491 157382 -8446
rect 157481 -8457 157482 -8446
rect 157492 -8491 157527 -8457
rect 157537 -8491 157538 -8446
rect 157637 -8457 157638 -8446
rect 158213 -8451 158248 -8417
rect 158390 -8451 158425 -8417
rect 157648 -8491 157683 -8457
rect 155750 -8537 155785 -8503
rect 157029 -8505 157030 -8494
rect 155396 -8577 155431 -8543
rect 154309 -8621 154344 -8587
rect 154510 -8666 154545 -8632
rect 154633 -8637 154634 -8595
rect 154955 -8624 154990 -8590
rect 155594 -8620 155629 -8586
rect 155639 -8620 155640 -8575
rect 155739 -8586 155740 -8575
rect 155984 -8580 156019 -8546
rect 156029 -8580 156030 -8535
rect 156129 -8546 156130 -8535
rect 156140 -8580 156175 -8546
rect 156185 -8580 156186 -8535
rect 156285 -8546 156286 -8535
rect 156863 -8539 156898 -8505
rect 157040 -8539 157075 -8505
rect 156296 -8580 156331 -8546
rect 157183 -8565 157298 -8499
rect 157481 -8525 157482 -8499
rect 157878 -8517 157913 -8483
rect 157923 -8517 157924 -8472
rect 158023 -8483 158024 -8472
rect 158034 -8517 158069 -8483
rect 158079 -8517 158080 -8472
rect 158379 -8500 158380 -8489
rect 158584 -8494 158619 -8460
rect 158629 -8494 158630 -8449
rect 158729 -8460 158730 -8449
rect 158938 -8453 158973 -8419
rect 158983 -8453 158984 -8408
rect 159083 -8419 159084 -8408
rect 159264 -8413 159299 -8379
rect 159328 -8413 159371 -8379
rect 159373 -8413 159374 -8371
rect 159473 -8379 159474 -8371
rect 159408 -8413 159443 -8379
rect 159484 -8413 159519 -8379
rect 159529 -8413 159530 -8371
rect 159629 -8379 159630 -8371
rect 159578 -8413 159613 -8379
rect 159640 -8413 159685 -8379
rect 160680 -8408 160715 -8374
rect 160725 -8408 160726 -8363
rect 160825 -8374 160826 -8363
rect 160836 -8408 160871 -8374
rect 160881 -8408 160882 -8363
rect 160981 -8374 160982 -8363
rect 161557 -8367 161592 -8333
rect 161734 -8367 161769 -8333
rect 162327 -8336 162328 -8328
rect 162427 -8336 162428 -8328
rect 160992 -8408 161027 -8374
rect 159094 -8453 159129 -8419
rect 160373 -8422 160374 -8414
rect 161723 -8417 161724 -8406
rect 161928 -8410 161963 -8376
rect 161973 -8410 161974 -8365
rect 162073 -8376 162074 -8365
rect 162254 -8370 162317 -8336
rect 162326 -8370 162361 -8336
rect 162438 -8370 162473 -8336
rect 163163 -8360 163198 -8326
rect 163259 -8360 163294 -8326
rect 163355 -8360 163390 -8326
rect 163451 -8360 163486 -8326
rect 163547 -8360 163582 -8326
rect 163643 -8360 163678 -8326
rect 163739 -8360 163774 -8326
rect 165067 -8333 165068 -8322
rect 165244 -8327 165307 -8293
rect 165316 -8327 165351 -8293
rect 165428 -8327 165463 -8293
rect 165959 -8317 165994 -8283
rect 166055 -8317 166090 -8283
rect 166151 -8317 166186 -8283
rect 166247 -8317 166282 -8283
rect 166343 -8317 166378 -8283
rect 167368 -8324 167403 -8290
rect 167413 -8324 167414 -8279
rect 167513 -8290 167514 -8279
rect 167524 -8324 167559 -8290
rect 167569 -8324 167570 -8279
rect 167669 -8290 167670 -8279
rect 167848 -8284 167883 -8250
rect 167920 -8284 167955 -8250
rect 167992 -8284 168027 -8250
rect 168136 -8284 168171 -8250
rect 168208 -8284 168243 -8250
rect 168245 -8284 168315 -8250
rect 168352 -8284 168387 -8250
rect 168422 -8284 168457 -8250
rect 168949 -8274 168984 -8240
rect 169045 -8274 169080 -8240
rect 169141 -8274 169176 -8240
rect 170648 -8241 170683 -8207
rect 170712 -8241 170755 -8207
rect 170757 -8241 170758 -8199
rect 170857 -8207 170858 -8199
rect 170792 -8241 170827 -8207
rect 170868 -8241 170903 -8207
rect 170913 -8241 170914 -8199
rect 171013 -8207 171014 -8199
rect 170962 -8241 170997 -8207
rect 171024 -8241 171069 -8207
rect 171939 -8231 171974 -8197
rect 172035 -8231 172070 -8197
rect 172131 -8231 172166 -8197
rect 171755 -8250 171756 -8242
rect 167680 -8324 167715 -8290
rect 168661 -8293 168662 -8285
rect 168761 -8293 168762 -8285
rect 162084 -8410 162119 -8376
rect 158740 -8494 158775 -8460
rect 155750 -8620 155785 -8586
rect 157029 -8589 157030 -8578
rect 154279 -8689 154280 -8681
rect 154290 -8723 154325 -8689
rect 154510 -8734 154545 -8700
rect 152957 -8793 152992 -8759
rect 153160 -8838 153195 -8804
rect 153283 -8809 153284 -8767
rect 153605 -8796 153640 -8762
rect 152927 -8861 152928 -8853
rect 152938 -8895 152973 -8861
rect 153160 -8906 153195 -8872
rect 152927 -8961 152928 -8950
rect 152938 -8995 152973 -8961
rect 151875 -9045 151910 -9011
rect 151971 -9045 152006 -9011
rect 152067 -9045 152102 -9011
rect 152576 -9035 152611 -9001
rect 152648 -9035 152683 -9001
rect 152720 -9035 152755 -9001
rect 152792 -9029 152828 -9001
rect 153138 -9025 153173 -8991
rect 153183 -9025 153184 -8980
rect 152792 -9035 152827 -9029
rect 152229 -9088 152264 -9054
rect 152325 -9088 152360 -9054
rect 152421 -9088 152456 -9054
rect 153325 -9076 153326 -8809
rect 153954 -8819 154341 -8753
rect 153341 -8860 153376 -8826
rect 153690 -8832 153701 -8819
rect 153624 -8874 153701 -8832
rect 153752 -8874 154341 -8819
rect 154488 -8853 154523 -8819
rect 154533 -8853 154534 -8808
rect 153624 -8877 154341 -8874
rect 153341 -8928 153376 -8894
rect 153544 -8942 153579 -8908
rect 153589 -8942 153590 -8900
rect 153425 -8991 153426 -8980
rect 153436 -9025 153471 -8991
rect 153544 -9042 153579 -9008
rect 153589 -9042 153590 -8997
rect 153437 -9078 153472 -9044
rect 153509 -9078 153544 -9044
rect 153581 -9078 153616 -9044
rect 152583 -9131 152618 -9097
rect 152679 -9131 152714 -9097
rect 152775 -9131 152810 -9097
rect 152871 -9131 152906 -9097
rect 152967 -9131 153002 -9097
rect 153624 -9114 153769 -8877
rect 153954 -8899 154341 -8877
rect 153878 -8925 154341 -8899
rect 154675 -8904 154676 -8637
rect 154691 -8688 154726 -8654
rect 155305 -8691 155340 -8657
rect 155984 -8663 156019 -8629
rect 156029 -8663 156030 -8618
rect 156129 -8629 156130 -8618
rect 156140 -8663 156175 -8629
rect 156185 -8663 156186 -8618
rect 156285 -8629 156286 -8618
rect 156863 -8623 156898 -8589
rect 157040 -8623 157075 -8589
rect 157401 -8605 157436 -8571
rect 156296 -8663 156331 -8629
rect 156129 -8697 156130 -8671
rect 156528 -8689 156563 -8655
rect 156573 -8689 156574 -8644
rect 156673 -8655 156674 -8644
rect 156684 -8689 156719 -8655
rect 156729 -8689 156730 -8644
rect 157029 -8672 157030 -8661
rect 154691 -8756 154726 -8722
rect 154894 -8770 154929 -8736
rect 154939 -8770 154940 -8728
rect 155039 -8740 155040 -8729
rect 155659 -8734 155694 -8700
rect 155050 -8774 155085 -8740
rect 154775 -8819 154776 -8808
rect 155244 -8813 155279 -8779
rect 155289 -8813 155290 -8771
rect 155389 -8779 155390 -8771
rect 156049 -8777 156084 -8743
rect 155400 -8813 155435 -8779
rect 154786 -8853 154821 -8819
rect 154894 -8870 154929 -8836
rect 154939 -8870 154940 -8825
rect 155039 -8832 155040 -8821
rect 155050 -8866 155085 -8832
rect 155598 -8856 155633 -8822
rect 155643 -8856 155644 -8814
rect 155743 -8822 155744 -8814
rect 155754 -8856 155789 -8822
rect 154787 -8906 154822 -8872
rect 154859 -8906 154894 -8872
rect 154931 -8906 154966 -8872
rect 155244 -8913 155279 -8879
rect 155289 -8913 155290 -8868
rect 155389 -8879 155390 -8868
rect 155400 -8913 155435 -8879
rect 155984 -8895 156019 -8861
rect 156029 -8895 156030 -8853
rect 153878 -8959 154354 -8925
rect 155212 -8949 155247 -8915
rect 155284 -8949 155319 -8915
rect 155598 -8956 155633 -8922
rect 155643 -8956 155644 -8911
rect 155743 -8922 155744 -8911
rect 155754 -8956 155789 -8922
rect 153878 -8985 154341 -8959
rect 153882 -8993 154083 -8985
rect 153898 -9003 154067 -8993
rect 153624 -9140 153799 -9114
rect 153131 -9174 153166 -9140
rect 153227 -9174 153262 -9140
rect 153323 -9174 153358 -9140
rect 153419 -9174 153454 -9140
rect 153515 -9174 153550 -9140
rect 153611 -9174 153799 -9140
rect 153624 -9200 153799 -9174
rect 153824 -9174 153925 -9050
rect 153702 -9870 153737 -9200
rect 153824 -9228 153827 -9174
rect 153509 -9936 153654 -9924
rect 153177 -9970 153654 -9936
rect 153509 -9971 153654 -9970
rect 153690 -9971 153737 -9870
rect 153836 -9971 153871 -9174
rect 154094 -9971 154129 -9062
rect 154228 -9971 154263 -8985
rect 154481 -9002 154516 -8968
rect 154577 -9002 154612 -8968
rect 154673 -9002 154708 -8968
rect 154769 -9002 154804 -8968
rect 154865 -9002 154900 -8968
rect 154961 -9002 154996 -8968
rect 155057 -9002 155092 -8968
rect 155566 -8992 155601 -8958
rect 155638 -8992 155673 -8958
rect 155984 -8995 156019 -8961
rect 156029 -8995 156030 -8950
rect 156171 -9001 156172 -8697
rect 156863 -8706 156898 -8672
rect 157040 -8706 157075 -8672
rect 157336 -8723 157371 -8689
rect 157381 -8723 157382 -8681
rect 157523 -8753 157524 -8525
rect 158213 -8534 158248 -8500
rect 158390 -8534 158425 -8500
rect 158584 -8577 158619 -8543
rect 158629 -8577 158630 -8532
rect 158729 -8543 158730 -8532
rect 158938 -8537 158973 -8503
rect 158983 -8537 158984 -8492
rect 159083 -8503 159084 -8492
rect 159328 -8496 159363 -8462
rect 159373 -8496 159374 -8451
rect 159473 -8462 159474 -8451
rect 159484 -8496 159519 -8462
rect 159529 -8496 159530 -8451
rect 159629 -8462 159630 -8451
rect 159810 -8456 159845 -8422
rect 159882 -8456 159917 -8422
rect 159954 -8456 159989 -8422
rect 160098 -8456 160133 -8422
rect 160170 -8456 160205 -8422
rect 160207 -8456 160277 -8422
rect 160314 -8456 160349 -8422
rect 160384 -8456 160419 -8422
rect 159640 -8496 159675 -8462
rect 160680 -8491 160715 -8457
rect 160725 -8491 160726 -8446
rect 160825 -8457 160826 -8446
rect 160836 -8491 160871 -8457
rect 160881 -8491 160882 -8446
rect 160981 -8457 160982 -8446
rect 161557 -8451 161592 -8417
rect 161734 -8451 161769 -8417
rect 160992 -8491 161027 -8457
rect 159094 -8537 159129 -8503
rect 160373 -8505 160374 -8494
rect 158740 -8577 158775 -8543
rect 157653 -8621 157688 -8587
rect 157854 -8666 157889 -8632
rect 157977 -8637 157978 -8595
rect 158299 -8624 158334 -8590
rect 158938 -8620 158973 -8586
rect 158983 -8620 158984 -8575
rect 159083 -8586 159084 -8575
rect 159328 -8580 159363 -8546
rect 159373 -8580 159374 -8535
rect 159473 -8546 159474 -8535
rect 159484 -8580 159519 -8546
rect 159529 -8580 159530 -8535
rect 159629 -8546 159630 -8535
rect 160207 -8539 160242 -8505
rect 160384 -8539 160419 -8505
rect 159640 -8580 159675 -8546
rect 160527 -8565 160642 -8499
rect 160825 -8525 160826 -8499
rect 161222 -8517 161257 -8483
rect 161267 -8517 161268 -8472
rect 161367 -8483 161368 -8472
rect 161378 -8517 161413 -8483
rect 161423 -8517 161424 -8472
rect 161723 -8500 161724 -8489
rect 161928 -8494 161963 -8460
rect 161973 -8494 161974 -8449
rect 162073 -8460 162074 -8449
rect 162282 -8453 162317 -8419
rect 162327 -8453 162328 -8408
rect 162427 -8419 162428 -8408
rect 162608 -8413 162643 -8379
rect 162672 -8413 162715 -8379
rect 162717 -8413 162718 -8371
rect 162817 -8379 162818 -8371
rect 162752 -8413 162787 -8379
rect 162828 -8413 162863 -8379
rect 162873 -8413 162874 -8371
rect 162973 -8379 162974 -8371
rect 162922 -8413 162957 -8379
rect 162984 -8413 163029 -8379
rect 164024 -8408 164059 -8374
rect 164069 -8408 164070 -8363
rect 164169 -8374 164170 -8363
rect 164180 -8408 164215 -8374
rect 164225 -8408 164226 -8363
rect 164325 -8374 164326 -8363
rect 164901 -8367 164936 -8333
rect 165078 -8367 165113 -8333
rect 165671 -8336 165672 -8328
rect 165771 -8336 165772 -8328
rect 164336 -8408 164371 -8374
rect 162438 -8453 162473 -8419
rect 163717 -8422 163718 -8414
rect 165067 -8417 165068 -8406
rect 165272 -8410 165307 -8376
rect 165317 -8410 165318 -8365
rect 165417 -8376 165418 -8365
rect 165598 -8370 165661 -8336
rect 165670 -8370 165705 -8336
rect 165782 -8370 165817 -8336
rect 166507 -8360 166542 -8326
rect 166603 -8360 166638 -8326
rect 166699 -8360 166734 -8326
rect 166795 -8360 166830 -8326
rect 166891 -8360 166926 -8326
rect 166987 -8360 167022 -8326
rect 167083 -8360 167118 -8326
rect 168411 -8333 168412 -8322
rect 168588 -8327 168651 -8293
rect 168660 -8327 168695 -8293
rect 168772 -8327 168807 -8293
rect 169303 -8317 169338 -8283
rect 169399 -8317 169434 -8283
rect 169495 -8317 169530 -8283
rect 169591 -8317 169626 -8283
rect 169687 -8317 169722 -8283
rect 170712 -8324 170747 -8290
rect 170757 -8324 170758 -8279
rect 170857 -8290 170858 -8279
rect 170868 -8324 170903 -8290
rect 170913 -8324 170914 -8279
rect 171013 -8290 171014 -8279
rect 171192 -8284 171227 -8250
rect 171264 -8284 171299 -8250
rect 171336 -8284 171371 -8250
rect 171480 -8284 171515 -8250
rect 171552 -8284 171587 -8250
rect 171589 -8284 171659 -8250
rect 171696 -8284 171731 -8250
rect 171766 -8284 171801 -8250
rect 172293 -8274 172328 -8240
rect 172389 -8274 172424 -8240
rect 172485 -8274 172520 -8240
rect 173992 -8241 174027 -8207
rect 174056 -8241 174099 -8207
rect 174101 -8241 174102 -8199
rect 174201 -8207 174202 -8199
rect 174136 -8241 174171 -8207
rect 174212 -8241 174247 -8207
rect 174257 -8241 174258 -8199
rect 174357 -8207 174358 -8199
rect 174306 -8241 174341 -8207
rect 174368 -8241 174413 -8207
rect 175283 -8231 175318 -8197
rect 175379 -8231 175414 -8197
rect 175475 -8231 175510 -8197
rect 175099 -8250 175100 -8242
rect 171024 -8324 171059 -8290
rect 172005 -8293 172006 -8285
rect 172105 -8293 172106 -8285
rect 165428 -8410 165463 -8376
rect 162084 -8494 162119 -8460
rect 159094 -8620 159129 -8586
rect 160373 -8589 160374 -8578
rect 157623 -8689 157624 -8681
rect 157634 -8723 157669 -8689
rect 157854 -8734 157889 -8700
rect 156301 -8793 156336 -8759
rect 156504 -8838 156539 -8804
rect 156627 -8809 156628 -8767
rect 156949 -8796 156984 -8762
rect 156271 -8861 156272 -8853
rect 156282 -8895 156317 -8861
rect 156504 -8906 156539 -8872
rect 156271 -8961 156272 -8950
rect 156282 -8995 156317 -8961
rect 155219 -9045 155254 -9011
rect 155315 -9045 155350 -9011
rect 155411 -9045 155446 -9011
rect 155920 -9035 155955 -9001
rect 155992 -9035 156027 -9001
rect 156064 -9035 156099 -9001
rect 156136 -9029 156172 -9001
rect 156482 -9025 156517 -8991
rect 156527 -9025 156528 -8980
rect 156136 -9035 156171 -9029
rect 155573 -9088 155608 -9054
rect 155669 -9088 155704 -9054
rect 155765 -9088 155800 -9054
rect 156669 -9076 156670 -8809
rect 157298 -8819 157685 -8753
rect 156685 -8860 156720 -8826
rect 157034 -8832 157045 -8819
rect 156968 -8874 157045 -8832
rect 157096 -8874 157685 -8819
rect 157832 -8853 157867 -8819
rect 157877 -8853 157878 -8808
rect 156968 -8877 157685 -8874
rect 156685 -8928 156720 -8894
rect 156888 -8942 156923 -8908
rect 156933 -8942 156934 -8900
rect 156769 -8991 156770 -8980
rect 156780 -9025 156815 -8991
rect 156888 -9042 156923 -9008
rect 156933 -9042 156934 -8997
rect 156781 -9078 156816 -9044
rect 156853 -9078 156888 -9044
rect 156925 -9078 156960 -9044
rect 155927 -9131 155962 -9097
rect 156023 -9131 156058 -9097
rect 156119 -9131 156154 -9097
rect 156215 -9131 156250 -9097
rect 156311 -9131 156346 -9097
rect 156968 -9114 157113 -8877
rect 157298 -8899 157685 -8877
rect 157222 -8925 157685 -8899
rect 158019 -8904 158020 -8637
rect 158035 -8688 158070 -8654
rect 158649 -8691 158684 -8657
rect 159328 -8663 159363 -8629
rect 159373 -8663 159374 -8618
rect 159473 -8629 159474 -8618
rect 159484 -8663 159519 -8629
rect 159529 -8663 159530 -8618
rect 159629 -8629 159630 -8618
rect 160207 -8623 160242 -8589
rect 160384 -8623 160419 -8589
rect 160745 -8605 160780 -8571
rect 159640 -8663 159675 -8629
rect 159473 -8697 159474 -8671
rect 159872 -8689 159907 -8655
rect 159917 -8689 159918 -8644
rect 160017 -8655 160018 -8644
rect 160028 -8689 160063 -8655
rect 160073 -8689 160074 -8644
rect 160373 -8672 160374 -8661
rect 158035 -8756 158070 -8722
rect 158238 -8770 158273 -8736
rect 158283 -8770 158284 -8728
rect 158383 -8740 158384 -8729
rect 159003 -8734 159038 -8700
rect 158394 -8774 158429 -8740
rect 158119 -8819 158120 -8808
rect 158588 -8813 158623 -8779
rect 158633 -8813 158634 -8771
rect 158733 -8779 158734 -8771
rect 159393 -8777 159428 -8743
rect 158744 -8813 158779 -8779
rect 158130 -8853 158165 -8819
rect 158238 -8870 158273 -8836
rect 158283 -8870 158284 -8825
rect 158383 -8832 158384 -8821
rect 158394 -8866 158429 -8832
rect 158942 -8856 158977 -8822
rect 158987 -8856 158988 -8814
rect 159087 -8822 159088 -8814
rect 159098 -8856 159133 -8822
rect 158131 -8906 158166 -8872
rect 158203 -8906 158238 -8872
rect 158275 -8906 158310 -8872
rect 158588 -8913 158623 -8879
rect 158633 -8913 158634 -8868
rect 158733 -8879 158734 -8868
rect 158744 -8913 158779 -8879
rect 159328 -8895 159363 -8861
rect 159373 -8895 159374 -8853
rect 157222 -8959 157698 -8925
rect 158556 -8949 158591 -8915
rect 158628 -8949 158663 -8915
rect 158942 -8956 158977 -8922
rect 158987 -8956 158988 -8911
rect 159087 -8922 159088 -8911
rect 159098 -8956 159133 -8922
rect 157222 -8985 157685 -8959
rect 157226 -8993 157427 -8985
rect 157242 -9003 157411 -8993
rect 156968 -9140 157143 -9114
rect 156475 -9174 156510 -9140
rect 156571 -9174 156606 -9140
rect 156667 -9174 156702 -9140
rect 156763 -9174 156798 -9140
rect 156859 -9174 156894 -9140
rect 156955 -9174 157143 -9140
rect 156968 -9200 157143 -9174
rect 157168 -9174 157269 -9050
rect 157046 -9870 157081 -9200
rect 157168 -9228 157171 -9174
rect 156853 -9936 156998 -9924
rect 156521 -9970 156998 -9936
rect 156853 -9971 156998 -9970
rect 157034 -9971 157081 -9870
rect 157180 -9971 157215 -9174
rect 157438 -9971 157473 -9062
rect 157572 -9971 157607 -8985
rect 157825 -9002 157860 -8968
rect 157921 -9002 157956 -8968
rect 158017 -9002 158052 -8968
rect 158113 -9002 158148 -8968
rect 158209 -9002 158244 -8968
rect 158305 -9002 158340 -8968
rect 158401 -9002 158436 -8968
rect 158910 -8992 158945 -8958
rect 158982 -8992 159017 -8958
rect 159328 -8995 159363 -8961
rect 159373 -8995 159374 -8950
rect 159515 -9001 159516 -8697
rect 160207 -8706 160242 -8672
rect 160384 -8706 160419 -8672
rect 160680 -8723 160715 -8689
rect 160725 -8723 160726 -8681
rect 160867 -8753 160868 -8525
rect 161557 -8534 161592 -8500
rect 161734 -8534 161769 -8500
rect 161928 -8577 161963 -8543
rect 161973 -8577 161974 -8532
rect 162073 -8543 162074 -8532
rect 162282 -8537 162317 -8503
rect 162327 -8537 162328 -8492
rect 162427 -8503 162428 -8492
rect 162672 -8496 162707 -8462
rect 162717 -8496 162718 -8451
rect 162817 -8462 162818 -8451
rect 162828 -8496 162863 -8462
rect 162873 -8496 162874 -8451
rect 162973 -8462 162974 -8451
rect 163154 -8456 163189 -8422
rect 163226 -8456 163261 -8422
rect 163298 -8456 163333 -8422
rect 163442 -8456 163477 -8422
rect 163514 -8456 163549 -8422
rect 163551 -8456 163621 -8422
rect 163658 -8456 163693 -8422
rect 163728 -8456 163763 -8422
rect 162984 -8496 163019 -8462
rect 164024 -8491 164059 -8457
rect 164069 -8491 164070 -8446
rect 164169 -8457 164170 -8446
rect 164180 -8491 164215 -8457
rect 164225 -8491 164226 -8446
rect 164325 -8457 164326 -8446
rect 164901 -8451 164936 -8417
rect 165078 -8451 165113 -8417
rect 164336 -8491 164371 -8457
rect 162438 -8537 162473 -8503
rect 163717 -8505 163718 -8494
rect 162084 -8577 162119 -8543
rect 160997 -8621 161032 -8587
rect 161198 -8666 161233 -8632
rect 161321 -8637 161322 -8595
rect 161643 -8624 161678 -8590
rect 162282 -8620 162317 -8586
rect 162327 -8620 162328 -8575
rect 162427 -8586 162428 -8575
rect 162672 -8580 162707 -8546
rect 162717 -8580 162718 -8535
rect 162817 -8546 162818 -8535
rect 162828 -8580 162863 -8546
rect 162873 -8580 162874 -8535
rect 162973 -8546 162974 -8535
rect 163551 -8539 163586 -8505
rect 163728 -8539 163763 -8505
rect 162984 -8580 163019 -8546
rect 163871 -8565 163986 -8499
rect 164169 -8525 164170 -8499
rect 164566 -8517 164601 -8483
rect 164611 -8517 164612 -8472
rect 164711 -8483 164712 -8472
rect 164722 -8517 164757 -8483
rect 164767 -8517 164768 -8472
rect 165067 -8500 165068 -8489
rect 165272 -8494 165307 -8460
rect 165317 -8494 165318 -8449
rect 165417 -8460 165418 -8449
rect 165626 -8453 165661 -8419
rect 165671 -8453 165672 -8408
rect 165771 -8419 165772 -8408
rect 165952 -8413 165987 -8379
rect 166016 -8413 166059 -8379
rect 166061 -8413 166062 -8371
rect 166161 -8379 166162 -8371
rect 166096 -8413 166131 -8379
rect 166172 -8413 166207 -8379
rect 166217 -8413 166218 -8371
rect 166317 -8379 166318 -8371
rect 166266 -8413 166301 -8379
rect 166328 -8413 166373 -8379
rect 167368 -8408 167403 -8374
rect 167413 -8408 167414 -8363
rect 167513 -8374 167514 -8363
rect 167524 -8408 167559 -8374
rect 167569 -8408 167570 -8363
rect 167669 -8374 167670 -8363
rect 168245 -8367 168280 -8333
rect 168422 -8367 168457 -8333
rect 169015 -8336 169016 -8328
rect 169115 -8336 169116 -8328
rect 167680 -8408 167715 -8374
rect 165782 -8453 165817 -8419
rect 167061 -8422 167062 -8414
rect 168411 -8417 168412 -8406
rect 168616 -8410 168651 -8376
rect 168661 -8410 168662 -8365
rect 168761 -8376 168762 -8365
rect 168942 -8370 169005 -8336
rect 169014 -8370 169049 -8336
rect 169126 -8370 169161 -8336
rect 169851 -8360 169886 -8326
rect 169947 -8360 169982 -8326
rect 170043 -8360 170078 -8326
rect 170139 -8360 170174 -8326
rect 170235 -8360 170270 -8326
rect 170331 -8360 170366 -8326
rect 170427 -8360 170462 -8326
rect 171755 -8333 171756 -8322
rect 171932 -8327 171995 -8293
rect 172004 -8327 172039 -8293
rect 172116 -8327 172151 -8293
rect 172647 -8317 172682 -8283
rect 172743 -8317 172778 -8283
rect 172839 -8317 172874 -8283
rect 172935 -8317 172970 -8283
rect 173031 -8317 173066 -8283
rect 174056 -8324 174091 -8290
rect 174101 -8324 174102 -8279
rect 174201 -8290 174202 -8279
rect 174212 -8324 174247 -8290
rect 174257 -8324 174258 -8279
rect 174357 -8290 174358 -8279
rect 174536 -8284 174571 -8250
rect 174608 -8284 174643 -8250
rect 174680 -8284 174715 -8250
rect 174824 -8284 174859 -8250
rect 174896 -8284 174931 -8250
rect 174933 -8284 175003 -8250
rect 175040 -8284 175075 -8250
rect 175110 -8284 175145 -8250
rect 175637 -8274 175672 -8240
rect 175733 -8274 175768 -8240
rect 175829 -8274 175864 -8240
rect 177336 -8241 177371 -8207
rect 177400 -8241 177443 -8207
rect 177445 -8241 177446 -8199
rect 177545 -8207 177546 -8199
rect 177480 -8241 177515 -8207
rect 177556 -8241 177591 -8207
rect 177601 -8241 177602 -8199
rect 177701 -8207 177702 -8199
rect 177650 -8241 177685 -8207
rect 177712 -8241 177757 -8207
rect 178627 -8231 178662 -8197
rect 178723 -8231 178758 -8197
rect 178819 -8231 178854 -8197
rect 178443 -8250 178444 -8242
rect 174368 -8324 174403 -8290
rect 175349 -8293 175350 -8285
rect 175449 -8293 175450 -8285
rect 168772 -8410 168807 -8376
rect 165428 -8494 165463 -8460
rect 162438 -8620 162473 -8586
rect 163717 -8589 163718 -8578
rect 160967 -8689 160968 -8681
rect 160978 -8723 161013 -8689
rect 161198 -8734 161233 -8700
rect 159645 -8793 159680 -8759
rect 159848 -8838 159883 -8804
rect 159971 -8809 159972 -8767
rect 160293 -8796 160328 -8762
rect 159615 -8861 159616 -8853
rect 159626 -8895 159661 -8861
rect 159848 -8906 159883 -8872
rect 159615 -8961 159616 -8950
rect 159626 -8995 159661 -8961
rect 158563 -9045 158598 -9011
rect 158659 -9045 158694 -9011
rect 158755 -9045 158790 -9011
rect 159264 -9035 159299 -9001
rect 159336 -9035 159371 -9001
rect 159408 -9035 159443 -9001
rect 159480 -9029 159516 -9001
rect 159826 -9025 159861 -8991
rect 159871 -9025 159872 -8980
rect 159480 -9035 159515 -9029
rect 158917 -9088 158952 -9054
rect 159013 -9088 159048 -9054
rect 159109 -9088 159144 -9054
rect 160013 -9076 160014 -8809
rect 160642 -8819 161029 -8753
rect 160029 -8860 160064 -8826
rect 160378 -8832 160389 -8819
rect 160312 -8874 160389 -8832
rect 160440 -8874 161029 -8819
rect 161176 -8853 161211 -8819
rect 161221 -8853 161222 -8808
rect 160312 -8877 161029 -8874
rect 160029 -8928 160064 -8894
rect 160232 -8942 160267 -8908
rect 160277 -8942 160278 -8900
rect 160113 -8991 160114 -8980
rect 160124 -9025 160159 -8991
rect 160232 -9042 160267 -9008
rect 160277 -9042 160278 -8997
rect 160125 -9078 160160 -9044
rect 160197 -9078 160232 -9044
rect 160269 -9078 160304 -9044
rect 159271 -9131 159306 -9097
rect 159367 -9131 159402 -9097
rect 159463 -9131 159498 -9097
rect 159559 -9131 159594 -9097
rect 159655 -9131 159690 -9097
rect 160312 -9114 160457 -8877
rect 160642 -8899 161029 -8877
rect 160566 -8925 161029 -8899
rect 161363 -8904 161364 -8637
rect 161379 -8688 161414 -8654
rect 161993 -8691 162028 -8657
rect 162672 -8663 162707 -8629
rect 162717 -8663 162718 -8618
rect 162817 -8629 162818 -8618
rect 162828 -8663 162863 -8629
rect 162873 -8663 162874 -8618
rect 162973 -8629 162974 -8618
rect 163551 -8623 163586 -8589
rect 163728 -8623 163763 -8589
rect 164089 -8605 164124 -8571
rect 162984 -8663 163019 -8629
rect 162817 -8697 162818 -8671
rect 163216 -8689 163251 -8655
rect 163261 -8689 163262 -8644
rect 163361 -8655 163362 -8644
rect 163372 -8689 163407 -8655
rect 163417 -8689 163418 -8644
rect 163717 -8672 163718 -8661
rect 161379 -8756 161414 -8722
rect 161582 -8770 161617 -8736
rect 161627 -8770 161628 -8728
rect 161727 -8740 161728 -8729
rect 162347 -8734 162382 -8700
rect 161738 -8774 161773 -8740
rect 161463 -8819 161464 -8808
rect 161932 -8813 161967 -8779
rect 161977 -8813 161978 -8771
rect 162077 -8779 162078 -8771
rect 162737 -8777 162772 -8743
rect 162088 -8813 162123 -8779
rect 161474 -8853 161509 -8819
rect 161582 -8870 161617 -8836
rect 161627 -8870 161628 -8825
rect 161727 -8832 161728 -8821
rect 161738 -8866 161773 -8832
rect 162286 -8856 162321 -8822
rect 162331 -8856 162332 -8814
rect 162431 -8822 162432 -8814
rect 162442 -8856 162477 -8822
rect 161475 -8906 161510 -8872
rect 161547 -8906 161582 -8872
rect 161619 -8906 161654 -8872
rect 161932 -8913 161967 -8879
rect 161977 -8913 161978 -8868
rect 162077 -8879 162078 -8868
rect 162088 -8913 162123 -8879
rect 162672 -8895 162707 -8861
rect 162717 -8895 162718 -8853
rect 160566 -8959 161042 -8925
rect 161900 -8949 161935 -8915
rect 161972 -8949 162007 -8915
rect 162286 -8956 162321 -8922
rect 162331 -8956 162332 -8911
rect 162431 -8922 162432 -8911
rect 162442 -8956 162477 -8922
rect 160566 -8985 161029 -8959
rect 160570 -8993 160771 -8985
rect 160586 -9003 160755 -8993
rect 160312 -9140 160487 -9114
rect 159819 -9174 159854 -9140
rect 159915 -9174 159950 -9140
rect 160011 -9174 160046 -9140
rect 160107 -9174 160142 -9140
rect 160203 -9174 160238 -9140
rect 160299 -9174 160487 -9140
rect 160312 -9200 160487 -9174
rect 160512 -9174 160613 -9050
rect 160390 -9870 160425 -9200
rect 160512 -9228 160515 -9174
rect 160197 -9936 160342 -9924
rect 159865 -9970 160342 -9936
rect 160197 -9971 160342 -9970
rect 160378 -9971 160425 -9870
rect 160524 -9971 160559 -9174
rect 160782 -9971 160817 -9062
rect 160916 -9971 160951 -8985
rect 161169 -9002 161204 -8968
rect 161265 -9002 161300 -8968
rect 161361 -9002 161396 -8968
rect 161457 -9002 161492 -8968
rect 161553 -9002 161588 -8968
rect 161649 -9002 161684 -8968
rect 161745 -9002 161780 -8968
rect 162254 -8992 162289 -8958
rect 162326 -8992 162361 -8958
rect 162672 -8995 162707 -8961
rect 162717 -8995 162718 -8950
rect 162859 -9001 162860 -8697
rect 163551 -8706 163586 -8672
rect 163728 -8706 163763 -8672
rect 164024 -8723 164059 -8689
rect 164069 -8723 164070 -8681
rect 164211 -8753 164212 -8525
rect 164901 -8534 164936 -8500
rect 165078 -8534 165113 -8500
rect 165272 -8577 165307 -8543
rect 165317 -8577 165318 -8532
rect 165417 -8543 165418 -8532
rect 165626 -8537 165661 -8503
rect 165671 -8537 165672 -8492
rect 165771 -8503 165772 -8492
rect 166016 -8496 166051 -8462
rect 166061 -8496 166062 -8451
rect 166161 -8462 166162 -8451
rect 166172 -8496 166207 -8462
rect 166217 -8496 166218 -8451
rect 166317 -8462 166318 -8451
rect 166498 -8456 166533 -8422
rect 166570 -8456 166605 -8422
rect 166642 -8456 166677 -8422
rect 166786 -8456 166821 -8422
rect 166858 -8456 166893 -8422
rect 166895 -8456 166965 -8422
rect 167002 -8456 167037 -8422
rect 167072 -8456 167107 -8422
rect 166328 -8496 166363 -8462
rect 167368 -8491 167403 -8457
rect 167413 -8491 167414 -8446
rect 167513 -8457 167514 -8446
rect 167524 -8491 167559 -8457
rect 167569 -8491 167570 -8446
rect 167669 -8457 167670 -8446
rect 168245 -8451 168280 -8417
rect 168422 -8451 168457 -8417
rect 167680 -8491 167715 -8457
rect 165782 -8537 165817 -8503
rect 167061 -8505 167062 -8494
rect 165428 -8577 165463 -8543
rect 164341 -8621 164376 -8587
rect 164542 -8666 164577 -8632
rect 164665 -8637 164666 -8595
rect 164987 -8624 165022 -8590
rect 165626 -8620 165661 -8586
rect 165671 -8620 165672 -8575
rect 165771 -8586 165772 -8575
rect 166016 -8580 166051 -8546
rect 166061 -8580 166062 -8535
rect 166161 -8546 166162 -8535
rect 166172 -8580 166207 -8546
rect 166217 -8580 166218 -8535
rect 166317 -8546 166318 -8535
rect 166895 -8539 166930 -8505
rect 167072 -8539 167107 -8505
rect 166328 -8580 166363 -8546
rect 167215 -8565 167330 -8499
rect 167513 -8525 167514 -8499
rect 167910 -8517 167945 -8483
rect 167955 -8517 167956 -8472
rect 168055 -8483 168056 -8472
rect 168066 -8517 168101 -8483
rect 168111 -8517 168112 -8472
rect 168411 -8500 168412 -8489
rect 168616 -8494 168651 -8460
rect 168661 -8494 168662 -8449
rect 168761 -8460 168762 -8449
rect 168970 -8453 169005 -8419
rect 169015 -8453 169016 -8408
rect 169115 -8419 169116 -8408
rect 169296 -8413 169331 -8379
rect 169360 -8413 169403 -8379
rect 169405 -8413 169406 -8371
rect 169505 -8379 169506 -8371
rect 169440 -8413 169475 -8379
rect 169516 -8413 169551 -8379
rect 169561 -8413 169562 -8371
rect 169661 -8379 169662 -8371
rect 169610 -8413 169645 -8379
rect 169672 -8413 169717 -8379
rect 170712 -8408 170747 -8374
rect 170757 -8408 170758 -8363
rect 170857 -8374 170858 -8363
rect 170868 -8408 170903 -8374
rect 170913 -8408 170914 -8363
rect 171013 -8374 171014 -8363
rect 171589 -8367 171624 -8333
rect 171766 -8367 171801 -8333
rect 172359 -8336 172360 -8328
rect 172459 -8336 172460 -8328
rect 171024 -8408 171059 -8374
rect 169126 -8453 169161 -8419
rect 170405 -8422 170406 -8414
rect 171755 -8417 171756 -8406
rect 171960 -8410 171995 -8376
rect 172005 -8410 172006 -8365
rect 172105 -8376 172106 -8365
rect 172286 -8370 172349 -8336
rect 172358 -8370 172393 -8336
rect 172470 -8370 172505 -8336
rect 173195 -8360 173230 -8326
rect 173291 -8360 173326 -8326
rect 173387 -8360 173422 -8326
rect 173483 -8360 173518 -8326
rect 173579 -8360 173614 -8326
rect 173675 -8360 173710 -8326
rect 173771 -8360 173806 -8326
rect 175099 -8333 175100 -8322
rect 175276 -8327 175339 -8293
rect 175348 -8327 175383 -8293
rect 175460 -8327 175495 -8293
rect 175991 -8317 176026 -8283
rect 176087 -8317 176122 -8283
rect 176183 -8317 176218 -8283
rect 176279 -8317 176314 -8283
rect 176375 -8317 176410 -8283
rect 177400 -8324 177435 -8290
rect 177445 -8324 177446 -8279
rect 177545 -8290 177546 -8279
rect 177556 -8324 177591 -8290
rect 177601 -8324 177602 -8279
rect 177701 -8290 177702 -8279
rect 177880 -8284 177915 -8250
rect 177952 -8284 177987 -8250
rect 178024 -8284 178059 -8250
rect 178168 -8284 178203 -8250
rect 178240 -8284 178275 -8250
rect 178277 -8284 178347 -8250
rect 178384 -8284 178419 -8250
rect 178454 -8284 178489 -8250
rect 178981 -8274 179016 -8240
rect 179077 -8274 179112 -8240
rect 179173 -8274 179208 -8240
rect 180680 -8241 180715 -8207
rect 180744 -8241 180787 -8207
rect 180789 -8241 180790 -8199
rect 180889 -8207 180890 -8199
rect 180824 -8241 180859 -8207
rect 180900 -8241 180935 -8207
rect 180945 -8241 180946 -8199
rect 181045 -8207 181046 -8199
rect 180994 -8241 181029 -8207
rect 181056 -8241 181101 -8207
rect 181971 -8231 182006 -8197
rect 182067 -8231 182102 -8197
rect 182163 -8231 182198 -8197
rect 181787 -8250 181788 -8242
rect 177712 -8324 177747 -8290
rect 178693 -8293 178694 -8285
rect 178793 -8293 178794 -8285
rect 172116 -8410 172151 -8376
rect 168772 -8494 168807 -8460
rect 165782 -8620 165817 -8586
rect 167061 -8589 167062 -8578
rect 164311 -8689 164312 -8681
rect 164322 -8723 164357 -8689
rect 164542 -8734 164577 -8700
rect 162989 -8793 163024 -8759
rect 163192 -8838 163227 -8804
rect 163315 -8809 163316 -8767
rect 163637 -8796 163672 -8762
rect 162959 -8861 162960 -8853
rect 162970 -8895 163005 -8861
rect 163192 -8906 163227 -8872
rect 162959 -8961 162960 -8950
rect 162970 -8995 163005 -8961
rect 161907 -9045 161942 -9011
rect 162003 -9045 162038 -9011
rect 162099 -9045 162134 -9011
rect 162608 -9035 162643 -9001
rect 162680 -9035 162715 -9001
rect 162752 -9035 162787 -9001
rect 162824 -9029 162860 -9001
rect 163170 -9025 163205 -8991
rect 163215 -9025 163216 -8980
rect 162824 -9035 162859 -9029
rect 162261 -9088 162296 -9054
rect 162357 -9088 162392 -9054
rect 162453 -9088 162488 -9054
rect 163357 -9076 163358 -8809
rect 163986 -8819 164373 -8753
rect 163373 -8860 163408 -8826
rect 163722 -8832 163733 -8819
rect 163656 -8874 163733 -8832
rect 163784 -8874 164373 -8819
rect 164520 -8853 164555 -8819
rect 164565 -8853 164566 -8808
rect 163656 -8877 164373 -8874
rect 163373 -8928 163408 -8894
rect 163576 -8942 163611 -8908
rect 163621 -8942 163622 -8900
rect 163457 -8991 163458 -8980
rect 163468 -9025 163503 -8991
rect 163576 -9042 163611 -9008
rect 163621 -9042 163622 -8997
rect 163469 -9078 163504 -9044
rect 163541 -9078 163576 -9044
rect 163613 -9078 163648 -9044
rect 162615 -9131 162650 -9097
rect 162711 -9131 162746 -9097
rect 162807 -9131 162842 -9097
rect 162903 -9131 162938 -9097
rect 162999 -9131 163034 -9097
rect 163656 -9114 163801 -8877
rect 163986 -8899 164373 -8877
rect 163910 -8925 164373 -8899
rect 164707 -8904 164708 -8637
rect 164723 -8688 164758 -8654
rect 165337 -8691 165372 -8657
rect 166016 -8663 166051 -8629
rect 166061 -8663 166062 -8618
rect 166161 -8629 166162 -8618
rect 166172 -8663 166207 -8629
rect 166217 -8663 166218 -8618
rect 166317 -8629 166318 -8618
rect 166895 -8623 166930 -8589
rect 167072 -8623 167107 -8589
rect 167433 -8605 167468 -8571
rect 166328 -8663 166363 -8629
rect 166161 -8697 166162 -8671
rect 166560 -8689 166595 -8655
rect 166605 -8689 166606 -8644
rect 166705 -8655 166706 -8644
rect 166716 -8689 166751 -8655
rect 166761 -8689 166762 -8644
rect 167061 -8672 167062 -8661
rect 164723 -8756 164758 -8722
rect 164926 -8770 164961 -8736
rect 164971 -8770 164972 -8728
rect 165071 -8740 165072 -8729
rect 165691 -8734 165726 -8700
rect 165082 -8774 165117 -8740
rect 164807 -8819 164808 -8808
rect 165276 -8813 165311 -8779
rect 165321 -8813 165322 -8771
rect 165421 -8779 165422 -8771
rect 166081 -8777 166116 -8743
rect 165432 -8813 165467 -8779
rect 164818 -8853 164853 -8819
rect 164926 -8870 164961 -8836
rect 164971 -8870 164972 -8825
rect 165071 -8832 165072 -8821
rect 165082 -8866 165117 -8832
rect 165630 -8856 165665 -8822
rect 165675 -8856 165676 -8814
rect 165775 -8822 165776 -8814
rect 165786 -8856 165821 -8822
rect 164819 -8906 164854 -8872
rect 164891 -8906 164926 -8872
rect 164963 -8906 164998 -8872
rect 165276 -8913 165311 -8879
rect 165321 -8913 165322 -8868
rect 165421 -8879 165422 -8868
rect 165432 -8913 165467 -8879
rect 166016 -8895 166051 -8861
rect 166061 -8895 166062 -8853
rect 163910 -8959 164386 -8925
rect 165244 -8949 165279 -8915
rect 165316 -8949 165351 -8915
rect 165630 -8956 165665 -8922
rect 165675 -8956 165676 -8911
rect 165775 -8922 165776 -8911
rect 165786 -8956 165821 -8922
rect 163910 -8985 164373 -8959
rect 163914 -8993 164115 -8985
rect 163930 -9003 164099 -8993
rect 163656 -9140 163831 -9114
rect 163163 -9174 163198 -9140
rect 163259 -9174 163294 -9140
rect 163355 -9174 163390 -9140
rect 163451 -9174 163486 -9140
rect 163547 -9174 163582 -9140
rect 163643 -9174 163831 -9140
rect 163656 -9200 163831 -9174
rect 163856 -9174 163957 -9050
rect 163734 -9870 163769 -9200
rect 163856 -9228 163859 -9174
rect 163541 -9936 163686 -9924
rect 163209 -9970 163686 -9936
rect 163541 -9971 163686 -9970
rect 163722 -9971 163769 -9870
rect 163868 -9971 163903 -9174
rect 164126 -9971 164161 -9062
rect 164260 -9971 164295 -8985
rect 164513 -9002 164548 -8968
rect 164609 -9002 164644 -8968
rect 164705 -9002 164740 -8968
rect 164801 -9002 164836 -8968
rect 164897 -9002 164932 -8968
rect 164993 -9002 165028 -8968
rect 165089 -9002 165124 -8968
rect 165598 -8992 165633 -8958
rect 165670 -8992 165705 -8958
rect 166016 -8995 166051 -8961
rect 166061 -8995 166062 -8950
rect 166203 -9001 166204 -8697
rect 166895 -8706 166930 -8672
rect 167072 -8706 167107 -8672
rect 167368 -8723 167403 -8689
rect 167413 -8723 167414 -8681
rect 167555 -8753 167556 -8525
rect 168245 -8534 168280 -8500
rect 168422 -8534 168457 -8500
rect 168616 -8577 168651 -8543
rect 168661 -8577 168662 -8532
rect 168761 -8543 168762 -8532
rect 168970 -8537 169005 -8503
rect 169015 -8537 169016 -8492
rect 169115 -8503 169116 -8492
rect 169360 -8496 169395 -8462
rect 169405 -8496 169406 -8451
rect 169505 -8462 169506 -8451
rect 169516 -8496 169551 -8462
rect 169561 -8496 169562 -8451
rect 169661 -8462 169662 -8451
rect 169842 -8456 169877 -8422
rect 169914 -8456 169949 -8422
rect 169986 -8456 170021 -8422
rect 170130 -8456 170165 -8422
rect 170202 -8456 170237 -8422
rect 170239 -8456 170309 -8422
rect 170346 -8456 170381 -8422
rect 170416 -8456 170451 -8422
rect 169672 -8496 169707 -8462
rect 170712 -8491 170747 -8457
rect 170757 -8491 170758 -8446
rect 170857 -8457 170858 -8446
rect 170868 -8491 170903 -8457
rect 170913 -8491 170914 -8446
rect 171013 -8457 171014 -8446
rect 171589 -8451 171624 -8417
rect 171766 -8451 171801 -8417
rect 171024 -8491 171059 -8457
rect 169126 -8537 169161 -8503
rect 170405 -8505 170406 -8494
rect 168772 -8577 168807 -8543
rect 167685 -8621 167720 -8587
rect 167886 -8666 167921 -8632
rect 168009 -8637 168010 -8595
rect 168331 -8624 168366 -8590
rect 168970 -8620 169005 -8586
rect 169015 -8620 169016 -8575
rect 169115 -8586 169116 -8575
rect 169360 -8580 169395 -8546
rect 169405 -8580 169406 -8535
rect 169505 -8546 169506 -8535
rect 169516 -8580 169551 -8546
rect 169561 -8580 169562 -8535
rect 169661 -8546 169662 -8535
rect 170239 -8539 170274 -8505
rect 170416 -8539 170451 -8505
rect 169672 -8580 169707 -8546
rect 170559 -8565 170674 -8499
rect 170857 -8525 170858 -8499
rect 171254 -8517 171289 -8483
rect 171299 -8517 171300 -8472
rect 171399 -8483 171400 -8472
rect 171410 -8517 171445 -8483
rect 171455 -8517 171456 -8472
rect 171755 -8500 171756 -8489
rect 171960 -8494 171995 -8460
rect 172005 -8494 172006 -8449
rect 172105 -8460 172106 -8449
rect 172314 -8453 172349 -8419
rect 172359 -8453 172360 -8408
rect 172459 -8419 172460 -8408
rect 172640 -8413 172675 -8379
rect 172704 -8413 172747 -8379
rect 172749 -8413 172750 -8371
rect 172849 -8379 172850 -8371
rect 172784 -8413 172819 -8379
rect 172860 -8413 172895 -8379
rect 172905 -8413 172906 -8371
rect 173005 -8379 173006 -8371
rect 172954 -8413 172989 -8379
rect 173016 -8413 173061 -8379
rect 174056 -8408 174091 -8374
rect 174101 -8408 174102 -8363
rect 174201 -8374 174202 -8363
rect 174212 -8408 174247 -8374
rect 174257 -8408 174258 -8363
rect 174357 -8374 174358 -8363
rect 174933 -8367 174968 -8333
rect 175110 -8367 175145 -8333
rect 175703 -8336 175704 -8328
rect 175803 -8336 175804 -8328
rect 174368 -8408 174403 -8374
rect 172470 -8453 172505 -8419
rect 173749 -8422 173750 -8414
rect 175099 -8417 175100 -8406
rect 175304 -8410 175339 -8376
rect 175349 -8410 175350 -8365
rect 175449 -8376 175450 -8365
rect 175630 -8370 175693 -8336
rect 175702 -8370 175737 -8336
rect 175814 -8370 175849 -8336
rect 176539 -8360 176574 -8326
rect 176635 -8360 176670 -8326
rect 176731 -8360 176766 -8326
rect 176827 -8360 176862 -8326
rect 176923 -8360 176958 -8326
rect 177019 -8360 177054 -8326
rect 177115 -8360 177150 -8326
rect 178443 -8333 178444 -8322
rect 178620 -8327 178683 -8293
rect 178692 -8327 178727 -8293
rect 178804 -8327 178839 -8293
rect 179335 -8317 179370 -8283
rect 179431 -8317 179466 -8283
rect 179527 -8317 179562 -8283
rect 179623 -8317 179658 -8283
rect 179719 -8317 179754 -8283
rect 180744 -8324 180779 -8290
rect 180789 -8324 180790 -8279
rect 180889 -8290 180890 -8279
rect 180900 -8324 180935 -8290
rect 180945 -8324 180946 -8279
rect 181045 -8290 181046 -8279
rect 181224 -8284 181259 -8250
rect 181296 -8284 181331 -8250
rect 181368 -8284 181403 -8250
rect 181512 -8284 181547 -8250
rect 181584 -8284 181619 -8250
rect 181621 -8284 181691 -8250
rect 181728 -8284 181763 -8250
rect 181798 -8284 181833 -8250
rect 182325 -8274 182360 -8240
rect 182421 -8274 182456 -8240
rect 182517 -8274 182552 -8240
rect 184024 -8241 184059 -8207
rect 184088 -8241 184131 -8207
rect 184133 -8241 184134 -8199
rect 184233 -8207 184234 -8199
rect 184168 -8241 184203 -8207
rect 184244 -8241 184279 -8207
rect 184289 -8241 184290 -8199
rect 184389 -8207 184390 -8199
rect 184338 -8241 184373 -8207
rect 184400 -8241 184445 -8207
rect 185315 -8231 185350 -8197
rect 185411 -8231 185446 -8197
rect 185507 -8231 185542 -8197
rect 185131 -8250 185132 -8242
rect 181056 -8324 181091 -8290
rect 182037 -8293 182038 -8285
rect 182137 -8293 182138 -8285
rect 175460 -8410 175495 -8376
rect 172116 -8494 172151 -8460
rect 169126 -8620 169161 -8586
rect 170405 -8589 170406 -8578
rect 167655 -8689 167656 -8681
rect 167666 -8723 167701 -8689
rect 167886 -8734 167921 -8700
rect 166333 -8793 166368 -8759
rect 166536 -8838 166571 -8804
rect 166659 -8809 166660 -8767
rect 166981 -8796 167016 -8762
rect 166303 -8861 166304 -8853
rect 166314 -8895 166349 -8861
rect 166536 -8906 166571 -8872
rect 166303 -8961 166304 -8950
rect 166314 -8995 166349 -8961
rect 165251 -9045 165286 -9011
rect 165347 -9045 165382 -9011
rect 165443 -9045 165478 -9011
rect 165952 -9035 165987 -9001
rect 166024 -9035 166059 -9001
rect 166096 -9035 166131 -9001
rect 166168 -9029 166204 -9001
rect 166514 -9025 166549 -8991
rect 166559 -9025 166560 -8980
rect 166168 -9035 166203 -9029
rect 165605 -9088 165640 -9054
rect 165701 -9088 165736 -9054
rect 165797 -9088 165832 -9054
rect 166701 -9076 166702 -8809
rect 167330 -8819 167717 -8753
rect 166717 -8860 166752 -8826
rect 167066 -8832 167077 -8819
rect 167000 -8874 167077 -8832
rect 167128 -8874 167717 -8819
rect 167864 -8853 167899 -8819
rect 167909 -8853 167910 -8808
rect 167000 -8877 167717 -8874
rect 166717 -8928 166752 -8894
rect 166920 -8942 166955 -8908
rect 166965 -8942 166966 -8900
rect 166801 -8991 166802 -8980
rect 166812 -9025 166847 -8991
rect 166920 -9042 166955 -9008
rect 166965 -9042 166966 -8997
rect 166813 -9078 166848 -9044
rect 166885 -9078 166920 -9044
rect 166957 -9078 166992 -9044
rect 165959 -9131 165994 -9097
rect 166055 -9131 166090 -9097
rect 166151 -9131 166186 -9097
rect 166247 -9131 166282 -9097
rect 166343 -9131 166378 -9097
rect 167000 -9114 167145 -8877
rect 167330 -8899 167717 -8877
rect 167254 -8925 167717 -8899
rect 168051 -8904 168052 -8637
rect 168067 -8688 168102 -8654
rect 168681 -8691 168716 -8657
rect 169360 -8663 169395 -8629
rect 169405 -8663 169406 -8618
rect 169505 -8629 169506 -8618
rect 169516 -8663 169551 -8629
rect 169561 -8663 169562 -8618
rect 169661 -8629 169662 -8618
rect 170239 -8623 170274 -8589
rect 170416 -8623 170451 -8589
rect 170777 -8605 170812 -8571
rect 169672 -8663 169707 -8629
rect 169505 -8697 169506 -8671
rect 169904 -8689 169939 -8655
rect 169949 -8689 169950 -8644
rect 170049 -8655 170050 -8644
rect 170060 -8689 170095 -8655
rect 170105 -8689 170106 -8644
rect 170405 -8672 170406 -8661
rect 168067 -8756 168102 -8722
rect 168270 -8770 168305 -8736
rect 168315 -8770 168316 -8728
rect 168415 -8740 168416 -8729
rect 169035 -8734 169070 -8700
rect 168426 -8774 168461 -8740
rect 168151 -8819 168152 -8808
rect 168620 -8813 168655 -8779
rect 168665 -8813 168666 -8771
rect 168765 -8779 168766 -8771
rect 169425 -8777 169460 -8743
rect 168776 -8813 168811 -8779
rect 168162 -8853 168197 -8819
rect 168270 -8870 168305 -8836
rect 168315 -8870 168316 -8825
rect 168415 -8832 168416 -8821
rect 168426 -8866 168461 -8832
rect 168974 -8856 169009 -8822
rect 169019 -8856 169020 -8814
rect 169119 -8822 169120 -8814
rect 169130 -8856 169165 -8822
rect 168163 -8906 168198 -8872
rect 168235 -8906 168270 -8872
rect 168307 -8906 168342 -8872
rect 168620 -8913 168655 -8879
rect 168665 -8913 168666 -8868
rect 168765 -8879 168766 -8868
rect 168776 -8913 168811 -8879
rect 169360 -8895 169395 -8861
rect 169405 -8895 169406 -8853
rect 167254 -8959 167730 -8925
rect 168588 -8949 168623 -8915
rect 168660 -8949 168695 -8915
rect 168974 -8956 169009 -8922
rect 169019 -8956 169020 -8911
rect 169119 -8922 169120 -8911
rect 169130 -8956 169165 -8922
rect 167254 -8985 167717 -8959
rect 167258 -8993 167459 -8985
rect 167274 -9003 167443 -8993
rect 167000 -9140 167175 -9114
rect 166507 -9174 166542 -9140
rect 166603 -9174 166638 -9140
rect 166699 -9174 166734 -9140
rect 166795 -9174 166830 -9140
rect 166891 -9174 166926 -9140
rect 166987 -9174 167175 -9140
rect 167000 -9200 167175 -9174
rect 167200 -9174 167301 -9050
rect 167078 -9870 167113 -9200
rect 167200 -9228 167203 -9174
rect 166885 -9936 167030 -9924
rect 166553 -9970 167030 -9936
rect 166885 -9971 167030 -9970
rect 167066 -9971 167113 -9870
rect 167212 -9971 167247 -9174
rect 167470 -9971 167505 -9062
rect 167604 -9971 167639 -8985
rect 167857 -9002 167892 -8968
rect 167953 -9002 167988 -8968
rect 168049 -9002 168084 -8968
rect 168145 -9002 168180 -8968
rect 168241 -9002 168276 -8968
rect 168337 -9002 168372 -8968
rect 168433 -9002 168468 -8968
rect 168942 -8992 168977 -8958
rect 169014 -8992 169049 -8958
rect 169360 -8995 169395 -8961
rect 169405 -8995 169406 -8950
rect 169547 -9001 169548 -8697
rect 170239 -8706 170274 -8672
rect 170416 -8706 170451 -8672
rect 170712 -8723 170747 -8689
rect 170757 -8723 170758 -8681
rect 170899 -8753 170900 -8525
rect 171589 -8534 171624 -8500
rect 171766 -8534 171801 -8500
rect 171960 -8577 171995 -8543
rect 172005 -8577 172006 -8532
rect 172105 -8543 172106 -8532
rect 172314 -8537 172349 -8503
rect 172359 -8537 172360 -8492
rect 172459 -8503 172460 -8492
rect 172704 -8496 172739 -8462
rect 172749 -8496 172750 -8451
rect 172849 -8462 172850 -8451
rect 172860 -8496 172895 -8462
rect 172905 -8496 172906 -8451
rect 173005 -8462 173006 -8451
rect 173186 -8456 173221 -8422
rect 173258 -8456 173293 -8422
rect 173330 -8456 173365 -8422
rect 173474 -8456 173509 -8422
rect 173546 -8456 173581 -8422
rect 173583 -8456 173653 -8422
rect 173690 -8456 173725 -8422
rect 173760 -8456 173795 -8422
rect 173016 -8496 173051 -8462
rect 174056 -8491 174091 -8457
rect 174101 -8491 174102 -8446
rect 174201 -8457 174202 -8446
rect 174212 -8491 174247 -8457
rect 174257 -8491 174258 -8446
rect 174357 -8457 174358 -8446
rect 174933 -8451 174968 -8417
rect 175110 -8451 175145 -8417
rect 174368 -8491 174403 -8457
rect 172470 -8537 172505 -8503
rect 173749 -8505 173750 -8494
rect 172116 -8577 172151 -8543
rect 171029 -8621 171064 -8587
rect 171230 -8666 171265 -8632
rect 171353 -8637 171354 -8595
rect 171675 -8624 171710 -8590
rect 172314 -8620 172349 -8586
rect 172359 -8620 172360 -8575
rect 172459 -8586 172460 -8575
rect 172704 -8580 172739 -8546
rect 172749 -8580 172750 -8535
rect 172849 -8546 172850 -8535
rect 172860 -8580 172895 -8546
rect 172905 -8580 172906 -8535
rect 173005 -8546 173006 -8535
rect 173583 -8539 173618 -8505
rect 173760 -8539 173795 -8505
rect 173016 -8580 173051 -8546
rect 173903 -8565 174018 -8499
rect 174201 -8525 174202 -8499
rect 174598 -8517 174633 -8483
rect 174643 -8517 174644 -8472
rect 174743 -8483 174744 -8472
rect 174754 -8517 174789 -8483
rect 174799 -8517 174800 -8472
rect 175099 -8500 175100 -8489
rect 175304 -8494 175339 -8460
rect 175349 -8494 175350 -8449
rect 175449 -8460 175450 -8449
rect 175658 -8453 175693 -8419
rect 175703 -8453 175704 -8408
rect 175803 -8419 175804 -8408
rect 175984 -8413 176019 -8379
rect 176048 -8413 176091 -8379
rect 176093 -8413 176094 -8371
rect 176193 -8379 176194 -8371
rect 176128 -8413 176163 -8379
rect 176204 -8413 176239 -8379
rect 176249 -8413 176250 -8371
rect 176349 -8379 176350 -8371
rect 176298 -8413 176333 -8379
rect 176360 -8413 176405 -8379
rect 177400 -8408 177435 -8374
rect 177445 -8408 177446 -8363
rect 177545 -8374 177546 -8363
rect 177556 -8408 177591 -8374
rect 177601 -8408 177602 -8363
rect 177701 -8374 177702 -8363
rect 178277 -8367 178312 -8333
rect 178454 -8367 178489 -8333
rect 179047 -8336 179048 -8328
rect 179147 -8336 179148 -8328
rect 177712 -8408 177747 -8374
rect 175814 -8453 175849 -8419
rect 177093 -8422 177094 -8414
rect 178443 -8417 178444 -8406
rect 178648 -8410 178683 -8376
rect 178693 -8410 178694 -8365
rect 178793 -8376 178794 -8365
rect 178974 -8370 179037 -8336
rect 179046 -8370 179081 -8336
rect 179158 -8370 179193 -8336
rect 179883 -8360 179918 -8326
rect 179979 -8360 180014 -8326
rect 180075 -8360 180110 -8326
rect 180171 -8360 180206 -8326
rect 180267 -8360 180302 -8326
rect 180363 -8360 180398 -8326
rect 180459 -8360 180494 -8326
rect 181787 -8333 181788 -8322
rect 181964 -8327 182027 -8293
rect 182036 -8327 182071 -8293
rect 182148 -8327 182183 -8293
rect 182679 -8317 182714 -8283
rect 182775 -8317 182810 -8283
rect 182871 -8317 182906 -8283
rect 182967 -8317 183002 -8283
rect 183063 -8317 183098 -8283
rect 184088 -8324 184123 -8290
rect 184133 -8324 184134 -8279
rect 184233 -8290 184234 -8279
rect 184244 -8324 184279 -8290
rect 184289 -8324 184290 -8279
rect 184389 -8290 184390 -8279
rect 184568 -8284 184603 -8250
rect 184640 -8284 184675 -8250
rect 184712 -8284 184747 -8250
rect 184856 -8284 184891 -8250
rect 184928 -8284 184963 -8250
rect 184965 -8284 185035 -8250
rect 185072 -8284 185107 -8250
rect 185142 -8284 185177 -8250
rect 185669 -8274 185704 -8240
rect 185765 -8274 185800 -8240
rect 185861 -8274 185896 -8240
rect 187368 -8241 187403 -8207
rect 187432 -8241 187475 -8207
rect 187477 -8241 187478 -8199
rect 187577 -8207 187578 -8199
rect 187512 -8241 187547 -8207
rect 187588 -8241 187623 -8207
rect 187633 -8241 187634 -8199
rect 187733 -8207 187734 -8199
rect 187682 -8241 187717 -8207
rect 187744 -8241 187789 -8207
rect 188659 -8231 188694 -8197
rect 188755 -8231 188790 -8197
rect 188851 -8231 188886 -8197
rect 188475 -8250 188476 -8242
rect 184400 -8324 184435 -8290
rect 185381 -8293 185382 -8285
rect 185481 -8293 185482 -8285
rect 178804 -8410 178839 -8376
rect 175460 -8494 175495 -8460
rect 172470 -8620 172505 -8586
rect 173749 -8589 173750 -8578
rect 170999 -8689 171000 -8681
rect 171010 -8723 171045 -8689
rect 171230 -8734 171265 -8700
rect 169677 -8793 169712 -8759
rect 169880 -8838 169915 -8804
rect 170003 -8809 170004 -8767
rect 170325 -8796 170360 -8762
rect 169647 -8861 169648 -8853
rect 169658 -8895 169693 -8861
rect 169880 -8906 169915 -8872
rect 169647 -8961 169648 -8950
rect 169658 -8995 169693 -8961
rect 168595 -9045 168630 -9011
rect 168691 -9045 168726 -9011
rect 168787 -9045 168822 -9011
rect 169296 -9035 169331 -9001
rect 169368 -9035 169403 -9001
rect 169440 -9035 169475 -9001
rect 169512 -9029 169548 -9001
rect 169858 -9025 169893 -8991
rect 169903 -9025 169904 -8980
rect 169512 -9035 169547 -9029
rect 168949 -9088 168984 -9054
rect 169045 -9088 169080 -9054
rect 169141 -9088 169176 -9054
rect 170045 -9076 170046 -8809
rect 170674 -8819 171061 -8753
rect 170061 -8860 170096 -8826
rect 170410 -8832 170421 -8819
rect 170344 -8874 170421 -8832
rect 170472 -8874 171061 -8819
rect 171208 -8853 171243 -8819
rect 171253 -8853 171254 -8808
rect 170344 -8877 171061 -8874
rect 170061 -8928 170096 -8894
rect 170264 -8942 170299 -8908
rect 170309 -8942 170310 -8900
rect 170145 -8991 170146 -8980
rect 170156 -9025 170191 -8991
rect 170264 -9042 170299 -9008
rect 170309 -9042 170310 -8997
rect 170157 -9078 170192 -9044
rect 170229 -9078 170264 -9044
rect 170301 -9078 170336 -9044
rect 169303 -9131 169338 -9097
rect 169399 -9131 169434 -9097
rect 169495 -9131 169530 -9097
rect 169591 -9131 169626 -9097
rect 169687 -9131 169722 -9097
rect 170344 -9114 170489 -8877
rect 170674 -8899 171061 -8877
rect 170598 -8925 171061 -8899
rect 171395 -8904 171396 -8637
rect 171411 -8688 171446 -8654
rect 172025 -8691 172060 -8657
rect 172704 -8663 172739 -8629
rect 172749 -8663 172750 -8618
rect 172849 -8629 172850 -8618
rect 172860 -8663 172895 -8629
rect 172905 -8663 172906 -8618
rect 173005 -8629 173006 -8618
rect 173583 -8623 173618 -8589
rect 173760 -8623 173795 -8589
rect 174121 -8605 174156 -8571
rect 173016 -8663 173051 -8629
rect 172849 -8697 172850 -8671
rect 173248 -8689 173283 -8655
rect 173293 -8689 173294 -8644
rect 173393 -8655 173394 -8644
rect 173404 -8689 173439 -8655
rect 173449 -8689 173450 -8644
rect 173749 -8672 173750 -8661
rect 171411 -8756 171446 -8722
rect 171614 -8770 171649 -8736
rect 171659 -8770 171660 -8728
rect 171759 -8740 171760 -8729
rect 172379 -8734 172414 -8700
rect 171770 -8774 171805 -8740
rect 171495 -8819 171496 -8808
rect 171964 -8813 171999 -8779
rect 172009 -8813 172010 -8771
rect 172109 -8779 172110 -8771
rect 172769 -8777 172804 -8743
rect 172120 -8813 172155 -8779
rect 171506 -8853 171541 -8819
rect 171614 -8870 171649 -8836
rect 171659 -8870 171660 -8825
rect 171759 -8832 171760 -8821
rect 171770 -8866 171805 -8832
rect 172318 -8856 172353 -8822
rect 172363 -8856 172364 -8814
rect 172463 -8822 172464 -8814
rect 172474 -8856 172509 -8822
rect 171507 -8906 171542 -8872
rect 171579 -8906 171614 -8872
rect 171651 -8906 171686 -8872
rect 171964 -8913 171999 -8879
rect 172009 -8913 172010 -8868
rect 172109 -8879 172110 -8868
rect 172120 -8913 172155 -8879
rect 172704 -8895 172739 -8861
rect 172749 -8895 172750 -8853
rect 170598 -8959 171074 -8925
rect 171932 -8949 171967 -8915
rect 172004 -8949 172039 -8915
rect 172318 -8956 172353 -8922
rect 172363 -8956 172364 -8911
rect 172463 -8922 172464 -8911
rect 172474 -8956 172509 -8922
rect 170598 -8985 171061 -8959
rect 170602 -8993 170803 -8985
rect 170618 -9003 170787 -8993
rect 170344 -9140 170519 -9114
rect 169851 -9174 169886 -9140
rect 169947 -9174 169982 -9140
rect 170043 -9174 170078 -9140
rect 170139 -9174 170174 -9140
rect 170235 -9174 170270 -9140
rect 170331 -9174 170519 -9140
rect 170344 -9200 170519 -9174
rect 170544 -9174 170645 -9050
rect 170422 -9870 170457 -9200
rect 170544 -9228 170547 -9174
rect 170229 -9936 170374 -9924
rect 169897 -9970 170374 -9936
rect 170229 -9971 170374 -9970
rect 170410 -9971 170457 -9870
rect 170556 -9971 170591 -9174
rect 170814 -9971 170849 -9062
rect 170948 -9971 170983 -8985
rect 171201 -9002 171236 -8968
rect 171297 -9002 171332 -8968
rect 171393 -9002 171428 -8968
rect 171489 -9002 171524 -8968
rect 171585 -9002 171620 -8968
rect 171681 -9002 171716 -8968
rect 171777 -9002 171812 -8968
rect 172286 -8992 172321 -8958
rect 172358 -8992 172393 -8958
rect 172704 -8995 172739 -8961
rect 172749 -8995 172750 -8950
rect 172891 -9001 172892 -8697
rect 173583 -8706 173618 -8672
rect 173760 -8706 173795 -8672
rect 174056 -8723 174091 -8689
rect 174101 -8723 174102 -8681
rect 174243 -8753 174244 -8525
rect 174933 -8534 174968 -8500
rect 175110 -8534 175145 -8500
rect 175304 -8577 175339 -8543
rect 175349 -8577 175350 -8532
rect 175449 -8543 175450 -8532
rect 175658 -8537 175693 -8503
rect 175703 -8537 175704 -8492
rect 175803 -8503 175804 -8492
rect 176048 -8496 176083 -8462
rect 176093 -8496 176094 -8451
rect 176193 -8462 176194 -8451
rect 176204 -8496 176239 -8462
rect 176249 -8496 176250 -8451
rect 176349 -8462 176350 -8451
rect 176530 -8456 176565 -8422
rect 176602 -8456 176637 -8422
rect 176674 -8456 176709 -8422
rect 176818 -8456 176853 -8422
rect 176890 -8456 176925 -8422
rect 176927 -8456 176997 -8422
rect 177034 -8456 177069 -8422
rect 177104 -8456 177139 -8422
rect 176360 -8496 176395 -8462
rect 177400 -8491 177435 -8457
rect 177445 -8491 177446 -8446
rect 177545 -8457 177546 -8446
rect 177556 -8491 177591 -8457
rect 177601 -8491 177602 -8446
rect 177701 -8457 177702 -8446
rect 178277 -8451 178312 -8417
rect 178454 -8451 178489 -8417
rect 177712 -8491 177747 -8457
rect 175814 -8537 175849 -8503
rect 177093 -8505 177094 -8494
rect 175460 -8577 175495 -8543
rect 174373 -8621 174408 -8587
rect 174574 -8666 174609 -8632
rect 174697 -8637 174698 -8595
rect 175019 -8624 175054 -8590
rect 175658 -8620 175693 -8586
rect 175703 -8620 175704 -8575
rect 175803 -8586 175804 -8575
rect 176048 -8580 176083 -8546
rect 176093 -8580 176094 -8535
rect 176193 -8546 176194 -8535
rect 176204 -8580 176239 -8546
rect 176249 -8580 176250 -8535
rect 176349 -8546 176350 -8535
rect 176927 -8539 176962 -8505
rect 177104 -8539 177139 -8505
rect 176360 -8580 176395 -8546
rect 177247 -8565 177362 -8499
rect 177545 -8525 177546 -8499
rect 177942 -8517 177977 -8483
rect 177987 -8517 177988 -8472
rect 178087 -8483 178088 -8472
rect 178098 -8517 178133 -8483
rect 178143 -8517 178144 -8472
rect 178443 -8500 178444 -8489
rect 178648 -8494 178683 -8460
rect 178693 -8494 178694 -8449
rect 178793 -8460 178794 -8449
rect 179002 -8453 179037 -8419
rect 179047 -8453 179048 -8408
rect 179147 -8419 179148 -8408
rect 179328 -8413 179363 -8379
rect 179392 -8413 179435 -8379
rect 179437 -8413 179438 -8371
rect 179537 -8379 179538 -8371
rect 179472 -8413 179507 -8379
rect 179548 -8413 179583 -8379
rect 179593 -8413 179594 -8371
rect 179693 -8379 179694 -8371
rect 179642 -8413 179677 -8379
rect 179704 -8413 179749 -8379
rect 180744 -8408 180779 -8374
rect 180789 -8408 180790 -8363
rect 180889 -8374 180890 -8363
rect 180900 -8408 180935 -8374
rect 180945 -8408 180946 -8363
rect 181045 -8374 181046 -8363
rect 181621 -8367 181656 -8333
rect 181798 -8367 181833 -8333
rect 182391 -8336 182392 -8328
rect 182491 -8336 182492 -8328
rect 181056 -8408 181091 -8374
rect 179158 -8453 179193 -8419
rect 180437 -8422 180438 -8414
rect 181787 -8417 181788 -8406
rect 181992 -8410 182027 -8376
rect 182037 -8410 182038 -8365
rect 182137 -8376 182138 -8365
rect 182318 -8370 182381 -8336
rect 182390 -8370 182425 -8336
rect 182502 -8370 182537 -8336
rect 183227 -8360 183262 -8326
rect 183323 -8360 183358 -8326
rect 183419 -8360 183454 -8326
rect 183515 -8360 183550 -8326
rect 183611 -8360 183646 -8326
rect 183707 -8360 183742 -8326
rect 183803 -8360 183838 -8326
rect 185131 -8333 185132 -8322
rect 185308 -8327 185371 -8293
rect 185380 -8327 185415 -8293
rect 185492 -8327 185527 -8293
rect 186023 -8317 186058 -8283
rect 186119 -8317 186154 -8283
rect 186215 -8317 186250 -8283
rect 186311 -8317 186346 -8283
rect 186407 -8317 186442 -8283
rect 187432 -8324 187467 -8290
rect 187477 -8324 187478 -8279
rect 187577 -8290 187578 -8279
rect 187588 -8324 187623 -8290
rect 187633 -8324 187634 -8279
rect 187733 -8290 187734 -8279
rect 187912 -8284 187947 -8250
rect 187984 -8284 188019 -8250
rect 188056 -8284 188091 -8250
rect 188200 -8284 188235 -8250
rect 188272 -8284 188307 -8250
rect 188309 -8284 188379 -8250
rect 188416 -8284 188451 -8250
rect 188486 -8284 188521 -8250
rect 189013 -8274 189048 -8240
rect 189109 -8274 189144 -8240
rect 189205 -8274 189240 -8240
rect 190712 -8241 190747 -8207
rect 190776 -8241 190819 -8207
rect 190821 -8241 190822 -8199
rect 190921 -8207 190922 -8199
rect 190856 -8241 190891 -8207
rect 190932 -8241 190967 -8207
rect 190977 -8241 190978 -8199
rect 191077 -8207 191078 -8199
rect 191026 -8241 191061 -8207
rect 191088 -8241 191133 -8207
rect 192003 -8231 192038 -8197
rect 192099 -8231 192134 -8197
rect 192195 -8231 192230 -8197
rect 191819 -8250 191820 -8242
rect 187744 -8324 187779 -8290
rect 188725 -8293 188726 -8285
rect 188825 -8293 188826 -8285
rect 182148 -8410 182183 -8376
rect 178804 -8494 178839 -8460
rect 175814 -8620 175849 -8586
rect 177093 -8589 177094 -8578
rect 174343 -8689 174344 -8681
rect 174354 -8723 174389 -8689
rect 174574 -8734 174609 -8700
rect 173021 -8793 173056 -8759
rect 173224 -8838 173259 -8804
rect 173347 -8809 173348 -8767
rect 173669 -8796 173704 -8762
rect 172991 -8861 172992 -8853
rect 173002 -8895 173037 -8861
rect 173224 -8906 173259 -8872
rect 172991 -8961 172992 -8950
rect 173002 -8995 173037 -8961
rect 171939 -9045 171974 -9011
rect 172035 -9045 172070 -9011
rect 172131 -9045 172166 -9011
rect 172640 -9035 172675 -9001
rect 172712 -9035 172747 -9001
rect 172784 -9035 172819 -9001
rect 172856 -9029 172892 -9001
rect 173202 -9025 173237 -8991
rect 173247 -9025 173248 -8980
rect 172856 -9035 172891 -9029
rect 172293 -9088 172328 -9054
rect 172389 -9088 172424 -9054
rect 172485 -9088 172520 -9054
rect 173389 -9076 173390 -8809
rect 174018 -8819 174405 -8753
rect 173405 -8860 173440 -8826
rect 173754 -8832 173765 -8819
rect 173688 -8874 173765 -8832
rect 173816 -8874 174405 -8819
rect 174552 -8853 174587 -8819
rect 174597 -8853 174598 -8808
rect 173688 -8877 174405 -8874
rect 173405 -8928 173440 -8894
rect 173608 -8942 173643 -8908
rect 173653 -8942 173654 -8900
rect 173489 -8991 173490 -8980
rect 173500 -9025 173535 -8991
rect 173608 -9042 173643 -9008
rect 173653 -9042 173654 -8997
rect 173501 -9078 173536 -9044
rect 173573 -9078 173608 -9044
rect 173645 -9078 173680 -9044
rect 172647 -9131 172682 -9097
rect 172743 -9131 172778 -9097
rect 172839 -9131 172874 -9097
rect 172935 -9131 172970 -9097
rect 173031 -9131 173066 -9097
rect 173688 -9114 173833 -8877
rect 174018 -8899 174405 -8877
rect 173942 -8925 174405 -8899
rect 174739 -8904 174740 -8637
rect 174755 -8688 174790 -8654
rect 175369 -8691 175404 -8657
rect 176048 -8663 176083 -8629
rect 176093 -8663 176094 -8618
rect 176193 -8629 176194 -8618
rect 176204 -8663 176239 -8629
rect 176249 -8663 176250 -8618
rect 176349 -8629 176350 -8618
rect 176927 -8623 176962 -8589
rect 177104 -8623 177139 -8589
rect 177465 -8605 177500 -8571
rect 176360 -8663 176395 -8629
rect 176193 -8697 176194 -8671
rect 176592 -8689 176627 -8655
rect 176637 -8689 176638 -8644
rect 176737 -8655 176738 -8644
rect 176748 -8689 176783 -8655
rect 176793 -8689 176794 -8644
rect 177093 -8672 177094 -8661
rect 174755 -8756 174790 -8722
rect 174958 -8770 174993 -8736
rect 175003 -8770 175004 -8728
rect 175103 -8740 175104 -8729
rect 175723 -8734 175758 -8700
rect 175114 -8774 175149 -8740
rect 174839 -8819 174840 -8808
rect 175308 -8813 175343 -8779
rect 175353 -8813 175354 -8771
rect 175453 -8779 175454 -8771
rect 176113 -8777 176148 -8743
rect 175464 -8813 175499 -8779
rect 174850 -8853 174885 -8819
rect 174958 -8870 174993 -8836
rect 175003 -8870 175004 -8825
rect 175103 -8832 175104 -8821
rect 175114 -8866 175149 -8832
rect 175662 -8856 175697 -8822
rect 175707 -8856 175708 -8814
rect 175807 -8822 175808 -8814
rect 175818 -8856 175853 -8822
rect 174851 -8906 174886 -8872
rect 174923 -8906 174958 -8872
rect 174995 -8906 175030 -8872
rect 175308 -8913 175343 -8879
rect 175353 -8913 175354 -8868
rect 175453 -8879 175454 -8868
rect 175464 -8913 175499 -8879
rect 176048 -8895 176083 -8861
rect 176093 -8895 176094 -8853
rect 173942 -8959 174418 -8925
rect 175276 -8949 175311 -8915
rect 175348 -8949 175383 -8915
rect 175662 -8956 175697 -8922
rect 175707 -8956 175708 -8911
rect 175807 -8922 175808 -8911
rect 175818 -8956 175853 -8922
rect 173942 -8985 174405 -8959
rect 173946 -8993 174147 -8985
rect 173962 -9003 174131 -8993
rect 173688 -9140 173863 -9114
rect 173195 -9174 173230 -9140
rect 173291 -9174 173326 -9140
rect 173387 -9174 173422 -9140
rect 173483 -9174 173518 -9140
rect 173579 -9174 173614 -9140
rect 173675 -9174 173863 -9140
rect 173688 -9200 173863 -9174
rect 173888 -9174 173989 -9050
rect 173766 -9870 173801 -9200
rect 173888 -9228 173891 -9174
rect 173573 -9936 173718 -9924
rect 173241 -9970 173718 -9936
rect 173573 -9971 173718 -9970
rect 173754 -9971 173801 -9870
rect 173900 -9971 173935 -9174
rect 174158 -9971 174193 -9062
rect 174292 -9971 174327 -8985
rect 174545 -9002 174580 -8968
rect 174641 -9002 174676 -8968
rect 174737 -9002 174772 -8968
rect 174833 -9002 174868 -8968
rect 174929 -9002 174964 -8968
rect 175025 -9002 175060 -8968
rect 175121 -9002 175156 -8968
rect 175630 -8992 175665 -8958
rect 175702 -8992 175737 -8958
rect 176048 -8995 176083 -8961
rect 176093 -8995 176094 -8950
rect 176235 -9001 176236 -8697
rect 176927 -8706 176962 -8672
rect 177104 -8706 177139 -8672
rect 177400 -8723 177435 -8689
rect 177445 -8723 177446 -8681
rect 177587 -8753 177588 -8525
rect 178277 -8534 178312 -8500
rect 178454 -8534 178489 -8500
rect 178648 -8577 178683 -8543
rect 178693 -8577 178694 -8532
rect 178793 -8543 178794 -8532
rect 179002 -8537 179037 -8503
rect 179047 -8537 179048 -8492
rect 179147 -8503 179148 -8492
rect 179392 -8496 179427 -8462
rect 179437 -8496 179438 -8451
rect 179537 -8462 179538 -8451
rect 179548 -8496 179583 -8462
rect 179593 -8496 179594 -8451
rect 179693 -8462 179694 -8451
rect 179874 -8456 179909 -8422
rect 179946 -8456 179981 -8422
rect 180018 -8456 180053 -8422
rect 180162 -8456 180197 -8422
rect 180234 -8456 180269 -8422
rect 180271 -8456 180341 -8422
rect 180378 -8456 180413 -8422
rect 180448 -8456 180483 -8422
rect 179704 -8496 179739 -8462
rect 180744 -8491 180779 -8457
rect 180789 -8491 180790 -8446
rect 180889 -8457 180890 -8446
rect 180900 -8491 180935 -8457
rect 180945 -8491 180946 -8446
rect 181045 -8457 181046 -8446
rect 181621 -8451 181656 -8417
rect 181798 -8451 181833 -8417
rect 181056 -8491 181091 -8457
rect 179158 -8537 179193 -8503
rect 180437 -8505 180438 -8494
rect 178804 -8577 178839 -8543
rect 177717 -8621 177752 -8587
rect 177918 -8666 177953 -8632
rect 178041 -8637 178042 -8595
rect 178363 -8624 178398 -8590
rect 179002 -8620 179037 -8586
rect 179047 -8620 179048 -8575
rect 179147 -8586 179148 -8575
rect 179392 -8580 179427 -8546
rect 179437 -8580 179438 -8535
rect 179537 -8546 179538 -8535
rect 179548 -8580 179583 -8546
rect 179593 -8580 179594 -8535
rect 179693 -8546 179694 -8535
rect 180271 -8539 180306 -8505
rect 180448 -8539 180483 -8505
rect 179704 -8580 179739 -8546
rect 180591 -8565 180706 -8499
rect 180889 -8525 180890 -8499
rect 181286 -8517 181321 -8483
rect 181331 -8517 181332 -8472
rect 181431 -8483 181432 -8472
rect 181442 -8517 181477 -8483
rect 181487 -8517 181488 -8472
rect 181787 -8500 181788 -8489
rect 181992 -8494 182027 -8460
rect 182037 -8494 182038 -8449
rect 182137 -8460 182138 -8449
rect 182346 -8453 182381 -8419
rect 182391 -8453 182392 -8408
rect 182491 -8419 182492 -8408
rect 182672 -8413 182707 -8379
rect 182736 -8413 182779 -8379
rect 182781 -8413 182782 -8371
rect 182881 -8379 182882 -8371
rect 182816 -8413 182851 -8379
rect 182892 -8413 182927 -8379
rect 182937 -8413 182938 -8371
rect 183037 -8379 183038 -8371
rect 182986 -8413 183021 -8379
rect 183048 -8413 183093 -8379
rect 184088 -8408 184123 -8374
rect 184133 -8408 184134 -8363
rect 184233 -8374 184234 -8363
rect 184244 -8408 184279 -8374
rect 184289 -8408 184290 -8363
rect 184389 -8374 184390 -8363
rect 184965 -8367 185000 -8333
rect 185142 -8367 185177 -8333
rect 185735 -8336 185736 -8328
rect 185835 -8336 185836 -8328
rect 184400 -8408 184435 -8374
rect 182502 -8453 182537 -8419
rect 183781 -8422 183782 -8414
rect 185131 -8417 185132 -8406
rect 185336 -8410 185371 -8376
rect 185381 -8410 185382 -8365
rect 185481 -8376 185482 -8365
rect 185662 -8370 185725 -8336
rect 185734 -8370 185769 -8336
rect 185846 -8370 185881 -8336
rect 186571 -8360 186606 -8326
rect 186667 -8360 186702 -8326
rect 186763 -8360 186798 -8326
rect 186859 -8360 186894 -8326
rect 186955 -8360 186990 -8326
rect 187051 -8360 187086 -8326
rect 187147 -8360 187182 -8326
rect 188475 -8333 188476 -8322
rect 188652 -8327 188715 -8293
rect 188724 -8327 188759 -8293
rect 188836 -8327 188871 -8293
rect 189367 -8317 189402 -8283
rect 189463 -8317 189498 -8283
rect 189559 -8317 189594 -8283
rect 189655 -8317 189690 -8283
rect 189751 -8317 189786 -8283
rect 190776 -8324 190811 -8290
rect 190821 -8324 190822 -8279
rect 190921 -8290 190922 -8279
rect 190932 -8324 190967 -8290
rect 190977 -8324 190978 -8279
rect 191077 -8290 191078 -8279
rect 191256 -8284 191291 -8250
rect 191328 -8284 191363 -8250
rect 191400 -8284 191435 -8250
rect 191544 -8284 191579 -8250
rect 191616 -8284 191651 -8250
rect 191653 -8284 191723 -8250
rect 191760 -8284 191795 -8250
rect 191830 -8284 191865 -8250
rect 192357 -8274 192392 -8240
rect 192453 -8274 192488 -8240
rect 192549 -8274 192584 -8240
rect 194056 -8241 194091 -8207
rect 194120 -8241 194163 -8207
rect 194165 -8241 194166 -8199
rect 194265 -8207 194266 -8199
rect 194200 -8241 194235 -8207
rect 194276 -8241 194311 -8207
rect 194321 -8241 194322 -8199
rect 194421 -8207 194422 -8199
rect 194370 -8241 194405 -8207
rect 194432 -8241 194477 -8207
rect 195347 -8231 195382 -8197
rect 195443 -8231 195478 -8197
rect 195539 -8231 195574 -8197
rect 195163 -8250 195164 -8242
rect 191088 -8324 191123 -8290
rect 192069 -8293 192070 -8285
rect 192169 -8293 192170 -8285
rect 185492 -8410 185527 -8376
rect 182148 -8494 182183 -8460
rect 179158 -8620 179193 -8586
rect 180437 -8589 180438 -8578
rect 177687 -8689 177688 -8681
rect 177698 -8723 177733 -8689
rect 177918 -8734 177953 -8700
rect 176365 -8793 176400 -8759
rect 176568 -8838 176603 -8804
rect 176691 -8809 176692 -8767
rect 177013 -8796 177048 -8762
rect 176335 -8861 176336 -8853
rect 176346 -8895 176381 -8861
rect 176568 -8906 176603 -8872
rect 176335 -8961 176336 -8950
rect 176346 -8995 176381 -8961
rect 175283 -9045 175318 -9011
rect 175379 -9045 175414 -9011
rect 175475 -9045 175510 -9011
rect 175984 -9035 176019 -9001
rect 176056 -9035 176091 -9001
rect 176128 -9035 176163 -9001
rect 176200 -9029 176236 -9001
rect 176546 -9025 176581 -8991
rect 176591 -9025 176592 -8980
rect 176200 -9035 176235 -9029
rect 175637 -9088 175672 -9054
rect 175733 -9088 175768 -9054
rect 175829 -9088 175864 -9054
rect 176733 -9076 176734 -8809
rect 177362 -8819 177749 -8753
rect 176749 -8860 176784 -8826
rect 177098 -8832 177109 -8819
rect 177032 -8874 177109 -8832
rect 177160 -8874 177749 -8819
rect 177896 -8853 177931 -8819
rect 177941 -8853 177942 -8808
rect 177032 -8877 177749 -8874
rect 176749 -8928 176784 -8894
rect 176952 -8942 176987 -8908
rect 176997 -8942 176998 -8900
rect 176833 -8991 176834 -8980
rect 176844 -9025 176879 -8991
rect 176952 -9042 176987 -9008
rect 176997 -9042 176998 -8997
rect 176845 -9078 176880 -9044
rect 176917 -9078 176952 -9044
rect 176989 -9078 177024 -9044
rect 175991 -9131 176026 -9097
rect 176087 -9131 176122 -9097
rect 176183 -9131 176218 -9097
rect 176279 -9131 176314 -9097
rect 176375 -9131 176410 -9097
rect 177032 -9114 177177 -8877
rect 177362 -8899 177749 -8877
rect 177286 -8925 177749 -8899
rect 178083 -8904 178084 -8637
rect 178099 -8688 178134 -8654
rect 178713 -8691 178748 -8657
rect 179392 -8663 179427 -8629
rect 179437 -8663 179438 -8618
rect 179537 -8629 179538 -8618
rect 179548 -8663 179583 -8629
rect 179593 -8663 179594 -8618
rect 179693 -8629 179694 -8618
rect 180271 -8623 180306 -8589
rect 180448 -8623 180483 -8589
rect 180809 -8605 180844 -8571
rect 179704 -8663 179739 -8629
rect 179537 -8697 179538 -8671
rect 179936 -8689 179971 -8655
rect 179981 -8689 179982 -8644
rect 180081 -8655 180082 -8644
rect 180092 -8689 180127 -8655
rect 180137 -8689 180138 -8644
rect 180437 -8672 180438 -8661
rect 178099 -8756 178134 -8722
rect 178302 -8770 178337 -8736
rect 178347 -8770 178348 -8728
rect 178447 -8740 178448 -8729
rect 179067 -8734 179102 -8700
rect 178458 -8774 178493 -8740
rect 178183 -8819 178184 -8808
rect 178652 -8813 178687 -8779
rect 178697 -8813 178698 -8771
rect 178797 -8779 178798 -8771
rect 179457 -8777 179492 -8743
rect 178808 -8813 178843 -8779
rect 178194 -8853 178229 -8819
rect 178302 -8870 178337 -8836
rect 178347 -8870 178348 -8825
rect 178447 -8832 178448 -8821
rect 178458 -8866 178493 -8832
rect 179006 -8856 179041 -8822
rect 179051 -8856 179052 -8814
rect 179151 -8822 179152 -8814
rect 179162 -8856 179197 -8822
rect 178195 -8906 178230 -8872
rect 178267 -8906 178302 -8872
rect 178339 -8906 178374 -8872
rect 178652 -8913 178687 -8879
rect 178697 -8913 178698 -8868
rect 178797 -8879 178798 -8868
rect 178808 -8913 178843 -8879
rect 179392 -8895 179427 -8861
rect 179437 -8895 179438 -8853
rect 177286 -8959 177762 -8925
rect 178620 -8949 178655 -8915
rect 178692 -8949 178727 -8915
rect 179006 -8956 179041 -8922
rect 179051 -8956 179052 -8911
rect 179151 -8922 179152 -8911
rect 179162 -8956 179197 -8922
rect 177286 -8985 177749 -8959
rect 177290 -8993 177491 -8985
rect 177306 -9003 177475 -8993
rect 177032 -9140 177207 -9114
rect 176539 -9174 176574 -9140
rect 176635 -9174 176670 -9140
rect 176731 -9174 176766 -9140
rect 176827 -9174 176862 -9140
rect 176923 -9174 176958 -9140
rect 177019 -9174 177207 -9140
rect 177032 -9200 177207 -9174
rect 177232 -9174 177333 -9050
rect 177110 -9870 177145 -9200
rect 177232 -9228 177235 -9174
rect 176917 -9936 177062 -9924
rect 176585 -9970 177062 -9936
rect 176917 -9971 177062 -9970
rect 177098 -9971 177145 -9870
rect 177244 -9971 177279 -9174
rect 177502 -9971 177537 -9062
rect 177636 -9971 177671 -8985
rect 177889 -9002 177924 -8968
rect 177985 -9002 178020 -8968
rect 178081 -9002 178116 -8968
rect 178177 -9002 178212 -8968
rect 178273 -9002 178308 -8968
rect 178369 -9002 178404 -8968
rect 178465 -9002 178500 -8968
rect 178974 -8992 179009 -8958
rect 179046 -8992 179081 -8958
rect 179392 -8995 179427 -8961
rect 179437 -8995 179438 -8950
rect 179579 -9001 179580 -8697
rect 180271 -8706 180306 -8672
rect 180448 -8706 180483 -8672
rect 180744 -8723 180779 -8689
rect 180789 -8723 180790 -8681
rect 180931 -8753 180932 -8525
rect 181621 -8534 181656 -8500
rect 181798 -8534 181833 -8500
rect 181992 -8577 182027 -8543
rect 182037 -8577 182038 -8532
rect 182137 -8543 182138 -8532
rect 182346 -8537 182381 -8503
rect 182391 -8537 182392 -8492
rect 182491 -8503 182492 -8492
rect 182736 -8496 182771 -8462
rect 182781 -8496 182782 -8451
rect 182881 -8462 182882 -8451
rect 182892 -8496 182927 -8462
rect 182937 -8496 182938 -8451
rect 183037 -8462 183038 -8451
rect 183218 -8456 183253 -8422
rect 183290 -8456 183325 -8422
rect 183362 -8456 183397 -8422
rect 183506 -8456 183541 -8422
rect 183578 -8456 183613 -8422
rect 183615 -8456 183685 -8422
rect 183722 -8456 183757 -8422
rect 183792 -8456 183827 -8422
rect 183048 -8496 183083 -8462
rect 184088 -8491 184123 -8457
rect 184133 -8491 184134 -8446
rect 184233 -8457 184234 -8446
rect 184244 -8491 184279 -8457
rect 184289 -8491 184290 -8446
rect 184389 -8457 184390 -8446
rect 184965 -8451 185000 -8417
rect 185142 -8451 185177 -8417
rect 184400 -8491 184435 -8457
rect 182502 -8537 182537 -8503
rect 183781 -8505 183782 -8494
rect 182148 -8577 182183 -8543
rect 181061 -8621 181096 -8587
rect 181262 -8666 181297 -8632
rect 181385 -8637 181386 -8595
rect 181707 -8624 181742 -8590
rect 182346 -8620 182381 -8586
rect 182391 -8620 182392 -8575
rect 182491 -8586 182492 -8575
rect 182736 -8580 182771 -8546
rect 182781 -8580 182782 -8535
rect 182881 -8546 182882 -8535
rect 182892 -8580 182927 -8546
rect 182937 -8580 182938 -8535
rect 183037 -8546 183038 -8535
rect 183615 -8539 183650 -8505
rect 183792 -8539 183827 -8505
rect 183048 -8580 183083 -8546
rect 183935 -8565 184050 -8499
rect 184233 -8525 184234 -8499
rect 184630 -8517 184665 -8483
rect 184675 -8517 184676 -8472
rect 184775 -8483 184776 -8472
rect 184786 -8517 184821 -8483
rect 184831 -8517 184832 -8472
rect 185131 -8500 185132 -8489
rect 185336 -8494 185371 -8460
rect 185381 -8494 185382 -8449
rect 185481 -8460 185482 -8449
rect 185690 -8453 185725 -8419
rect 185735 -8453 185736 -8408
rect 185835 -8419 185836 -8408
rect 186016 -8413 186051 -8379
rect 186080 -8413 186123 -8379
rect 186125 -8413 186126 -8371
rect 186225 -8379 186226 -8371
rect 186160 -8413 186195 -8379
rect 186236 -8413 186271 -8379
rect 186281 -8413 186282 -8371
rect 186381 -8379 186382 -8371
rect 186330 -8413 186365 -8379
rect 186392 -8413 186437 -8379
rect 187432 -8408 187467 -8374
rect 187477 -8408 187478 -8363
rect 187577 -8374 187578 -8363
rect 187588 -8408 187623 -8374
rect 187633 -8408 187634 -8363
rect 187733 -8374 187734 -8363
rect 188309 -8367 188344 -8333
rect 188486 -8367 188521 -8333
rect 189079 -8336 189080 -8328
rect 189179 -8336 189180 -8328
rect 187744 -8408 187779 -8374
rect 185846 -8453 185881 -8419
rect 187125 -8422 187126 -8414
rect 188475 -8417 188476 -8406
rect 188680 -8410 188715 -8376
rect 188725 -8410 188726 -8365
rect 188825 -8376 188826 -8365
rect 189006 -8370 189069 -8336
rect 189078 -8370 189113 -8336
rect 189190 -8370 189225 -8336
rect 189915 -8360 189950 -8326
rect 190011 -8360 190046 -8326
rect 190107 -8360 190142 -8326
rect 190203 -8360 190238 -8326
rect 190299 -8360 190334 -8326
rect 190395 -8360 190430 -8326
rect 190491 -8360 190526 -8326
rect 191819 -8333 191820 -8322
rect 191996 -8327 192059 -8293
rect 192068 -8327 192103 -8293
rect 192180 -8327 192215 -8293
rect 192711 -8317 192746 -8283
rect 192807 -8317 192842 -8283
rect 192903 -8317 192938 -8283
rect 192999 -8317 193034 -8283
rect 193095 -8317 193130 -8283
rect 194120 -8324 194155 -8290
rect 194165 -8324 194166 -8279
rect 194265 -8290 194266 -8279
rect 194276 -8324 194311 -8290
rect 194321 -8324 194322 -8279
rect 194421 -8290 194422 -8279
rect 194600 -8284 194635 -8250
rect 194672 -8284 194707 -8250
rect 194744 -8284 194779 -8250
rect 194888 -8284 194923 -8250
rect 194960 -8284 194995 -8250
rect 194997 -8284 195067 -8250
rect 195104 -8284 195139 -8250
rect 195174 -8284 195209 -8250
rect 195701 -8274 195736 -8240
rect 195797 -8274 195832 -8240
rect 195893 -8274 195928 -8240
rect 197400 -8241 197435 -8207
rect 197464 -8241 197507 -8207
rect 197509 -8241 197510 -8199
rect 197609 -8207 197610 -8199
rect 197544 -8241 197579 -8207
rect 197620 -8241 197655 -8207
rect 197665 -8241 197666 -8199
rect 197765 -8207 197766 -8199
rect 197714 -8241 197749 -8207
rect 197776 -8241 197821 -8207
rect 198691 -8231 198726 -8197
rect 198787 -8231 198822 -8197
rect 198883 -8231 198918 -8197
rect 198507 -8250 198508 -8242
rect 194432 -8324 194467 -8290
rect 195413 -8293 195414 -8285
rect 195513 -8293 195514 -8285
rect 188836 -8410 188871 -8376
rect 185492 -8494 185527 -8460
rect 182502 -8620 182537 -8586
rect 183781 -8589 183782 -8578
rect 181031 -8689 181032 -8681
rect 181042 -8723 181077 -8689
rect 181262 -8734 181297 -8700
rect 179709 -8793 179744 -8759
rect 179912 -8838 179947 -8804
rect 180035 -8809 180036 -8767
rect 180357 -8796 180392 -8762
rect 179679 -8861 179680 -8853
rect 179690 -8895 179725 -8861
rect 179912 -8906 179947 -8872
rect 179679 -8961 179680 -8950
rect 179690 -8995 179725 -8961
rect 178627 -9045 178662 -9011
rect 178723 -9045 178758 -9011
rect 178819 -9045 178854 -9011
rect 179328 -9035 179363 -9001
rect 179400 -9035 179435 -9001
rect 179472 -9035 179507 -9001
rect 179544 -9029 179580 -9001
rect 179890 -9025 179925 -8991
rect 179935 -9025 179936 -8980
rect 179544 -9035 179579 -9029
rect 178981 -9088 179016 -9054
rect 179077 -9088 179112 -9054
rect 179173 -9088 179208 -9054
rect 180077 -9076 180078 -8809
rect 180706 -8819 181093 -8753
rect 180093 -8860 180128 -8826
rect 180442 -8832 180453 -8819
rect 180376 -8874 180453 -8832
rect 180504 -8874 181093 -8819
rect 181240 -8853 181275 -8819
rect 181285 -8853 181286 -8808
rect 180376 -8877 181093 -8874
rect 180093 -8928 180128 -8894
rect 180296 -8942 180331 -8908
rect 180341 -8942 180342 -8900
rect 180177 -8991 180178 -8980
rect 180188 -9025 180223 -8991
rect 180296 -9042 180331 -9008
rect 180341 -9042 180342 -8997
rect 180189 -9078 180224 -9044
rect 180261 -9078 180296 -9044
rect 180333 -9078 180368 -9044
rect 179335 -9131 179370 -9097
rect 179431 -9131 179466 -9097
rect 179527 -9131 179562 -9097
rect 179623 -9131 179658 -9097
rect 179719 -9131 179754 -9097
rect 180376 -9114 180521 -8877
rect 180706 -8899 181093 -8877
rect 180630 -8925 181093 -8899
rect 181427 -8904 181428 -8637
rect 181443 -8688 181478 -8654
rect 182057 -8691 182092 -8657
rect 182736 -8663 182771 -8629
rect 182781 -8663 182782 -8618
rect 182881 -8629 182882 -8618
rect 182892 -8663 182927 -8629
rect 182937 -8663 182938 -8618
rect 183037 -8629 183038 -8618
rect 183615 -8623 183650 -8589
rect 183792 -8623 183827 -8589
rect 184153 -8605 184188 -8571
rect 183048 -8663 183083 -8629
rect 182881 -8697 182882 -8671
rect 183280 -8689 183315 -8655
rect 183325 -8689 183326 -8644
rect 183425 -8655 183426 -8644
rect 183436 -8689 183471 -8655
rect 183481 -8689 183482 -8644
rect 183781 -8672 183782 -8661
rect 181443 -8756 181478 -8722
rect 181646 -8770 181681 -8736
rect 181691 -8770 181692 -8728
rect 181791 -8740 181792 -8729
rect 182411 -8734 182446 -8700
rect 181802 -8774 181837 -8740
rect 181527 -8819 181528 -8808
rect 181996 -8813 182031 -8779
rect 182041 -8813 182042 -8771
rect 182141 -8779 182142 -8771
rect 182801 -8777 182836 -8743
rect 182152 -8813 182187 -8779
rect 181538 -8853 181573 -8819
rect 181646 -8870 181681 -8836
rect 181691 -8870 181692 -8825
rect 181791 -8832 181792 -8821
rect 181802 -8866 181837 -8832
rect 182350 -8856 182385 -8822
rect 182395 -8856 182396 -8814
rect 182495 -8822 182496 -8814
rect 182506 -8856 182541 -8822
rect 181539 -8906 181574 -8872
rect 181611 -8906 181646 -8872
rect 181683 -8906 181718 -8872
rect 181996 -8913 182031 -8879
rect 182041 -8913 182042 -8868
rect 182141 -8879 182142 -8868
rect 182152 -8913 182187 -8879
rect 182736 -8895 182771 -8861
rect 182781 -8895 182782 -8853
rect 180630 -8959 181106 -8925
rect 181964 -8949 181999 -8915
rect 182036 -8949 182071 -8915
rect 182350 -8956 182385 -8922
rect 182395 -8956 182396 -8911
rect 182495 -8922 182496 -8911
rect 182506 -8956 182541 -8922
rect 180630 -8985 181093 -8959
rect 180634 -8993 180835 -8985
rect 180650 -9003 180819 -8993
rect 180376 -9140 180551 -9114
rect 179883 -9174 179918 -9140
rect 179979 -9174 180014 -9140
rect 180075 -9174 180110 -9140
rect 180171 -9174 180206 -9140
rect 180267 -9174 180302 -9140
rect 180363 -9174 180551 -9140
rect 180376 -9200 180551 -9174
rect 180576 -9174 180677 -9050
rect 180454 -9870 180489 -9200
rect 180576 -9228 180579 -9174
rect 180261 -9936 180406 -9924
rect 179929 -9970 180406 -9936
rect 180261 -9971 180406 -9970
rect 180442 -9971 180489 -9870
rect 180588 -9971 180623 -9174
rect 180846 -9971 180881 -9062
rect 180980 -9971 181015 -8985
rect 181233 -9002 181268 -8968
rect 181329 -9002 181364 -8968
rect 181425 -9002 181460 -8968
rect 181521 -9002 181556 -8968
rect 181617 -9002 181652 -8968
rect 181713 -9002 181748 -8968
rect 181809 -9002 181844 -8968
rect 182318 -8992 182353 -8958
rect 182390 -8992 182425 -8958
rect 182736 -8995 182771 -8961
rect 182781 -8995 182782 -8950
rect 182923 -9001 182924 -8697
rect 183615 -8706 183650 -8672
rect 183792 -8706 183827 -8672
rect 184088 -8723 184123 -8689
rect 184133 -8723 184134 -8681
rect 184275 -8753 184276 -8525
rect 184965 -8534 185000 -8500
rect 185142 -8534 185177 -8500
rect 185336 -8577 185371 -8543
rect 185381 -8577 185382 -8532
rect 185481 -8543 185482 -8532
rect 185690 -8537 185725 -8503
rect 185735 -8537 185736 -8492
rect 185835 -8503 185836 -8492
rect 186080 -8496 186115 -8462
rect 186125 -8496 186126 -8451
rect 186225 -8462 186226 -8451
rect 186236 -8496 186271 -8462
rect 186281 -8496 186282 -8451
rect 186381 -8462 186382 -8451
rect 186562 -8456 186597 -8422
rect 186634 -8456 186669 -8422
rect 186706 -8456 186741 -8422
rect 186850 -8456 186885 -8422
rect 186922 -8456 186957 -8422
rect 186959 -8456 187029 -8422
rect 187066 -8456 187101 -8422
rect 187136 -8456 187171 -8422
rect 186392 -8496 186427 -8462
rect 187432 -8491 187467 -8457
rect 187477 -8491 187478 -8446
rect 187577 -8457 187578 -8446
rect 187588 -8491 187623 -8457
rect 187633 -8491 187634 -8446
rect 187733 -8457 187734 -8446
rect 188309 -8451 188344 -8417
rect 188486 -8451 188521 -8417
rect 187744 -8491 187779 -8457
rect 185846 -8537 185881 -8503
rect 187125 -8505 187126 -8494
rect 185492 -8577 185527 -8543
rect 184405 -8621 184440 -8587
rect 184606 -8666 184641 -8632
rect 184729 -8637 184730 -8595
rect 185051 -8624 185086 -8590
rect 185690 -8620 185725 -8586
rect 185735 -8620 185736 -8575
rect 185835 -8586 185836 -8575
rect 186080 -8580 186115 -8546
rect 186125 -8580 186126 -8535
rect 186225 -8546 186226 -8535
rect 186236 -8580 186271 -8546
rect 186281 -8580 186282 -8535
rect 186381 -8546 186382 -8535
rect 186959 -8539 186994 -8505
rect 187136 -8539 187171 -8505
rect 186392 -8580 186427 -8546
rect 187279 -8565 187394 -8499
rect 187577 -8525 187578 -8499
rect 187974 -8517 188009 -8483
rect 188019 -8517 188020 -8472
rect 188119 -8483 188120 -8472
rect 188130 -8517 188165 -8483
rect 188175 -8517 188176 -8472
rect 188475 -8500 188476 -8489
rect 188680 -8494 188715 -8460
rect 188725 -8494 188726 -8449
rect 188825 -8460 188826 -8449
rect 189034 -8453 189069 -8419
rect 189079 -8453 189080 -8408
rect 189179 -8419 189180 -8408
rect 189360 -8413 189395 -8379
rect 189424 -8413 189467 -8379
rect 189469 -8413 189470 -8371
rect 189569 -8379 189570 -8371
rect 189504 -8413 189539 -8379
rect 189580 -8413 189615 -8379
rect 189625 -8413 189626 -8371
rect 189725 -8379 189726 -8371
rect 189674 -8413 189709 -8379
rect 189736 -8413 189781 -8379
rect 190776 -8408 190811 -8374
rect 190821 -8408 190822 -8363
rect 190921 -8374 190922 -8363
rect 190932 -8408 190967 -8374
rect 190977 -8408 190978 -8363
rect 191077 -8374 191078 -8363
rect 191653 -8367 191688 -8333
rect 191830 -8367 191865 -8333
rect 192423 -8336 192424 -8328
rect 192523 -8336 192524 -8328
rect 191088 -8408 191123 -8374
rect 189190 -8453 189225 -8419
rect 190469 -8422 190470 -8414
rect 191819 -8417 191820 -8406
rect 192024 -8410 192059 -8376
rect 192069 -8410 192070 -8365
rect 192169 -8376 192170 -8365
rect 192350 -8370 192413 -8336
rect 192422 -8370 192457 -8336
rect 192534 -8370 192569 -8336
rect 193259 -8360 193294 -8326
rect 193355 -8360 193390 -8326
rect 193451 -8360 193486 -8326
rect 193547 -8360 193582 -8326
rect 193643 -8360 193678 -8326
rect 193739 -8360 193774 -8326
rect 193835 -8360 193870 -8326
rect 195163 -8333 195164 -8322
rect 195340 -8327 195403 -8293
rect 195412 -8327 195447 -8293
rect 195524 -8327 195559 -8293
rect 196055 -8317 196090 -8283
rect 196151 -8317 196186 -8283
rect 196247 -8317 196282 -8283
rect 196343 -8317 196378 -8283
rect 196439 -8317 196474 -8283
rect 197464 -8324 197499 -8290
rect 197509 -8324 197510 -8279
rect 197609 -8290 197610 -8279
rect 197620 -8324 197655 -8290
rect 197665 -8324 197666 -8279
rect 197765 -8290 197766 -8279
rect 197944 -8284 197979 -8250
rect 198016 -8284 198051 -8250
rect 198088 -8284 198123 -8250
rect 198232 -8284 198267 -8250
rect 198304 -8284 198339 -8250
rect 198341 -8284 198411 -8250
rect 198448 -8284 198483 -8250
rect 198518 -8284 198553 -8250
rect 199045 -8274 199080 -8240
rect 199141 -8274 199176 -8240
rect 199237 -8274 199272 -8240
rect 200744 -8241 200779 -8207
rect 200808 -8241 200851 -8207
rect 200853 -8241 200854 -8199
rect 200953 -8207 200954 -8199
rect 200888 -8241 200923 -8207
rect 200964 -8241 200999 -8207
rect 201009 -8241 201010 -8199
rect 201109 -8207 201110 -8199
rect 201058 -8241 201093 -8207
rect 201120 -8241 201165 -8207
rect 202035 -8231 202070 -8197
rect 202131 -8231 202166 -8197
rect 202227 -8231 202262 -8197
rect 201851 -8250 201852 -8242
rect 197776 -8324 197811 -8290
rect 198757 -8293 198758 -8285
rect 198857 -8293 198858 -8285
rect 192180 -8410 192215 -8376
rect 188836 -8494 188871 -8460
rect 185846 -8620 185881 -8586
rect 187125 -8589 187126 -8578
rect 184375 -8689 184376 -8681
rect 184386 -8723 184421 -8689
rect 184606 -8734 184641 -8700
rect 183053 -8793 183088 -8759
rect 183256 -8838 183291 -8804
rect 183379 -8809 183380 -8767
rect 183701 -8796 183736 -8762
rect 183023 -8861 183024 -8853
rect 183034 -8895 183069 -8861
rect 183256 -8906 183291 -8872
rect 183023 -8961 183024 -8950
rect 183034 -8995 183069 -8961
rect 181971 -9045 182006 -9011
rect 182067 -9045 182102 -9011
rect 182163 -9045 182198 -9011
rect 182672 -9035 182707 -9001
rect 182744 -9035 182779 -9001
rect 182816 -9035 182851 -9001
rect 182888 -9029 182924 -9001
rect 183234 -9025 183269 -8991
rect 183279 -9025 183280 -8980
rect 182888 -9035 182923 -9029
rect 182325 -9088 182360 -9054
rect 182421 -9088 182456 -9054
rect 182517 -9088 182552 -9054
rect 183421 -9076 183422 -8809
rect 184050 -8819 184437 -8753
rect 183437 -8860 183472 -8826
rect 183786 -8832 183797 -8819
rect 183720 -8874 183797 -8832
rect 183848 -8874 184437 -8819
rect 184584 -8853 184619 -8819
rect 184629 -8853 184630 -8808
rect 183720 -8877 184437 -8874
rect 183437 -8928 183472 -8894
rect 183640 -8942 183675 -8908
rect 183685 -8942 183686 -8900
rect 183521 -8991 183522 -8980
rect 183532 -9025 183567 -8991
rect 183640 -9042 183675 -9008
rect 183685 -9042 183686 -8997
rect 183533 -9078 183568 -9044
rect 183605 -9078 183640 -9044
rect 183677 -9078 183712 -9044
rect 182679 -9131 182714 -9097
rect 182775 -9131 182810 -9097
rect 182871 -9131 182906 -9097
rect 182967 -9131 183002 -9097
rect 183063 -9131 183098 -9097
rect 183720 -9114 183865 -8877
rect 184050 -8899 184437 -8877
rect 183974 -8925 184437 -8899
rect 184771 -8904 184772 -8637
rect 184787 -8688 184822 -8654
rect 185401 -8691 185436 -8657
rect 186080 -8663 186115 -8629
rect 186125 -8663 186126 -8618
rect 186225 -8629 186226 -8618
rect 186236 -8663 186271 -8629
rect 186281 -8663 186282 -8618
rect 186381 -8629 186382 -8618
rect 186959 -8623 186994 -8589
rect 187136 -8623 187171 -8589
rect 187497 -8605 187532 -8571
rect 186392 -8663 186427 -8629
rect 186225 -8697 186226 -8671
rect 186624 -8689 186659 -8655
rect 186669 -8689 186670 -8644
rect 186769 -8655 186770 -8644
rect 186780 -8689 186815 -8655
rect 186825 -8689 186826 -8644
rect 187125 -8672 187126 -8661
rect 184787 -8756 184822 -8722
rect 184990 -8770 185025 -8736
rect 185035 -8770 185036 -8728
rect 185135 -8740 185136 -8729
rect 185755 -8734 185790 -8700
rect 185146 -8774 185181 -8740
rect 184871 -8819 184872 -8808
rect 185340 -8813 185375 -8779
rect 185385 -8813 185386 -8771
rect 185485 -8779 185486 -8771
rect 186145 -8777 186180 -8743
rect 185496 -8813 185531 -8779
rect 184882 -8853 184917 -8819
rect 184990 -8870 185025 -8836
rect 185035 -8870 185036 -8825
rect 185135 -8832 185136 -8821
rect 185146 -8866 185181 -8832
rect 185694 -8856 185729 -8822
rect 185739 -8856 185740 -8814
rect 185839 -8822 185840 -8814
rect 185850 -8856 185885 -8822
rect 184883 -8906 184918 -8872
rect 184955 -8906 184990 -8872
rect 185027 -8906 185062 -8872
rect 185340 -8913 185375 -8879
rect 185385 -8913 185386 -8868
rect 185485 -8879 185486 -8868
rect 185496 -8913 185531 -8879
rect 186080 -8895 186115 -8861
rect 186125 -8895 186126 -8853
rect 183974 -8959 184450 -8925
rect 185308 -8949 185343 -8915
rect 185380 -8949 185415 -8915
rect 185694 -8956 185729 -8922
rect 185739 -8956 185740 -8911
rect 185839 -8922 185840 -8911
rect 185850 -8956 185885 -8922
rect 183974 -8985 184437 -8959
rect 183978 -8993 184179 -8985
rect 183994 -9003 184163 -8993
rect 183720 -9140 183895 -9114
rect 183227 -9174 183262 -9140
rect 183323 -9174 183358 -9140
rect 183419 -9174 183454 -9140
rect 183515 -9174 183550 -9140
rect 183611 -9174 183646 -9140
rect 183707 -9174 183895 -9140
rect 183720 -9200 183895 -9174
rect 183920 -9174 184021 -9050
rect 183798 -9870 183833 -9200
rect 183920 -9228 183923 -9174
rect 183605 -9936 183750 -9924
rect 183273 -9970 183750 -9936
rect 183605 -9971 183750 -9970
rect 183786 -9971 183833 -9870
rect 183932 -9971 183967 -9174
rect 184190 -9971 184225 -9062
rect 184324 -9971 184359 -8985
rect 184577 -9002 184612 -8968
rect 184673 -9002 184708 -8968
rect 184769 -9002 184804 -8968
rect 184865 -9002 184900 -8968
rect 184961 -9002 184996 -8968
rect 185057 -9002 185092 -8968
rect 185153 -9002 185188 -8968
rect 185662 -8992 185697 -8958
rect 185734 -8992 185769 -8958
rect 186080 -8995 186115 -8961
rect 186125 -8995 186126 -8950
rect 186267 -9001 186268 -8697
rect 186959 -8706 186994 -8672
rect 187136 -8706 187171 -8672
rect 187432 -8723 187467 -8689
rect 187477 -8723 187478 -8681
rect 187619 -8753 187620 -8525
rect 188309 -8534 188344 -8500
rect 188486 -8534 188521 -8500
rect 188680 -8577 188715 -8543
rect 188725 -8577 188726 -8532
rect 188825 -8543 188826 -8532
rect 189034 -8537 189069 -8503
rect 189079 -8537 189080 -8492
rect 189179 -8503 189180 -8492
rect 189424 -8496 189459 -8462
rect 189469 -8496 189470 -8451
rect 189569 -8462 189570 -8451
rect 189580 -8496 189615 -8462
rect 189625 -8496 189626 -8451
rect 189725 -8462 189726 -8451
rect 189906 -8456 189941 -8422
rect 189978 -8456 190013 -8422
rect 190050 -8456 190085 -8422
rect 190194 -8456 190229 -8422
rect 190266 -8456 190301 -8422
rect 190303 -8456 190373 -8422
rect 190410 -8456 190445 -8422
rect 190480 -8456 190515 -8422
rect 189736 -8496 189771 -8462
rect 190776 -8491 190811 -8457
rect 190821 -8491 190822 -8446
rect 190921 -8457 190922 -8446
rect 190932 -8491 190967 -8457
rect 190977 -8491 190978 -8446
rect 191077 -8457 191078 -8446
rect 191653 -8451 191688 -8417
rect 191830 -8451 191865 -8417
rect 191088 -8491 191123 -8457
rect 189190 -8537 189225 -8503
rect 190469 -8505 190470 -8494
rect 188836 -8577 188871 -8543
rect 187749 -8621 187784 -8587
rect 187950 -8666 187985 -8632
rect 188073 -8637 188074 -8595
rect 188395 -8624 188430 -8590
rect 189034 -8620 189069 -8586
rect 189079 -8620 189080 -8575
rect 189179 -8586 189180 -8575
rect 189424 -8580 189459 -8546
rect 189469 -8580 189470 -8535
rect 189569 -8546 189570 -8535
rect 189580 -8580 189615 -8546
rect 189625 -8580 189626 -8535
rect 189725 -8546 189726 -8535
rect 190303 -8539 190338 -8505
rect 190480 -8539 190515 -8505
rect 189736 -8580 189771 -8546
rect 190623 -8565 190738 -8499
rect 190921 -8525 190922 -8499
rect 191318 -8517 191353 -8483
rect 191363 -8517 191364 -8472
rect 191463 -8483 191464 -8472
rect 191474 -8517 191509 -8483
rect 191519 -8517 191520 -8472
rect 191819 -8500 191820 -8489
rect 192024 -8494 192059 -8460
rect 192069 -8494 192070 -8449
rect 192169 -8460 192170 -8449
rect 192378 -8453 192413 -8419
rect 192423 -8453 192424 -8408
rect 192523 -8419 192524 -8408
rect 192704 -8413 192739 -8379
rect 192768 -8413 192811 -8379
rect 192813 -8413 192814 -8371
rect 192913 -8379 192914 -8371
rect 192848 -8413 192883 -8379
rect 192924 -8413 192959 -8379
rect 192969 -8413 192970 -8371
rect 193069 -8379 193070 -8371
rect 193018 -8413 193053 -8379
rect 193080 -8413 193125 -8379
rect 194120 -8408 194155 -8374
rect 194165 -8408 194166 -8363
rect 194265 -8374 194266 -8363
rect 194276 -8408 194311 -8374
rect 194321 -8408 194322 -8363
rect 194421 -8374 194422 -8363
rect 194997 -8367 195032 -8333
rect 195174 -8367 195209 -8333
rect 195767 -8336 195768 -8328
rect 195867 -8336 195868 -8328
rect 194432 -8408 194467 -8374
rect 192534 -8453 192569 -8419
rect 193813 -8422 193814 -8414
rect 195163 -8417 195164 -8406
rect 195368 -8410 195403 -8376
rect 195413 -8410 195414 -8365
rect 195513 -8376 195514 -8365
rect 195694 -8370 195757 -8336
rect 195766 -8370 195801 -8336
rect 195878 -8370 195913 -8336
rect 196603 -8360 196638 -8326
rect 196699 -8360 196734 -8326
rect 196795 -8360 196830 -8326
rect 196891 -8360 196926 -8326
rect 196987 -8360 197022 -8326
rect 197083 -8360 197118 -8326
rect 197179 -8360 197214 -8326
rect 198507 -8333 198508 -8322
rect 198684 -8327 198747 -8293
rect 198756 -8327 198791 -8293
rect 198868 -8327 198903 -8293
rect 199399 -8317 199434 -8283
rect 199495 -8317 199530 -8283
rect 199591 -8317 199626 -8283
rect 199687 -8317 199722 -8283
rect 199783 -8317 199818 -8283
rect 200808 -8324 200843 -8290
rect 200853 -8324 200854 -8279
rect 200953 -8290 200954 -8279
rect 200964 -8324 200999 -8290
rect 201009 -8324 201010 -8279
rect 201109 -8290 201110 -8279
rect 201288 -8284 201323 -8250
rect 201360 -8284 201395 -8250
rect 201432 -8284 201467 -8250
rect 201576 -8284 201611 -8250
rect 201648 -8284 201683 -8250
rect 201685 -8284 201755 -8250
rect 201792 -8284 201827 -8250
rect 201862 -8284 201897 -8250
rect 202389 -8274 202424 -8240
rect 202485 -8274 202520 -8240
rect 202581 -8274 202616 -8240
rect 204088 -8241 204123 -8207
rect 204152 -8241 204195 -8207
rect 204197 -8241 204198 -8199
rect 204297 -8207 204298 -8199
rect 204232 -8241 204267 -8207
rect 204308 -8241 204343 -8207
rect 204353 -8241 204354 -8199
rect 204453 -8207 204454 -8199
rect 204402 -8241 204437 -8207
rect 204464 -8241 204509 -8207
rect 205379 -8231 205414 -8197
rect 205475 -8231 205510 -8197
rect 205571 -8231 205606 -8197
rect 205195 -8250 205196 -8242
rect 201120 -8324 201155 -8290
rect 202101 -8293 202102 -8285
rect 202201 -8293 202202 -8285
rect 195524 -8410 195559 -8376
rect 192180 -8494 192215 -8460
rect 189190 -8620 189225 -8586
rect 190469 -8589 190470 -8578
rect 187719 -8689 187720 -8681
rect 187730 -8723 187765 -8689
rect 187950 -8734 187985 -8700
rect 186397 -8793 186432 -8759
rect 186600 -8838 186635 -8804
rect 186723 -8809 186724 -8767
rect 187045 -8796 187080 -8762
rect 186367 -8861 186368 -8853
rect 186378 -8895 186413 -8861
rect 186600 -8906 186635 -8872
rect 186367 -8961 186368 -8950
rect 186378 -8995 186413 -8961
rect 185315 -9045 185350 -9011
rect 185411 -9045 185446 -9011
rect 185507 -9045 185542 -9011
rect 186016 -9035 186051 -9001
rect 186088 -9035 186123 -9001
rect 186160 -9035 186195 -9001
rect 186232 -9029 186268 -9001
rect 186578 -9025 186613 -8991
rect 186623 -9025 186624 -8980
rect 186232 -9035 186267 -9029
rect 185669 -9088 185704 -9054
rect 185765 -9088 185800 -9054
rect 185861 -9088 185896 -9054
rect 186765 -9076 186766 -8809
rect 187394 -8819 187781 -8753
rect 186781 -8860 186816 -8826
rect 187130 -8832 187141 -8819
rect 187064 -8874 187141 -8832
rect 187192 -8874 187781 -8819
rect 187928 -8853 187963 -8819
rect 187973 -8853 187974 -8808
rect 187064 -8877 187781 -8874
rect 186781 -8928 186816 -8894
rect 186984 -8942 187019 -8908
rect 187029 -8942 187030 -8900
rect 186865 -8991 186866 -8980
rect 186876 -9025 186911 -8991
rect 186984 -9042 187019 -9008
rect 187029 -9042 187030 -8997
rect 186877 -9078 186912 -9044
rect 186949 -9078 186984 -9044
rect 187021 -9078 187056 -9044
rect 186023 -9131 186058 -9097
rect 186119 -9131 186154 -9097
rect 186215 -9131 186250 -9097
rect 186311 -9131 186346 -9097
rect 186407 -9131 186442 -9097
rect 187064 -9114 187209 -8877
rect 187394 -8899 187781 -8877
rect 187318 -8925 187781 -8899
rect 188115 -8904 188116 -8637
rect 188131 -8688 188166 -8654
rect 188745 -8691 188780 -8657
rect 189424 -8663 189459 -8629
rect 189469 -8663 189470 -8618
rect 189569 -8629 189570 -8618
rect 189580 -8663 189615 -8629
rect 189625 -8663 189626 -8618
rect 189725 -8629 189726 -8618
rect 190303 -8623 190338 -8589
rect 190480 -8623 190515 -8589
rect 190841 -8605 190876 -8571
rect 189736 -8663 189771 -8629
rect 189569 -8697 189570 -8671
rect 189968 -8689 190003 -8655
rect 190013 -8689 190014 -8644
rect 190113 -8655 190114 -8644
rect 190124 -8689 190159 -8655
rect 190169 -8689 190170 -8644
rect 190469 -8672 190470 -8661
rect 188131 -8756 188166 -8722
rect 188334 -8770 188369 -8736
rect 188379 -8770 188380 -8728
rect 188479 -8740 188480 -8729
rect 189099 -8734 189134 -8700
rect 188490 -8774 188525 -8740
rect 188215 -8819 188216 -8808
rect 188684 -8813 188719 -8779
rect 188729 -8813 188730 -8771
rect 188829 -8779 188830 -8771
rect 189489 -8777 189524 -8743
rect 188840 -8813 188875 -8779
rect 188226 -8853 188261 -8819
rect 188334 -8870 188369 -8836
rect 188379 -8870 188380 -8825
rect 188479 -8832 188480 -8821
rect 188490 -8866 188525 -8832
rect 189038 -8856 189073 -8822
rect 189083 -8856 189084 -8814
rect 189183 -8822 189184 -8814
rect 189194 -8856 189229 -8822
rect 188227 -8906 188262 -8872
rect 188299 -8906 188334 -8872
rect 188371 -8906 188406 -8872
rect 188684 -8913 188719 -8879
rect 188729 -8913 188730 -8868
rect 188829 -8879 188830 -8868
rect 188840 -8913 188875 -8879
rect 189424 -8895 189459 -8861
rect 189469 -8895 189470 -8853
rect 187318 -8959 187794 -8925
rect 188652 -8949 188687 -8915
rect 188724 -8949 188759 -8915
rect 189038 -8956 189073 -8922
rect 189083 -8956 189084 -8911
rect 189183 -8922 189184 -8911
rect 189194 -8956 189229 -8922
rect 187318 -8985 187781 -8959
rect 187322 -8993 187523 -8985
rect 187338 -9003 187507 -8993
rect 187064 -9140 187239 -9114
rect 186571 -9174 186606 -9140
rect 186667 -9174 186702 -9140
rect 186763 -9174 186798 -9140
rect 186859 -9174 186894 -9140
rect 186955 -9174 186990 -9140
rect 187051 -9174 187239 -9140
rect 187064 -9200 187239 -9174
rect 187264 -9174 187365 -9050
rect 187142 -9870 187177 -9200
rect 187264 -9228 187267 -9174
rect 186949 -9936 187094 -9924
rect 186617 -9970 187094 -9936
rect 186949 -9971 187094 -9970
rect 187130 -9971 187177 -9870
rect 187276 -9971 187311 -9174
rect 187534 -9971 187569 -9062
rect 187668 -9971 187703 -8985
rect 187921 -9002 187956 -8968
rect 188017 -9002 188052 -8968
rect 188113 -9002 188148 -8968
rect 188209 -9002 188244 -8968
rect 188305 -9002 188340 -8968
rect 188401 -9002 188436 -8968
rect 188497 -9002 188532 -8968
rect 189006 -8992 189041 -8958
rect 189078 -8992 189113 -8958
rect 189424 -8995 189459 -8961
rect 189469 -8995 189470 -8950
rect 189611 -9001 189612 -8697
rect 190303 -8706 190338 -8672
rect 190480 -8706 190515 -8672
rect 190776 -8723 190811 -8689
rect 190821 -8723 190822 -8681
rect 190963 -8753 190964 -8525
rect 191653 -8534 191688 -8500
rect 191830 -8534 191865 -8500
rect 192024 -8577 192059 -8543
rect 192069 -8577 192070 -8532
rect 192169 -8543 192170 -8532
rect 192378 -8537 192413 -8503
rect 192423 -8537 192424 -8492
rect 192523 -8503 192524 -8492
rect 192768 -8496 192803 -8462
rect 192813 -8496 192814 -8451
rect 192913 -8462 192914 -8451
rect 192924 -8496 192959 -8462
rect 192969 -8496 192970 -8451
rect 193069 -8462 193070 -8451
rect 193250 -8456 193285 -8422
rect 193322 -8456 193357 -8422
rect 193394 -8456 193429 -8422
rect 193538 -8456 193573 -8422
rect 193610 -8456 193645 -8422
rect 193647 -8456 193717 -8422
rect 193754 -8456 193789 -8422
rect 193824 -8456 193859 -8422
rect 193080 -8496 193115 -8462
rect 194120 -8491 194155 -8457
rect 194165 -8491 194166 -8446
rect 194265 -8457 194266 -8446
rect 194276 -8491 194311 -8457
rect 194321 -8491 194322 -8446
rect 194421 -8457 194422 -8446
rect 194997 -8451 195032 -8417
rect 195174 -8451 195209 -8417
rect 194432 -8491 194467 -8457
rect 192534 -8537 192569 -8503
rect 193813 -8505 193814 -8494
rect 192180 -8577 192215 -8543
rect 191093 -8621 191128 -8587
rect 191294 -8666 191329 -8632
rect 191417 -8637 191418 -8595
rect 191739 -8624 191774 -8590
rect 192378 -8620 192413 -8586
rect 192423 -8620 192424 -8575
rect 192523 -8586 192524 -8575
rect 192768 -8580 192803 -8546
rect 192813 -8580 192814 -8535
rect 192913 -8546 192914 -8535
rect 192924 -8580 192959 -8546
rect 192969 -8580 192970 -8535
rect 193069 -8546 193070 -8535
rect 193647 -8539 193682 -8505
rect 193824 -8539 193859 -8505
rect 193080 -8580 193115 -8546
rect 193967 -8565 194082 -8499
rect 194265 -8525 194266 -8499
rect 194662 -8517 194697 -8483
rect 194707 -8517 194708 -8472
rect 194807 -8483 194808 -8472
rect 194818 -8517 194853 -8483
rect 194863 -8517 194864 -8472
rect 195163 -8500 195164 -8489
rect 195368 -8494 195403 -8460
rect 195413 -8494 195414 -8449
rect 195513 -8460 195514 -8449
rect 195722 -8453 195757 -8419
rect 195767 -8453 195768 -8408
rect 195867 -8419 195868 -8408
rect 196048 -8413 196083 -8379
rect 196112 -8413 196155 -8379
rect 196157 -8413 196158 -8371
rect 196257 -8379 196258 -8371
rect 196192 -8413 196227 -8379
rect 196268 -8413 196303 -8379
rect 196313 -8413 196314 -8371
rect 196413 -8379 196414 -8371
rect 196362 -8413 196397 -8379
rect 196424 -8413 196469 -8379
rect 197464 -8408 197499 -8374
rect 197509 -8408 197510 -8363
rect 197609 -8374 197610 -8363
rect 197620 -8408 197655 -8374
rect 197665 -8408 197666 -8363
rect 197765 -8374 197766 -8363
rect 198341 -8367 198376 -8333
rect 198518 -8367 198553 -8333
rect 199111 -8336 199112 -8328
rect 199211 -8336 199212 -8328
rect 197776 -8408 197811 -8374
rect 195878 -8453 195913 -8419
rect 197157 -8422 197158 -8414
rect 198507 -8417 198508 -8406
rect 198712 -8410 198747 -8376
rect 198757 -8410 198758 -8365
rect 198857 -8376 198858 -8365
rect 199038 -8370 199101 -8336
rect 199110 -8370 199145 -8336
rect 199222 -8370 199257 -8336
rect 199947 -8360 199982 -8326
rect 200043 -8360 200078 -8326
rect 200139 -8360 200174 -8326
rect 200235 -8360 200270 -8326
rect 200331 -8360 200366 -8326
rect 200427 -8360 200462 -8326
rect 200523 -8360 200558 -8326
rect 201851 -8333 201852 -8322
rect 202028 -8327 202091 -8293
rect 202100 -8327 202135 -8293
rect 202212 -8327 202247 -8293
rect 202743 -8317 202778 -8283
rect 202839 -8317 202874 -8283
rect 202935 -8317 202970 -8283
rect 203031 -8317 203066 -8283
rect 203127 -8317 203162 -8283
rect 204152 -8324 204187 -8290
rect 204197 -8324 204198 -8279
rect 204297 -8290 204298 -8279
rect 204308 -8324 204343 -8290
rect 204353 -8324 204354 -8279
rect 204453 -8290 204454 -8279
rect 204632 -8284 204667 -8250
rect 204704 -8284 204739 -8250
rect 204776 -8284 204811 -8250
rect 204920 -8284 204955 -8250
rect 204992 -8284 205027 -8250
rect 205029 -8284 205099 -8250
rect 205136 -8284 205171 -8250
rect 205206 -8284 205241 -8250
rect 205733 -8274 205768 -8240
rect 205829 -8274 205864 -8240
rect 205925 -8274 205960 -8240
rect 207432 -8241 207467 -8207
rect 207496 -8241 207539 -8207
rect 207541 -8241 207542 -8199
rect 207641 -8207 207642 -8199
rect 207576 -8241 207611 -8207
rect 207652 -8241 207687 -8207
rect 207697 -8241 207698 -8199
rect 207797 -8207 207798 -8199
rect 207746 -8241 207781 -8207
rect 207808 -8241 207853 -8207
rect 208723 -8231 208758 -8197
rect 208819 -8231 208854 -8197
rect 208915 -8231 208950 -8197
rect 208539 -8250 208540 -8242
rect 204464 -8324 204499 -8290
rect 205445 -8293 205446 -8285
rect 205545 -8293 205546 -8285
rect 198868 -8410 198903 -8376
rect 195524 -8494 195559 -8460
rect 192534 -8620 192569 -8586
rect 193813 -8589 193814 -8578
rect 191063 -8689 191064 -8681
rect 191074 -8723 191109 -8689
rect 191294 -8734 191329 -8700
rect 189741 -8793 189776 -8759
rect 189944 -8838 189979 -8804
rect 190067 -8809 190068 -8767
rect 190389 -8796 190424 -8762
rect 189711 -8861 189712 -8853
rect 189722 -8895 189757 -8861
rect 189944 -8906 189979 -8872
rect 189711 -8961 189712 -8950
rect 189722 -8995 189757 -8961
rect 188659 -9045 188694 -9011
rect 188755 -9045 188790 -9011
rect 188851 -9045 188886 -9011
rect 189360 -9035 189395 -9001
rect 189432 -9035 189467 -9001
rect 189504 -9035 189539 -9001
rect 189576 -9029 189612 -9001
rect 189922 -9025 189957 -8991
rect 189967 -9025 189968 -8980
rect 189576 -9035 189611 -9029
rect 189013 -9088 189048 -9054
rect 189109 -9088 189144 -9054
rect 189205 -9088 189240 -9054
rect 190109 -9076 190110 -8809
rect 190738 -8819 191125 -8753
rect 190125 -8860 190160 -8826
rect 190474 -8832 190485 -8819
rect 190408 -8874 190485 -8832
rect 190536 -8874 191125 -8819
rect 191272 -8853 191307 -8819
rect 191317 -8853 191318 -8808
rect 190408 -8877 191125 -8874
rect 190125 -8928 190160 -8894
rect 190328 -8942 190363 -8908
rect 190373 -8942 190374 -8900
rect 190209 -8991 190210 -8980
rect 190220 -9025 190255 -8991
rect 190328 -9042 190363 -9008
rect 190373 -9042 190374 -8997
rect 190221 -9078 190256 -9044
rect 190293 -9078 190328 -9044
rect 190365 -9078 190400 -9044
rect 189367 -9131 189402 -9097
rect 189463 -9131 189498 -9097
rect 189559 -9131 189594 -9097
rect 189655 -9131 189690 -9097
rect 189751 -9131 189786 -9097
rect 190408 -9114 190553 -8877
rect 190738 -8899 191125 -8877
rect 190662 -8925 191125 -8899
rect 191459 -8904 191460 -8637
rect 191475 -8688 191510 -8654
rect 192089 -8691 192124 -8657
rect 192768 -8663 192803 -8629
rect 192813 -8663 192814 -8618
rect 192913 -8629 192914 -8618
rect 192924 -8663 192959 -8629
rect 192969 -8663 192970 -8618
rect 193069 -8629 193070 -8618
rect 193647 -8623 193682 -8589
rect 193824 -8623 193859 -8589
rect 194185 -8605 194220 -8571
rect 193080 -8663 193115 -8629
rect 192913 -8697 192914 -8671
rect 193312 -8689 193347 -8655
rect 193357 -8689 193358 -8644
rect 193457 -8655 193458 -8644
rect 193468 -8689 193503 -8655
rect 193513 -8689 193514 -8644
rect 193813 -8672 193814 -8661
rect 191475 -8756 191510 -8722
rect 191678 -8770 191713 -8736
rect 191723 -8770 191724 -8728
rect 191823 -8740 191824 -8729
rect 192443 -8734 192478 -8700
rect 191834 -8774 191869 -8740
rect 191559 -8819 191560 -8808
rect 192028 -8813 192063 -8779
rect 192073 -8813 192074 -8771
rect 192173 -8779 192174 -8771
rect 192833 -8777 192868 -8743
rect 192184 -8813 192219 -8779
rect 191570 -8853 191605 -8819
rect 191678 -8870 191713 -8836
rect 191723 -8870 191724 -8825
rect 191823 -8832 191824 -8821
rect 191834 -8866 191869 -8832
rect 192382 -8856 192417 -8822
rect 192427 -8856 192428 -8814
rect 192527 -8822 192528 -8814
rect 192538 -8856 192573 -8822
rect 191571 -8906 191606 -8872
rect 191643 -8906 191678 -8872
rect 191715 -8906 191750 -8872
rect 192028 -8913 192063 -8879
rect 192073 -8913 192074 -8868
rect 192173 -8879 192174 -8868
rect 192184 -8913 192219 -8879
rect 192768 -8895 192803 -8861
rect 192813 -8895 192814 -8853
rect 190662 -8959 191138 -8925
rect 191996 -8949 192031 -8915
rect 192068 -8949 192103 -8915
rect 192382 -8956 192417 -8922
rect 192427 -8956 192428 -8911
rect 192527 -8922 192528 -8911
rect 192538 -8956 192573 -8922
rect 190662 -8985 191125 -8959
rect 190666 -8993 190867 -8985
rect 190682 -9003 190851 -8993
rect 190408 -9140 190583 -9114
rect 189915 -9174 189950 -9140
rect 190011 -9174 190046 -9140
rect 190107 -9174 190142 -9140
rect 190203 -9174 190238 -9140
rect 190299 -9174 190334 -9140
rect 190395 -9174 190583 -9140
rect 190408 -9200 190583 -9174
rect 190608 -9174 190709 -9050
rect 190486 -9870 190521 -9200
rect 190608 -9228 190611 -9174
rect 190293 -9936 190438 -9924
rect 189961 -9970 190438 -9936
rect 190293 -9971 190438 -9970
rect 190474 -9971 190521 -9870
rect 190620 -9971 190655 -9174
rect 190878 -9971 190913 -9062
rect 191012 -9971 191047 -8985
rect 191265 -9002 191300 -8968
rect 191361 -9002 191396 -8968
rect 191457 -9002 191492 -8968
rect 191553 -9002 191588 -8968
rect 191649 -9002 191684 -8968
rect 191745 -9002 191780 -8968
rect 191841 -9002 191876 -8968
rect 192350 -8992 192385 -8958
rect 192422 -8992 192457 -8958
rect 192768 -8995 192803 -8961
rect 192813 -8995 192814 -8950
rect 192955 -9001 192956 -8697
rect 193647 -8706 193682 -8672
rect 193824 -8706 193859 -8672
rect 194120 -8723 194155 -8689
rect 194165 -8723 194166 -8681
rect 194307 -8753 194308 -8525
rect 194997 -8534 195032 -8500
rect 195174 -8534 195209 -8500
rect 195368 -8577 195403 -8543
rect 195413 -8577 195414 -8532
rect 195513 -8543 195514 -8532
rect 195722 -8537 195757 -8503
rect 195767 -8537 195768 -8492
rect 195867 -8503 195868 -8492
rect 196112 -8496 196147 -8462
rect 196157 -8496 196158 -8451
rect 196257 -8462 196258 -8451
rect 196268 -8496 196303 -8462
rect 196313 -8496 196314 -8451
rect 196413 -8462 196414 -8451
rect 196594 -8456 196629 -8422
rect 196666 -8456 196701 -8422
rect 196738 -8456 196773 -8422
rect 196882 -8456 196917 -8422
rect 196954 -8456 196989 -8422
rect 196991 -8456 197061 -8422
rect 197098 -8456 197133 -8422
rect 197168 -8456 197203 -8422
rect 196424 -8496 196459 -8462
rect 197464 -8491 197499 -8457
rect 197509 -8491 197510 -8446
rect 197609 -8457 197610 -8446
rect 197620 -8491 197655 -8457
rect 197665 -8491 197666 -8446
rect 197765 -8457 197766 -8446
rect 198341 -8451 198376 -8417
rect 198518 -8451 198553 -8417
rect 197776 -8491 197811 -8457
rect 195878 -8537 195913 -8503
rect 197157 -8505 197158 -8494
rect 195524 -8577 195559 -8543
rect 194437 -8621 194472 -8587
rect 194638 -8666 194673 -8632
rect 194761 -8637 194762 -8595
rect 195083 -8624 195118 -8590
rect 195722 -8620 195757 -8586
rect 195767 -8620 195768 -8575
rect 195867 -8586 195868 -8575
rect 196112 -8580 196147 -8546
rect 196157 -8580 196158 -8535
rect 196257 -8546 196258 -8535
rect 196268 -8580 196303 -8546
rect 196313 -8580 196314 -8535
rect 196413 -8546 196414 -8535
rect 196991 -8539 197026 -8505
rect 197168 -8539 197203 -8505
rect 196424 -8580 196459 -8546
rect 197311 -8565 197426 -8499
rect 197609 -8525 197610 -8499
rect 198006 -8517 198041 -8483
rect 198051 -8517 198052 -8472
rect 198151 -8483 198152 -8472
rect 198162 -8517 198197 -8483
rect 198207 -8517 198208 -8472
rect 198507 -8500 198508 -8489
rect 198712 -8494 198747 -8460
rect 198757 -8494 198758 -8449
rect 198857 -8460 198858 -8449
rect 199066 -8453 199101 -8419
rect 199111 -8453 199112 -8408
rect 199211 -8419 199212 -8408
rect 199392 -8413 199427 -8379
rect 199456 -8413 199499 -8379
rect 199501 -8413 199502 -8371
rect 199601 -8379 199602 -8371
rect 199536 -8413 199571 -8379
rect 199612 -8413 199647 -8379
rect 199657 -8413 199658 -8371
rect 199757 -8379 199758 -8371
rect 199706 -8413 199741 -8379
rect 199768 -8413 199813 -8379
rect 200808 -8408 200843 -8374
rect 200853 -8408 200854 -8363
rect 200953 -8374 200954 -8363
rect 200964 -8408 200999 -8374
rect 201009 -8408 201010 -8363
rect 201109 -8374 201110 -8363
rect 201685 -8367 201720 -8333
rect 201862 -8367 201897 -8333
rect 202455 -8336 202456 -8328
rect 202555 -8336 202556 -8328
rect 201120 -8408 201155 -8374
rect 199222 -8453 199257 -8419
rect 200501 -8422 200502 -8414
rect 201851 -8417 201852 -8406
rect 202056 -8410 202091 -8376
rect 202101 -8410 202102 -8365
rect 202201 -8376 202202 -8365
rect 202382 -8370 202445 -8336
rect 202454 -8370 202489 -8336
rect 202566 -8370 202601 -8336
rect 203291 -8360 203326 -8326
rect 203387 -8360 203422 -8326
rect 203483 -8360 203518 -8326
rect 203579 -8360 203614 -8326
rect 203675 -8360 203710 -8326
rect 203771 -8360 203806 -8326
rect 203867 -8360 203902 -8326
rect 205195 -8333 205196 -8322
rect 205372 -8327 205435 -8293
rect 205444 -8327 205479 -8293
rect 205556 -8327 205591 -8293
rect 206087 -8317 206122 -8283
rect 206183 -8317 206218 -8283
rect 206279 -8317 206314 -8283
rect 206375 -8317 206410 -8283
rect 206471 -8317 206506 -8283
rect 207496 -8324 207531 -8290
rect 207541 -8324 207542 -8279
rect 207641 -8290 207642 -8279
rect 207652 -8324 207687 -8290
rect 207697 -8324 207698 -8279
rect 207797 -8290 207798 -8279
rect 207976 -8284 208011 -8250
rect 208048 -8284 208083 -8250
rect 208120 -8284 208155 -8250
rect 208264 -8284 208299 -8250
rect 208336 -8284 208371 -8250
rect 208373 -8284 208443 -8250
rect 208480 -8284 208515 -8250
rect 208550 -8284 208585 -8250
rect 209077 -8274 209112 -8240
rect 209173 -8274 209208 -8240
rect 209269 -8274 209304 -8240
rect 210776 -8241 210811 -8207
rect 210840 -8241 210883 -8207
rect 210885 -8241 210886 -8199
rect 210985 -8207 210986 -8199
rect 210920 -8241 210955 -8207
rect 210996 -8241 211031 -8207
rect 211041 -8241 211042 -8199
rect 211141 -8207 211142 -8199
rect 211090 -8241 211125 -8207
rect 211152 -8241 211197 -8207
rect 212067 -8231 212102 -8197
rect 212163 -8231 212198 -8197
rect 212259 -8231 212294 -8197
rect 211883 -8250 211884 -8242
rect 207808 -8324 207843 -8290
rect 208789 -8293 208790 -8285
rect 208889 -8293 208890 -8285
rect 202212 -8410 202247 -8376
rect 198868 -8494 198903 -8460
rect 195878 -8620 195913 -8586
rect 197157 -8589 197158 -8578
rect 194407 -8689 194408 -8681
rect 194418 -8723 194453 -8689
rect 194638 -8734 194673 -8700
rect 193085 -8793 193120 -8759
rect 193288 -8838 193323 -8804
rect 193411 -8809 193412 -8767
rect 193733 -8796 193768 -8762
rect 193055 -8861 193056 -8853
rect 193066 -8895 193101 -8861
rect 193288 -8906 193323 -8872
rect 193055 -8961 193056 -8950
rect 193066 -8995 193101 -8961
rect 192003 -9045 192038 -9011
rect 192099 -9045 192134 -9011
rect 192195 -9045 192230 -9011
rect 192704 -9035 192739 -9001
rect 192776 -9035 192811 -9001
rect 192848 -9035 192883 -9001
rect 192920 -9029 192956 -9001
rect 193266 -9025 193301 -8991
rect 193311 -9025 193312 -8980
rect 192920 -9035 192955 -9029
rect 192357 -9088 192392 -9054
rect 192453 -9088 192488 -9054
rect 192549 -9088 192584 -9054
rect 193453 -9076 193454 -8809
rect 194082 -8819 194469 -8753
rect 193469 -8860 193504 -8826
rect 193818 -8832 193829 -8819
rect 193752 -8874 193829 -8832
rect 193880 -8874 194469 -8819
rect 194616 -8853 194651 -8819
rect 194661 -8853 194662 -8808
rect 193752 -8877 194469 -8874
rect 193469 -8928 193504 -8894
rect 193672 -8942 193707 -8908
rect 193717 -8942 193718 -8900
rect 193553 -8991 193554 -8980
rect 193564 -9025 193599 -8991
rect 193672 -9042 193707 -9008
rect 193717 -9042 193718 -8997
rect 193565 -9078 193600 -9044
rect 193637 -9078 193672 -9044
rect 193709 -9078 193744 -9044
rect 192711 -9131 192746 -9097
rect 192807 -9131 192842 -9097
rect 192903 -9131 192938 -9097
rect 192999 -9131 193034 -9097
rect 193095 -9131 193130 -9097
rect 193752 -9114 193897 -8877
rect 194082 -8899 194469 -8877
rect 194006 -8925 194469 -8899
rect 194803 -8904 194804 -8637
rect 194819 -8688 194854 -8654
rect 195433 -8691 195468 -8657
rect 196112 -8663 196147 -8629
rect 196157 -8663 196158 -8618
rect 196257 -8629 196258 -8618
rect 196268 -8663 196303 -8629
rect 196313 -8663 196314 -8618
rect 196413 -8629 196414 -8618
rect 196991 -8623 197026 -8589
rect 197168 -8623 197203 -8589
rect 197529 -8605 197564 -8571
rect 196424 -8663 196459 -8629
rect 196257 -8697 196258 -8671
rect 196656 -8689 196691 -8655
rect 196701 -8689 196702 -8644
rect 196801 -8655 196802 -8644
rect 196812 -8689 196847 -8655
rect 196857 -8689 196858 -8644
rect 197157 -8672 197158 -8661
rect 194819 -8756 194854 -8722
rect 195022 -8770 195057 -8736
rect 195067 -8770 195068 -8728
rect 195167 -8740 195168 -8729
rect 195787 -8734 195822 -8700
rect 195178 -8774 195213 -8740
rect 194903 -8819 194904 -8808
rect 195372 -8813 195407 -8779
rect 195417 -8813 195418 -8771
rect 195517 -8779 195518 -8771
rect 196177 -8777 196212 -8743
rect 195528 -8813 195563 -8779
rect 194914 -8853 194949 -8819
rect 195022 -8870 195057 -8836
rect 195067 -8870 195068 -8825
rect 195167 -8832 195168 -8821
rect 195178 -8866 195213 -8832
rect 195726 -8856 195761 -8822
rect 195771 -8856 195772 -8814
rect 195871 -8822 195872 -8814
rect 195882 -8856 195917 -8822
rect 194915 -8906 194950 -8872
rect 194987 -8906 195022 -8872
rect 195059 -8906 195094 -8872
rect 195372 -8913 195407 -8879
rect 195417 -8913 195418 -8868
rect 195517 -8879 195518 -8868
rect 195528 -8913 195563 -8879
rect 196112 -8895 196147 -8861
rect 196157 -8895 196158 -8853
rect 194006 -8959 194482 -8925
rect 195340 -8949 195375 -8915
rect 195412 -8949 195447 -8915
rect 195726 -8956 195761 -8922
rect 195771 -8956 195772 -8911
rect 195871 -8922 195872 -8911
rect 195882 -8956 195917 -8922
rect 194006 -8985 194469 -8959
rect 194010 -8993 194211 -8985
rect 194026 -9003 194195 -8993
rect 193752 -9140 193927 -9114
rect 193259 -9174 193294 -9140
rect 193355 -9174 193390 -9140
rect 193451 -9174 193486 -9140
rect 193547 -9174 193582 -9140
rect 193643 -9174 193678 -9140
rect 193739 -9174 193927 -9140
rect 193752 -9200 193927 -9174
rect 193952 -9174 194053 -9050
rect 193830 -9870 193865 -9200
rect 193952 -9228 193955 -9174
rect 193637 -9936 193782 -9924
rect 193305 -9970 193782 -9936
rect 193637 -9971 193782 -9970
rect 193818 -9971 193865 -9870
rect 193964 -9971 193999 -9174
rect 194222 -9971 194257 -9062
rect 194356 -9971 194391 -8985
rect 194609 -9002 194644 -8968
rect 194705 -9002 194740 -8968
rect 194801 -9002 194836 -8968
rect 194897 -9002 194932 -8968
rect 194993 -9002 195028 -8968
rect 195089 -9002 195124 -8968
rect 195185 -9002 195220 -8968
rect 195694 -8992 195729 -8958
rect 195766 -8992 195801 -8958
rect 196112 -8995 196147 -8961
rect 196157 -8995 196158 -8950
rect 196299 -9001 196300 -8697
rect 196991 -8706 197026 -8672
rect 197168 -8706 197203 -8672
rect 197464 -8723 197499 -8689
rect 197509 -8723 197510 -8681
rect 197651 -8753 197652 -8525
rect 198341 -8534 198376 -8500
rect 198518 -8534 198553 -8500
rect 198712 -8577 198747 -8543
rect 198757 -8577 198758 -8532
rect 198857 -8543 198858 -8532
rect 199066 -8537 199101 -8503
rect 199111 -8537 199112 -8492
rect 199211 -8503 199212 -8492
rect 199456 -8496 199491 -8462
rect 199501 -8496 199502 -8451
rect 199601 -8462 199602 -8451
rect 199612 -8496 199647 -8462
rect 199657 -8496 199658 -8451
rect 199757 -8462 199758 -8451
rect 199938 -8456 199973 -8422
rect 200010 -8456 200045 -8422
rect 200082 -8456 200117 -8422
rect 200226 -8456 200261 -8422
rect 200298 -8456 200333 -8422
rect 200335 -8456 200405 -8422
rect 200442 -8456 200477 -8422
rect 200512 -8456 200547 -8422
rect 199768 -8496 199803 -8462
rect 200808 -8491 200843 -8457
rect 200853 -8491 200854 -8446
rect 200953 -8457 200954 -8446
rect 200964 -8491 200999 -8457
rect 201009 -8491 201010 -8446
rect 201109 -8457 201110 -8446
rect 201685 -8451 201720 -8417
rect 201862 -8451 201897 -8417
rect 201120 -8491 201155 -8457
rect 199222 -8537 199257 -8503
rect 200501 -8505 200502 -8494
rect 198868 -8577 198903 -8543
rect 197781 -8621 197816 -8587
rect 197982 -8666 198017 -8632
rect 198105 -8637 198106 -8595
rect 198427 -8624 198462 -8590
rect 199066 -8620 199101 -8586
rect 199111 -8620 199112 -8575
rect 199211 -8586 199212 -8575
rect 199456 -8580 199491 -8546
rect 199501 -8580 199502 -8535
rect 199601 -8546 199602 -8535
rect 199612 -8580 199647 -8546
rect 199657 -8580 199658 -8535
rect 199757 -8546 199758 -8535
rect 200335 -8539 200370 -8505
rect 200512 -8539 200547 -8505
rect 199768 -8580 199803 -8546
rect 200655 -8565 200770 -8499
rect 200953 -8525 200954 -8499
rect 201350 -8517 201385 -8483
rect 201395 -8517 201396 -8472
rect 201495 -8483 201496 -8472
rect 201506 -8517 201541 -8483
rect 201551 -8517 201552 -8472
rect 201851 -8500 201852 -8489
rect 202056 -8494 202091 -8460
rect 202101 -8494 202102 -8449
rect 202201 -8460 202202 -8449
rect 202410 -8453 202445 -8419
rect 202455 -8453 202456 -8408
rect 202555 -8419 202556 -8408
rect 202736 -8413 202771 -8379
rect 202800 -8413 202843 -8379
rect 202845 -8413 202846 -8371
rect 202945 -8379 202946 -8371
rect 202880 -8413 202915 -8379
rect 202956 -8413 202991 -8379
rect 203001 -8413 203002 -8371
rect 203101 -8379 203102 -8371
rect 203050 -8413 203085 -8379
rect 203112 -8413 203157 -8379
rect 204152 -8408 204187 -8374
rect 204197 -8408 204198 -8363
rect 204297 -8374 204298 -8363
rect 204308 -8408 204343 -8374
rect 204353 -8408 204354 -8363
rect 204453 -8374 204454 -8363
rect 205029 -8367 205064 -8333
rect 205206 -8367 205241 -8333
rect 205799 -8336 205800 -8328
rect 205899 -8336 205900 -8328
rect 204464 -8408 204499 -8374
rect 202566 -8453 202601 -8419
rect 203845 -8422 203846 -8414
rect 205195 -8417 205196 -8406
rect 205400 -8410 205435 -8376
rect 205445 -8410 205446 -8365
rect 205545 -8376 205546 -8365
rect 205726 -8370 205789 -8336
rect 205798 -8370 205833 -8336
rect 205910 -8370 205945 -8336
rect 206635 -8360 206670 -8326
rect 206731 -8360 206766 -8326
rect 206827 -8360 206862 -8326
rect 206923 -8360 206958 -8326
rect 207019 -8360 207054 -8326
rect 207115 -8360 207150 -8326
rect 207211 -8360 207246 -8326
rect 208539 -8333 208540 -8322
rect 208716 -8327 208779 -8293
rect 208788 -8327 208823 -8293
rect 208900 -8327 208935 -8293
rect 209431 -8317 209466 -8283
rect 209527 -8317 209562 -8283
rect 209623 -8317 209658 -8283
rect 209719 -8317 209754 -8283
rect 209815 -8317 209850 -8283
rect 210840 -8324 210875 -8290
rect 210885 -8324 210886 -8279
rect 210985 -8290 210986 -8279
rect 210996 -8324 211031 -8290
rect 211041 -8324 211042 -8279
rect 211141 -8290 211142 -8279
rect 211320 -8284 211355 -8250
rect 211392 -8284 211427 -8250
rect 211464 -8284 211499 -8250
rect 211608 -8284 211643 -8250
rect 211680 -8284 211715 -8250
rect 211717 -8284 211787 -8250
rect 211824 -8284 211859 -8250
rect 211894 -8284 211929 -8250
rect 212421 -8274 212456 -8240
rect 212517 -8274 212552 -8240
rect 212613 -8274 212648 -8240
rect 211152 -8324 211187 -8290
rect 212133 -8293 212134 -8285
rect 212233 -8293 212234 -8285
rect 205556 -8410 205591 -8376
rect 202212 -8494 202247 -8460
rect 199222 -8620 199257 -8586
rect 200501 -8589 200502 -8578
rect 197751 -8689 197752 -8681
rect 197762 -8723 197797 -8689
rect 197982 -8734 198017 -8700
rect 196429 -8793 196464 -8759
rect 196632 -8838 196667 -8804
rect 196755 -8809 196756 -8767
rect 197077 -8796 197112 -8762
rect 196399 -8861 196400 -8853
rect 196410 -8895 196445 -8861
rect 196632 -8906 196667 -8872
rect 196399 -8961 196400 -8950
rect 196410 -8995 196445 -8961
rect 195347 -9045 195382 -9011
rect 195443 -9045 195478 -9011
rect 195539 -9045 195574 -9011
rect 196048 -9035 196083 -9001
rect 196120 -9035 196155 -9001
rect 196192 -9035 196227 -9001
rect 196264 -9029 196300 -9001
rect 196610 -9025 196645 -8991
rect 196655 -9025 196656 -8980
rect 196264 -9035 196299 -9029
rect 195701 -9088 195736 -9054
rect 195797 -9088 195832 -9054
rect 195893 -9088 195928 -9054
rect 196797 -9076 196798 -8809
rect 197426 -8819 197813 -8753
rect 196813 -8860 196848 -8826
rect 197162 -8832 197173 -8819
rect 197096 -8874 197173 -8832
rect 197224 -8874 197813 -8819
rect 197960 -8853 197995 -8819
rect 198005 -8853 198006 -8808
rect 197096 -8877 197813 -8874
rect 196813 -8928 196848 -8894
rect 197016 -8942 197051 -8908
rect 197061 -8942 197062 -8900
rect 196897 -8991 196898 -8980
rect 196908 -9025 196943 -8991
rect 197016 -9042 197051 -9008
rect 197061 -9042 197062 -8997
rect 196909 -9078 196944 -9044
rect 196981 -9078 197016 -9044
rect 197053 -9078 197088 -9044
rect 196055 -9131 196090 -9097
rect 196151 -9131 196186 -9097
rect 196247 -9131 196282 -9097
rect 196343 -9131 196378 -9097
rect 196439 -9131 196474 -9097
rect 197096 -9114 197241 -8877
rect 197426 -8899 197813 -8877
rect 197350 -8925 197813 -8899
rect 198147 -8904 198148 -8637
rect 198163 -8688 198198 -8654
rect 198777 -8691 198812 -8657
rect 199456 -8663 199491 -8629
rect 199501 -8663 199502 -8618
rect 199601 -8629 199602 -8618
rect 199612 -8663 199647 -8629
rect 199657 -8663 199658 -8618
rect 199757 -8629 199758 -8618
rect 200335 -8623 200370 -8589
rect 200512 -8623 200547 -8589
rect 200873 -8605 200908 -8571
rect 199768 -8663 199803 -8629
rect 199601 -8697 199602 -8671
rect 200000 -8689 200035 -8655
rect 200045 -8689 200046 -8644
rect 200145 -8655 200146 -8644
rect 200156 -8689 200191 -8655
rect 200201 -8689 200202 -8644
rect 200501 -8672 200502 -8661
rect 198163 -8756 198198 -8722
rect 198366 -8770 198401 -8736
rect 198411 -8770 198412 -8728
rect 198511 -8740 198512 -8729
rect 199131 -8734 199166 -8700
rect 198522 -8774 198557 -8740
rect 198247 -8819 198248 -8808
rect 198716 -8813 198751 -8779
rect 198761 -8813 198762 -8771
rect 198861 -8779 198862 -8771
rect 199521 -8777 199556 -8743
rect 198872 -8813 198907 -8779
rect 198258 -8853 198293 -8819
rect 198366 -8870 198401 -8836
rect 198411 -8870 198412 -8825
rect 198511 -8832 198512 -8821
rect 198522 -8866 198557 -8832
rect 199070 -8856 199105 -8822
rect 199115 -8856 199116 -8814
rect 199215 -8822 199216 -8814
rect 199226 -8856 199261 -8822
rect 198259 -8906 198294 -8872
rect 198331 -8906 198366 -8872
rect 198403 -8906 198438 -8872
rect 198716 -8913 198751 -8879
rect 198761 -8913 198762 -8868
rect 198861 -8879 198862 -8868
rect 198872 -8913 198907 -8879
rect 199456 -8895 199491 -8861
rect 199501 -8895 199502 -8853
rect 197350 -8959 197826 -8925
rect 198684 -8949 198719 -8915
rect 198756 -8949 198791 -8915
rect 199070 -8956 199105 -8922
rect 199115 -8956 199116 -8911
rect 199215 -8922 199216 -8911
rect 199226 -8956 199261 -8922
rect 197350 -8985 197813 -8959
rect 197354 -8993 197555 -8985
rect 197370 -9003 197539 -8993
rect 197096 -9140 197271 -9114
rect 196603 -9174 196638 -9140
rect 196699 -9174 196734 -9140
rect 196795 -9174 196830 -9140
rect 196891 -9174 196926 -9140
rect 196987 -9174 197022 -9140
rect 197083 -9174 197271 -9140
rect 197096 -9200 197271 -9174
rect 197296 -9174 197397 -9050
rect 197174 -9870 197209 -9200
rect 197296 -9228 197299 -9174
rect 196981 -9936 197126 -9924
rect 196649 -9970 197126 -9936
rect 196981 -9971 197126 -9970
rect 197162 -9971 197209 -9870
rect 197308 -9971 197343 -9174
rect 197566 -9971 197601 -9062
rect 197700 -9971 197735 -8985
rect 197953 -9002 197988 -8968
rect 198049 -9002 198084 -8968
rect 198145 -9002 198180 -8968
rect 198241 -9002 198276 -8968
rect 198337 -9002 198372 -8968
rect 198433 -9002 198468 -8968
rect 198529 -9002 198564 -8968
rect 199038 -8992 199073 -8958
rect 199110 -8992 199145 -8958
rect 199456 -8995 199491 -8961
rect 199501 -8995 199502 -8950
rect 199643 -9001 199644 -8697
rect 200335 -8706 200370 -8672
rect 200512 -8706 200547 -8672
rect 200808 -8723 200843 -8689
rect 200853 -8723 200854 -8681
rect 200995 -8753 200996 -8525
rect 201685 -8534 201720 -8500
rect 201862 -8534 201897 -8500
rect 202056 -8577 202091 -8543
rect 202101 -8577 202102 -8532
rect 202201 -8543 202202 -8532
rect 202410 -8537 202445 -8503
rect 202455 -8537 202456 -8492
rect 202555 -8503 202556 -8492
rect 202800 -8496 202835 -8462
rect 202845 -8496 202846 -8451
rect 202945 -8462 202946 -8451
rect 202956 -8496 202991 -8462
rect 203001 -8496 203002 -8451
rect 203101 -8462 203102 -8451
rect 203282 -8456 203317 -8422
rect 203354 -8456 203389 -8422
rect 203426 -8456 203461 -8422
rect 203570 -8456 203605 -8422
rect 203642 -8456 203677 -8422
rect 203679 -8456 203749 -8422
rect 203786 -8456 203821 -8422
rect 203856 -8456 203891 -8422
rect 203112 -8496 203147 -8462
rect 204152 -8491 204187 -8457
rect 204197 -8491 204198 -8446
rect 204297 -8457 204298 -8446
rect 204308 -8491 204343 -8457
rect 204353 -8491 204354 -8446
rect 204453 -8457 204454 -8446
rect 205029 -8451 205064 -8417
rect 205206 -8451 205241 -8417
rect 204464 -8491 204499 -8457
rect 202566 -8537 202601 -8503
rect 203845 -8505 203846 -8494
rect 202212 -8577 202247 -8543
rect 201125 -8621 201160 -8587
rect 201326 -8666 201361 -8632
rect 201449 -8637 201450 -8595
rect 201771 -8624 201806 -8590
rect 202410 -8620 202445 -8586
rect 202455 -8620 202456 -8575
rect 202555 -8586 202556 -8575
rect 202800 -8580 202835 -8546
rect 202845 -8580 202846 -8535
rect 202945 -8546 202946 -8535
rect 202956 -8580 202991 -8546
rect 203001 -8580 203002 -8535
rect 203101 -8546 203102 -8535
rect 203679 -8539 203714 -8505
rect 203856 -8539 203891 -8505
rect 203112 -8580 203147 -8546
rect 203999 -8565 204114 -8499
rect 204297 -8525 204298 -8499
rect 204694 -8517 204729 -8483
rect 204739 -8517 204740 -8472
rect 204839 -8483 204840 -8472
rect 204850 -8517 204885 -8483
rect 204895 -8517 204896 -8472
rect 205195 -8500 205196 -8489
rect 205400 -8494 205435 -8460
rect 205445 -8494 205446 -8449
rect 205545 -8460 205546 -8449
rect 205754 -8453 205789 -8419
rect 205799 -8453 205800 -8408
rect 205899 -8419 205900 -8408
rect 206080 -8413 206115 -8379
rect 206144 -8413 206187 -8379
rect 206189 -8413 206190 -8371
rect 206289 -8379 206290 -8371
rect 206224 -8413 206259 -8379
rect 206300 -8413 206335 -8379
rect 206345 -8413 206346 -8371
rect 206445 -8379 206446 -8371
rect 206394 -8413 206429 -8379
rect 206456 -8413 206501 -8379
rect 207496 -8408 207531 -8374
rect 207541 -8408 207542 -8363
rect 207641 -8374 207642 -8363
rect 207652 -8408 207687 -8374
rect 207697 -8408 207698 -8363
rect 207797 -8374 207798 -8363
rect 208373 -8367 208408 -8333
rect 208550 -8367 208585 -8333
rect 209143 -8336 209144 -8328
rect 209243 -8336 209244 -8328
rect 207808 -8408 207843 -8374
rect 205910 -8453 205945 -8419
rect 207189 -8422 207190 -8414
rect 208539 -8417 208540 -8406
rect 208744 -8410 208779 -8376
rect 208789 -8410 208790 -8365
rect 208889 -8376 208890 -8365
rect 209070 -8370 209133 -8336
rect 209142 -8370 209177 -8336
rect 209254 -8370 209289 -8336
rect 209979 -8360 210014 -8326
rect 210075 -8360 210110 -8326
rect 210171 -8360 210206 -8326
rect 210267 -8360 210302 -8326
rect 210363 -8360 210398 -8326
rect 210459 -8360 210494 -8326
rect 210555 -8360 210590 -8326
rect 211883 -8333 211884 -8322
rect 212060 -8327 212123 -8293
rect 212132 -8327 212167 -8293
rect 212244 -8327 212279 -8293
rect 212775 -8317 212810 -8283
rect 212871 -8317 212906 -8283
rect 212967 -8317 213002 -8283
rect 213063 -8317 213098 -8283
rect 213159 -8317 213194 -8283
rect 208900 -8410 208935 -8376
rect 205556 -8494 205591 -8460
rect 202566 -8620 202601 -8586
rect 203845 -8589 203846 -8578
rect 201095 -8689 201096 -8681
rect 201106 -8723 201141 -8689
rect 201326 -8734 201361 -8700
rect 199773 -8793 199808 -8759
rect 199976 -8838 200011 -8804
rect 200099 -8809 200100 -8767
rect 200421 -8796 200456 -8762
rect 199743 -8861 199744 -8853
rect 199754 -8895 199789 -8861
rect 199976 -8906 200011 -8872
rect 199743 -8961 199744 -8950
rect 199754 -8995 199789 -8961
rect 198691 -9045 198726 -9011
rect 198787 -9045 198822 -9011
rect 198883 -9045 198918 -9011
rect 199392 -9035 199427 -9001
rect 199464 -9035 199499 -9001
rect 199536 -9035 199571 -9001
rect 199608 -9029 199644 -9001
rect 199954 -9025 199989 -8991
rect 199999 -9025 200000 -8980
rect 199608 -9035 199643 -9029
rect 199045 -9088 199080 -9054
rect 199141 -9088 199176 -9054
rect 199237 -9088 199272 -9054
rect 200141 -9076 200142 -8809
rect 200770 -8819 201157 -8753
rect 200157 -8860 200192 -8826
rect 200506 -8832 200517 -8819
rect 200440 -8874 200517 -8832
rect 200568 -8874 201157 -8819
rect 201304 -8853 201339 -8819
rect 201349 -8853 201350 -8808
rect 200440 -8877 201157 -8874
rect 200157 -8928 200192 -8894
rect 200360 -8942 200395 -8908
rect 200405 -8942 200406 -8900
rect 200241 -8991 200242 -8980
rect 200252 -9025 200287 -8991
rect 200360 -9042 200395 -9008
rect 200405 -9042 200406 -8997
rect 200253 -9078 200288 -9044
rect 200325 -9078 200360 -9044
rect 200397 -9078 200432 -9044
rect 199399 -9131 199434 -9097
rect 199495 -9131 199530 -9097
rect 199591 -9131 199626 -9097
rect 199687 -9131 199722 -9097
rect 199783 -9131 199818 -9097
rect 200440 -9114 200585 -8877
rect 200770 -8899 201157 -8877
rect 200694 -8925 201157 -8899
rect 201491 -8904 201492 -8637
rect 201507 -8688 201542 -8654
rect 202121 -8691 202156 -8657
rect 202800 -8663 202835 -8629
rect 202845 -8663 202846 -8618
rect 202945 -8629 202946 -8618
rect 202956 -8663 202991 -8629
rect 203001 -8663 203002 -8618
rect 203101 -8629 203102 -8618
rect 203679 -8623 203714 -8589
rect 203856 -8623 203891 -8589
rect 204217 -8605 204252 -8571
rect 203112 -8663 203147 -8629
rect 202945 -8697 202946 -8671
rect 203344 -8689 203379 -8655
rect 203389 -8689 203390 -8644
rect 203489 -8655 203490 -8644
rect 203500 -8689 203535 -8655
rect 203545 -8689 203546 -8644
rect 203845 -8672 203846 -8661
rect 201507 -8756 201542 -8722
rect 201710 -8770 201745 -8736
rect 201755 -8770 201756 -8728
rect 201855 -8740 201856 -8729
rect 202475 -8734 202510 -8700
rect 201866 -8774 201901 -8740
rect 201591 -8819 201592 -8808
rect 202060 -8813 202095 -8779
rect 202105 -8813 202106 -8771
rect 202205 -8779 202206 -8771
rect 202865 -8777 202900 -8743
rect 202216 -8813 202251 -8779
rect 201602 -8853 201637 -8819
rect 201710 -8870 201745 -8836
rect 201755 -8870 201756 -8825
rect 201855 -8832 201856 -8821
rect 201866 -8866 201901 -8832
rect 202414 -8856 202449 -8822
rect 202459 -8856 202460 -8814
rect 202559 -8822 202560 -8814
rect 202570 -8856 202605 -8822
rect 201603 -8906 201638 -8872
rect 201675 -8906 201710 -8872
rect 201747 -8906 201782 -8872
rect 202060 -8913 202095 -8879
rect 202105 -8913 202106 -8868
rect 202205 -8879 202206 -8868
rect 202216 -8913 202251 -8879
rect 202800 -8895 202835 -8861
rect 202845 -8895 202846 -8853
rect 200694 -8959 201170 -8925
rect 202028 -8949 202063 -8915
rect 202100 -8949 202135 -8915
rect 202414 -8956 202449 -8922
rect 202459 -8956 202460 -8911
rect 202559 -8922 202560 -8911
rect 202570 -8956 202605 -8922
rect 200694 -8985 201157 -8959
rect 200698 -8993 200899 -8985
rect 200714 -9003 200883 -8993
rect 200440 -9140 200615 -9114
rect 199947 -9174 199982 -9140
rect 200043 -9174 200078 -9140
rect 200139 -9174 200174 -9140
rect 200235 -9174 200270 -9140
rect 200331 -9174 200366 -9140
rect 200427 -9174 200615 -9140
rect 200440 -9200 200615 -9174
rect 200640 -9174 200741 -9050
rect 200518 -9870 200553 -9200
rect 200640 -9228 200643 -9174
rect 200325 -9936 200470 -9924
rect 199993 -9970 200470 -9936
rect 200325 -9971 200470 -9970
rect 200506 -9971 200553 -9870
rect 200652 -9971 200687 -9174
rect 200910 -9971 200945 -9062
rect 201044 -9971 201079 -8985
rect 201297 -9002 201332 -8968
rect 201393 -9002 201428 -8968
rect 201489 -9002 201524 -8968
rect 201585 -9002 201620 -8968
rect 201681 -9002 201716 -8968
rect 201777 -9002 201812 -8968
rect 201873 -9002 201908 -8968
rect 202382 -8992 202417 -8958
rect 202454 -8992 202489 -8958
rect 202800 -8995 202835 -8961
rect 202845 -8995 202846 -8950
rect 202987 -9001 202988 -8697
rect 203679 -8706 203714 -8672
rect 203856 -8706 203891 -8672
rect 204152 -8723 204187 -8689
rect 204197 -8723 204198 -8681
rect 204339 -8753 204340 -8525
rect 205029 -8534 205064 -8500
rect 205206 -8534 205241 -8500
rect 205400 -8577 205435 -8543
rect 205445 -8577 205446 -8532
rect 205545 -8543 205546 -8532
rect 205754 -8537 205789 -8503
rect 205799 -8537 205800 -8492
rect 205899 -8503 205900 -8492
rect 206144 -8496 206179 -8462
rect 206189 -8496 206190 -8451
rect 206289 -8462 206290 -8451
rect 206300 -8496 206335 -8462
rect 206345 -8496 206346 -8451
rect 206445 -8462 206446 -8451
rect 206626 -8456 206661 -8422
rect 206698 -8456 206733 -8422
rect 206770 -8456 206805 -8422
rect 206914 -8456 206949 -8422
rect 206986 -8456 207021 -8422
rect 207023 -8456 207093 -8422
rect 207130 -8456 207165 -8422
rect 207200 -8456 207235 -8422
rect 206456 -8496 206491 -8462
rect 207496 -8491 207531 -8457
rect 207541 -8491 207542 -8446
rect 207641 -8457 207642 -8446
rect 207652 -8491 207687 -8457
rect 207697 -8491 207698 -8446
rect 207797 -8457 207798 -8446
rect 208373 -8451 208408 -8417
rect 208550 -8451 208585 -8417
rect 207808 -8491 207843 -8457
rect 205910 -8537 205945 -8503
rect 207189 -8505 207190 -8494
rect 205556 -8577 205591 -8543
rect 204469 -8621 204504 -8587
rect 204670 -8666 204705 -8632
rect 204793 -8637 204794 -8595
rect 205115 -8624 205150 -8590
rect 205754 -8620 205789 -8586
rect 205799 -8620 205800 -8575
rect 205899 -8586 205900 -8575
rect 206144 -8580 206179 -8546
rect 206189 -8580 206190 -8535
rect 206289 -8546 206290 -8535
rect 206300 -8580 206335 -8546
rect 206345 -8580 206346 -8535
rect 206445 -8546 206446 -8535
rect 207023 -8539 207058 -8505
rect 207200 -8539 207235 -8505
rect 206456 -8580 206491 -8546
rect 207343 -8565 207458 -8499
rect 207641 -8525 207642 -8499
rect 208038 -8517 208073 -8483
rect 208083 -8517 208084 -8472
rect 208183 -8483 208184 -8472
rect 208194 -8517 208229 -8483
rect 208239 -8517 208240 -8472
rect 208539 -8500 208540 -8489
rect 208744 -8494 208779 -8460
rect 208789 -8494 208790 -8449
rect 208889 -8460 208890 -8449
rect 209098 -8453 209133 -8419
rect 209143 -8453 209144 -8408
rect 209243 -8419 209244 -8408
rect 209424 -8413 209459 -8379
rect 209488 -8413 209531 -8379
rect 209533 -8413 209534 -8371
rect 209633 -8379 209634 -8371
rect 209568 -8413 209603 -8379
rect 209644 -8413 209679 -8379
rect 209689 -8413 209690 -8371
rect 209789 -8379 209790 -8371
rect 209738 -8413 209773 -8379
rect 209800 -8413 209845 -8379
rect 210840 -8408 210875 -8374
rect 210885 -8408 210886 -8363
rect 210985 -8374 210986 -8363
rect 210996 -8408 211031 -8374
rect 211041 -8408 211042 -8363
rect 211141 -8374 211142 -8363
rect 211717 -8367 211752 -8333
rect 211894 -8367 211929 -8333
rect 212487 -8336 212488 -8328
rect 212587 -8336 212588 -8328
rect 211152 -8408 211187 -8374
rect 209254 -8453 209289 -8419
rect 210533 -8422 210534 -8414
rect 211883 -8417 211884 -8406
rect 212088 -8410 212123 -8376
rect 212133 -8410 212134 -8365
rect 212233 -8376 212234 -8365
rect 212414 -8370 212477 -8336
rect 212486 -8370 212521 -8336
rect 212598 -8370 212633 -8336
rect 213323 -8360 213358 -8326
rect 213419 -8360 213454 -8326
rect 213515 -8360 213550 -8326
rect 213611 -8360 213646 -8326
rect 213707 -8360 213742 -8326
rect 213803 -8360 213838 -8326
rect 213899 -8360 213934 -8326
rect 212244 -8410 212279 -8376
rect 208900 -8494 208935 -8460
rect 205910 -8620 205945 -8586
rect 207189 -8589 207190 -8578
rect 204439 -8689 204440 -8681
rect 204450 -8723 204485 -8689
rect 204670 -8734 204705 -8700
rect 203117 -8793 203152 -8759
rect 203320 -8838 203355 -8804
rect 203443 -8809 203444 -8767
rect 203765 -8796 203800 -8762
rect 203087 -8861 203088 -8853
rect 203098 -8895 203133 -8861
rect 203320 -8906 203355 -8872
rect 203087 -8961 203088 -8950
rect 203098 -8995 203133 -8961
rect 202035 -9045 202070 -9011
rect 202131 -9045 202166 -9011
rect 202227 -9045 202262 -9011
rect 202736 -9035 202771 -9001
rect 202808 -9035 202843 -9001
rect 202880 -9035 202915 -9001
rect 202952 -9029 202988 -9001
rect 203298 -9025 203333 -8991
rect 203343 -9025 203344 -8980
rect 202952 -9035 202987 -9029
rect 202389 -9088 202424 -9054
rect 202485 -9088 202520 -9054
rect 202581 -9088 202616 -9054
rect 203485 -9076 203486 -8809
rect 204114 -8819 204501 -8753
rect 203501 -8860 203536 -8826
rect 203850 -8832 203861 -8819
rect 203784 -8874 203861 -8832
rect 203912 -8874 204501 -8819
rect 204648 -8853 204683 -8819
rect 204693 -8853 204694 -8808
rect 203784 -8877 204501 -8874
rect 203501 -8928 203536 -8894
rect 203704 -8942 203739 -8908
rect 203749 -8942 203750 -8900
rect 203585 -8991 203586 -8980
rect 203596 -9025 203631 -8991
rect 203704 -9042 203739 -9008
rect 203749 -9042 203750 -8997
rect 203597 -9078 203632 -9044
rect 203669 -9078 203704 -9044
rect 203741 -9078 203776 -9044
rect 202743 -9131 202778 -9097
rect 202839 -9131 202874 -9097
rect 202935 -9131 202970 -9097
rect 203031 -9131 203066 -9097
rect 203127 -9131 203162 -9097
rect 203784 -9114 203929 -8877
rect 204114 -8899 204501 -8877
rect 204038 -8925 204501 -8899
rect 204835 -8904 204836 -8637
rect 204851 -8688 204886 -8654
rect 205465 -8691 205500 -8657
rect 206144 -8663 206179 -8629
rect 206189 -8663 206190 -8618
rect 206289 -8629 206290 -8618
rect 206300 -8663 206335 -8629
rect 206345 -8663 206346 -8618
rect 206445 -8629 206446 -8618
rect 207023 -8623 207058 -8589
rect 207200 -8623 207235 -8589
rect 207561 -8605 207596 -8571
rect 206456 -8663 206491 -8629
rect 206289 -8697 206290 -8671
rect 206688 -8689 206723 -8655
rect 206733 -8689 206734 -8644
rect 206833 -8655 206834 -8644
rect 206844 -8689 206879 -8655
rect 206889 -8689 206890 -8644
rect 207189 -8672 207190 -8661
rect 204851 -8756 204886 -8722
rect 205054 -8770 205089 -8736
rect 205099 -8770 205100 -8728
rect 205199 -8740 205200 -8729
rect 205819 -8734 205854 -8700
rect 205210 -8774 205245 -8740
rect 204935 -8819 204936 -8808
rect 205404 -8813 205439 -8779
rect 205449 -8813 205450 -8771
rect 205549 -8779 205550 -8771
rect 206209 -8777 206244 -8743
rect 205560 -8813 205595 -8779
rect 204946 -8853 204981 -8819
rect 205054 -8870 205089 -8836
rect 205099 -8870 205100 -8825
rect 205199 -8832 205200 -8821
rect 205210 -8866 205245 -8832
rect 205758 -8856 205793 -8822
rect 205803 -8856 205804 -8814
rect 205903 -8822 205904 -8814
rect 205914 -8856 205949 -8822
rect 204947 -8906 204982 -8872
rect 205019 -8906 205054 -8872
rect 205091 -8906 205126 -8872
rect 205404 -8913 205439 -8879
rect 205449 -8913 205450 -8868
rect 205549 -8879 205550 -8868
rect 205560 -8913 205595 -8879
rect 206144 -8895 206179 -8861
rect 206189 -8895 206190 -8853
rect 204038 -8959 204514 -8925
rect 205372 -8949 205407 -8915
rect 205444 -8949 205479 -8915
rect 205758 -8956 205793 -8922
rect 205803 -8956 205804 -8911
rect 205903 -8922 205904 -8911
rect 205914 -8956 205949 -8922
rect 204038 -8985 204501 -8959
rect 204042 -8993 204243 -8985
rect 204058 -9003 204227 -8993
rect 203784 -9140 203959 -9114
rect 203291 -9174 203326 -9140
rect 203387 -9174 203422 -9140
rect 203483 -9174 203518 -9140
rect 203579 -9174 203614 -9140
rect 203675 -9174 203710 -9140
rect 203771 -9174 203959 -9140
rect 203784 -9200 203959 -9174
rect 203984 -9174 204085 -9050
rect 203862 -9870 203897 -9200
rect 203984 -9228 203987 -9174
rect 203669 -9936 203814 -9924
rect 203337 -9970 203814 -9936
rect 203669 -9971 203814 -9970
rect 203850 -9971 203897 -9870
rect 203996 -9971 204031 -9174
rect 204254 -9971 204289 -9062
rect 204388 -9971 204423 -8985
rect 204641 -9002 204676 -8968
rect 204737 -9002 204772 -8968
rect 204833 -9002 204868 -8968
rect 204929 -9002 204964 -8968
rect 205025 -9002 205060 -8968
rect 205121 -9002 205156 -8968
rect 205217 -9002 205252 -8968
rect 205726 -8992 205761 -8958
rect 205798 -8992 205833 -8958
rect 206144 -8995 206179 -8961
rect 206189 -8995 206190 -8950
rect 206331 -9001 206332 -8697
rect 207023 -8706 207058 -8672
rect 207200 -8706 207235 -8672
rect 207496 -8723 207531 -8689
rect 207541 -8723 207542 -8681
rect 207683 -8753 207684 -8525
rect 208373 -8534 208408 -8500
rect 208550 -8534 208585 -8500
rect 208744 -8577 208779 -8543
rect 208789 -8577 208790 -8532
rect 208889 -8543 208890 -8532
rect 209098 -8537 209133 -8503
rect 209143 -8537 209144 -8492
rect 209243 -8503 209244 -8492
rect 209488 -8496 209523 -8462
rect 209533 -8496 209534 -8451
rect 209633 -8462 209634 -8451
rect 209644 -8496 209679 -8462
rect 209689 -8496 209690 -8451
rect 209789 -8462 209790 -8451
rect 209970 -8456 210005 -8422
rect 210042 -8456 210077 -8422
rect 210114 -8456 210149 -8422
rect 210258 -8456 210293 -8422
rect 210330 -8456 210365 -8422
rect 210367 -8456 210437 -8422
rect 210474 -8456 210509 -8422
rect 210544 -8456 210579 -8422
rect 209800 -8496 209835 -8462
rect 210840 -8491 210875 -8457
rect 210885 -8491 210886 -8446
rect 210985 -8457 210986 -8446
rect 210996 -8491 211031 -8457
rect 211041 -8491 211042 -8446
rect 211141 -8457 211142 -8446
rect 211717 -8451 211752 -8417
rect 211894 -8451 211929 -8417
rect 211152 -8491 211187 -8457
rect 209254 -8537 209289 -8503
rect 210533 -8505 210534 -8494
rect 208900 -8577 208935 -8543
rect 207813 -8621 207848 -8587
rect 208014 -8666 208049 -8632
rect 208137 -8637 208138 -8595
rect 208459 -8624 208494 -8590
rect 209098 -8620 209133 -8586
rect 209143 -8620 209144 -8575
rect 209243 -8586 209244 -8575
rect 209488 -8580 209523 -8546
rect 209533 -8580 209534 -8535
rect 209633 -8546 209634 -8535
rect 209644 -8580 209679 -8546
rect 209689 -8580 209690 -8535
rect 209789 -8546 209790 -8535
rect 210367 -8539 210402 -8505
rect 210544 -8539 210579 -8505
rect 209800 -8580 209835 -8546
rect 210687 -8565 210802 -8499
rect 210985 -8525 210986 -8499
rect 211382 -8517 211417 -8483
rect 211427 -8517 211428 -8472
rect 211527 -8483 211528 -8472
rect 211538 -8517 211573 -8483
rect 211583 -8517 211584 -8472
rect 211883 -8500 211884 -8489
rect 212088 -8494 212123 -8460
rect 212133 -8494 212134 -8449
rect 212233 -8460 212234 -8449
rect 212442 -8453 212477 -8419
rect 212487 -8453 212488 -8408
rect 212587 -8419 212588 -8408
rect 212768 -8413 212803 -8379
rect 212832 -8413 212875 -8379
rect 212877 -8413 212878 -8371
rect 212977 -8379 212978 -8371
rect 212912 -8413 212947 -8379
rect 212988 -8413 213023 -8379
rect 213033 -8413 213034 -8371
rect 213133 -8379 213134 -8371
rect 213082 -8413 213117 -8379
rect 213144 -8413 213189 -8379
rect 212598 -8453 212633 -8419
rect 213877 -8422 213878 -8414
rect 212244 -8494 212279 -8460
rect 209254 -8620 209289 -8586
rect 210533 -8589 210534 -8578
rect 207783 -8689 207784 -8681
rect 207794 -8723 207829 -8689
rect 208014 -8734 208049 -8700
rect 206461 -8793 206496 -8759
rect 206664 -8838 206699 -8804
rect 206787 -8809 206788 -8767
rect 207109 -8796 207144 -8762
rect 206431 -8861 206432 -8853
rect 206442 -8895 206477 -8861
rect 206664 -8906 206699 -8872
rect 206431 -8961 206432 -8950
rect 206442 -8995 206477 -8961
rect 205379 -9045 205414 -9011
rect 205475 -9045 205510 -9011
rect 205571 -9045 205606 -9011
rect 206080 -9035 206115 -9001
rect 206152 -9035 206187 -9001
rect 206224 -9035 206259 -9001
rect 206296 -9029 206332 -9001
rect 206642 -9025 206677 -8991
rect 206687 -9025 206688 -8980
rect 206296 -9035 206331 -9029
rect 205733 -9088 205768 -9054
rect 205829 -9088 205864 -9054
rect 205925 -9088 205960 -9054
rect 206829 -9076 206830 -8809
rect 207458 -8819 207845 -8753
rect 206845 -8860 206880 -8826
rect 207194 -8832 207205 -8819
rect 207128 -8874 207205 -8832
rect 207256 -8874 207845 -8819
rect 207992 -8853 208027 -8819
rect 208037 -8853 208038 -8808
rect 207128 -8877 207845 -8874
rect 206845 -8928 206880 -8894
rect 207048 -8942 207083 -8908
rect 207093 -8942 207094 -8900
rect 206929 -8991 206930 -8980
rect 206940 -9025 206975 -8991
rect 207048 -9042 207083 -9008
rect 207093 -9042 207094 -8997
rect 206941 -9078 206976 -9044
rect 207013 -9078 207048 -9044
rect 207085 -9078 207120 -9044
rect 206087 -9131 206122 -9097
rect 206183 -9131 206218 -9097
rect 206279 -9131 206314 -9097
rect 206375 -9131 206410 -9097
rect 206471 -9131 206506 -9097
rect 207128 -9114 207273 -8877
rect 207458 -8899 207845 -8877
rect 207382 -8925 207845 -8899
rect 208179 -8904 208180 -8637
rect 208195 -8688 208230 -8654
rect 208809 -8691 208844 -8657
rect 209488 -8663 209523 -8629
rect 209533 -8663 209534 -8618
rect 209633 -8629 209634 -8618
rect 209644 -8663 209679 -8629
rect 209689 -8663 209690 -8618
rect 209789 -8629 209790 -8618
rect 210367 -8623 210402 -8589
rect 210544 -8623 210579 -8589
rect 210905 -8605 210940 -8571
rect 209800 -8663 209835 -8629
rect 209633 -8697 209634 -8671
rect 210032 -8689 210067 -8655
rect 210077 -8689 210078 -8644
rect 210177 -8655 210178 -8644
rect 210188 -8689 210223 -8655
rect 210233 -8689 210234 -8644
rect 210533 -8672 210534 -8661
rect 208195 -8756 208230 -8722
rect 208398 -8770 208433 -8736
rect 208443 -8770 208444 -8728
rect 208543 -8740 208544 -8729
rect 209163 -8734 209198 -8700
rect 208554 -8774 208589 -8740
rect 208279 -8819 208280 -8808
rect 208748 -8813 208783 -8779
rect 208793 -8813 208794 -8771
rect 208893 -8779 208894 -8771
rect 209553 -8777 209588 -8743
rect 208904 -8813 208939 -8779
rect 208290 -8853 208325 -8819
rect 208398 -8870 208433 -8836
rect 208443 -8870 208444 -8825
rect 208543 -8832 208544 -8821
rect 208554 -8866 208589 -8832
rect 209102 -8856 209137 -8822
rect 209147 -8856 209148 -8814
rect 209247 -8822 209248 -8814
rect 209258 -8856 209293 -8822
rect 208291 -8906 208326 -8872
rect 208363 -8906 208398 -8872
rect 208435 -8906 208470 -8872
rect 208748 -8913 208783 -8879
rect 208793 -8913 208794 -8868
rect 208893 -8879 208894 -8868
rect 208904 -8913 208939 -8879
rect 209488 -8895 209523 -8861
rect 209533 -8895 209534 -8853
rect 207382 -8959 207858 -8925
rect 208716 -8949 208751 -8915
rect 208788 -8949 208823 -8915
rect 209102 -8956 209137 -8922
rect 209147 -8956 209148 -8911
rect 209247 -8922 209248 -8911
rect 209258 -8956 209293 -8922
rect 207382 -8985 207845 -8959
rect 207386 -8993 207587 -8985
rect 207402 -9003 207571 -8993
rect 207128 -9140 207303 -9114
rect 206635 -9174 206670 -9140
rect 206731 -9174 206766 -9140
rect 206827 -9174 206862 -9140
rect 206923 -9174 206958 -9140
rect 207019 -9174 207054 -9140
rect 207115 -9174 207303 -9140
rect 207128 -9200 207303 -9174
rect 207328 -9174 207429 -9050
rect 207206 -9870 207241 -9200
rect 207328 -9228 207331 -9174
rect 207013 -9936 207158 -9924
rect 206681 -9970 207158 -9936
rect 207013 -9971 207158 -9970
rect 207194 -9971 207241 -9870
rect 207340 -9971 207375 -9174
rect 207598 -9971 207633 -9062
rect 207732 -9971 207767 -8985
rect 207985 -9002 208020 -8968
rect 208081 -9002 208116 -8968
rect 208177 -9002 208212 -8968
rect 208273 -9002 208308 -8968
rect 208369 -9002 208404 -8968
rect 208465 -9002 208500 -8968
rect 208561 -9002 208596 -8968
rect 209070 -8992 209105 -8958
rect 209142 -8992 209177 -8958
rect 209488 -8995 209523 -8961
rect 209533 -8995 209534 -8950
rect 209675 -9001 209676 -8697
rect 210367 -8706 210402 -8672
rect 210544 -8706 210579 -8672
rect 210840 -8723 210875 -8689
rect 210885 -8723 210886 -8681
rect 211027 -8753 211028 -8525
rect 211717 -8534 211752 -8500
rect 211894 -8534 211929 -8500
rect 212088 -8577 212123 -8543
rect 212133 -8577 212134 -8532
rect 212233 -8543 212234 -8532
rect 212442 -8537 212477 -8503
rect 212487 -8537 212488 -8492
rect 212587 -8503 212588 -8492
rect 212832 -8496 212867 -8462
rect 212877 -8496 212878 -8451
rect 212977 -8462 212978 -8451
rect 212988 -8496 213023 -8462
rect 213033 -8496 213034 -8451
rect 213133 -8462 213134 -8451
rect 213314 -8456 213349 -8422
rect 213386 -8456 213421 -8422
rect 213458 -8456 213493 -8422
rect 213602 -8456 213637 -8422
rect 213674 -8456 213709 -8422
rect 213711 -8456 213781 -8422
rect 213818 -8456 213853 -8422
rect 213888 -8456 213923 -8422
rect 213144 -8496 213179 -8462
rect 212598 -8537 212633 -8503
rect 213877 -8505 213878 -8494
rect 212244 -8577 212279 -8543
rect 211157 -8621 211192 -8587
rect 211358 -8666 211393 -8632
rect 211481 -8637 211482 -8595
rect 211803 -8624 211838 -8590
rect 212442 -8620 212477 -8586
rect 212487 -8620 212488 -8575
rect 212587 -8586 212588 -8575
rect 212832 -8580 212867 -8546
rect 212877 -8580 212878 -8535
rect 212977 -8546 212978 -8535
rect 212988 -8580 213023 -8546
rect 213033 -8580 213034 -8535
rect 213133 -8546 213134 -8535
rect 213711 -8539 213746 -8505
rect 213888 -8539 213923 -8505
rect 213144 -8580 213179 -8546
rect 214031 -8565 214147 -8499
rect 212598 -8620 212633 -8586
rect 213877 -8589 213878 -8578
rect 211127 -8689 211128 -8681
rect 211138 -8723 211173 -8689
rect 211358 -8734 211393 -8700
rect 209805 -8793 209840 -8759
rect 210008 -8838 210043 -8804
rect 210131 -8809 210132 -8767
rect 210453 -8796 210488 -8762
rect 209775 -8861 209776 -8853
rect 209786 -8895 209821 -8861
rect 210008 -8906 210043 -8872
rect 209775 -8961 209776 -8950
rect 209786 -8995 209821 -8961
rect 208723 -9045 208758 -9011
rect 208819 -9045 208854 -9011
rect 208915 -9045 208950 -9011
rect 209424 -9035 209459 -9001
rect 209496 -9035 209531 -9001
rect 209568 -9035 209603 -9001
rect 209640 -9029 209676 -9001
rect 209986 -9025 210021 -8991
rect 210031 -9025 210032 -8980
rect 209640 -9035 209675 -9029
rect 209077 -9088 209112 -9054
rect 209173 -9088 209208 -9054
rect 209269 -9088 209304 -9054
rect 210173 -9076 210174 -8809
rect 210802 -8819 211189 -8753
rect 210189 -8860 210224 -8826
rect 210538 -8832 210549 -8819
rect 210472 -8874 210549 -8832
rect 210600 -8874 211189 -8819
rect 211336 -8853 211371 -8819
rect 211381 -8853 211382 -8808
rect 210472 -8877 211189 -8874
rect 210189 -8928 210224 -8894
rect 210392 -8942 210427 -8908
rect 210437 -8942 210438 -8900
rect 210273 -8991 210274 -8980
rect 210284 -9025 210319 -8991
rect 210392 -9042 210427 -9008
rect 210437 -9042 210438 -8997
rect 210285 -9078 210320 -9044
rect 210357 -9078 210392 -9044
rect 210429 -9078 210464 -9044
rect 209431 -9131 209466 -9097
rect 209527 -9131 209562 -9097
rect 209623 -9131 209658 -9097
rect 209719 -9131 209754 -9097
rect 209815 -9131 209850 -9097
rect 210472 -9114 210617 -8877
rect 210802 -8899 211189 -8877
rect 210726 -8925 211189 -8899
rect 211523 -8904 211524 -8637
rect 211539 -8688 211574 -8654
rect 212153 -8691 212188 -8657
rect 212832 -8663 212867 -8629
rect 212877 -8663 212878 -8618
rect 212977 -8629 212978 -8618
rect 212988 -8663 213023 -8629
rect 213033 -8663 213034 -8618
rect 213133 -8629 213134 -8618
rect 213711 -8623 213746 -8589
rect 213888 -8623 213923 -8589
rect 213144 -8663 213179 -8629
rect 212977 -8697 212978 -8671
rect 213376 -8689 213411 -8655
rect 213421 -8689 213422 -8644
rect 213521 -8655 213522 -8644
rect 213532 -8689 213567 -8655
rect 213577 -8689 213578 -8644
rect 213877 -8672 213878 -8661
rect 211539 -8756 211574 -8722
rect 211742 -8770 211777 -8736
rect 211787 -8770 211788 -8728
rect 211887 -8740 211888 -8729
rect 212507 -8734 212542 -8700
rect 211898 -8774 211933 -8740
rect 211623 -8819 211624 -8808
rect 212092 -8813 212127 -8779
rect 212137 -8813 212138 -8771
rect 212237 -8779 212238 -8771
rect 212897 -8777 212932 -8743
rect 212248 -8813 212283 -8779
rect 211634 -8853 211669 -8819
rect 211742 -8870 211777 -8836
rect 211787 -8870 211788 -8825
rect 211887 -8832 211888 -8821
rect 211898 -8866 211933 -8832
rect 212446 -8856 212481 -8822
rect 212491 -8856 212492 -8814
rect 212591 -8822 212592 -8814
rect 212602 -8856 212637 -8822
rect 211635 -8906 211670 -8872
rect 211707 -8906 211742 -8872
rect 211779 -8906 211814 -8872
rect 212092 -8913 212127 -8879
rect 212137 -8913 212138 -8868
rect 212237 -8879 212238 -8868
rect 212248 -8913 212283 -8879
rect 212832 -8895 212867 -8861
rect 212877 -8895 212878 -8853
rect 210726 -8959 211202 -8925
rect 212060 -8949 212095 -8915
rect 212132 -8949 212167 -8915
rect 212446 -8956 212481 -8922
rect 212491 -8956 212492 -8911
rect 212591 -8922 212592 -8911
rect 212602 -8956 212637 -8922
rect 210726 -8985 211189 -8959
rect 210730 -8993 210931 -8985
rect 210746 -9003 210915 -8993
rect 210472 -9140 210647 -9114
rect 209979 -9174 210014 -9140
rect 210075 -9174 210110 -9140
rect 210171 -9174 210206 -9140
rect 210267 -9174 210302 -9140
rect 210363 -9174 210398 -9140
rect 210459 -9174 210647 -9140
rect 210472 -9200 210647 -9174
rect 210672 -9174 210773 -9050
rect 210550 -9870 210585 -9200
rect 210672 -9228 210675 -9174
rect 210357 -9936 210502 -9924
rect 210025 -9970 210502 -9936
rect 210357 -9971 210502 -9970
rect 210538 -9971 210585 -9870
rect 210684 -9971 210719 -9174
rect 210942 -9971 210977 -9062
rect 211076 -9971 211111 -8985
rect 211329 -9002 211364 -8968
rect 211425 -9002 211460 -8968
rect 211521 -9002 211556 -8968
rect 211617 -9002 211652 -8968
rect 211713 -9002 211748 -8968
rect 211809 -9002 211844 -8968
rect 211905 -9002 211940 -8968
rect 212414 -8992 212449 -8958
rect 212486 -8992 212521 -8958
rect 212832 -8995 212867 -8961
rect 212877 -8995 212878 -8950
rect 213019 -9001 213020 -8697
rect 213711 -8706 213746 -8672
rect 213888 -8706 213923 -8672
rect 213149 -8793 213184 -8759
rect 213352 -8838 213387 -8804
rect 213475 -8809 213476 -8767
rect 213797 -8796 213832 -8762
rect 213119 -8861 213120 -8853
rect 213130 -8895 213165 -8861
rect 213352 -8906 213387 -8872
rect 213119 -8961 213120 -8950
rect 213130 -8995 213165 -8961
rect 212067 -9045 212102 -9011
rect 212163 -9045 212198 -9011
rect 212259 -9045 212294 -9011
rect 212768 -9035 212803 -9001
rect 212840 -9035 212875 -9001
rect 212912 -9035 212947 -9001
rect 212984 -9029 213020 -9001
rect 213330 -9025 213365 -8991
rect 213375 -9025 213376 -8980
rect 212984 -9035 213019 -9029
rect 212421 -9088 212456 -9054
rect 212517 -9088 212552 -9054
rect 212613 -9088 212648 -9054
rect 213517 -9076 213518 -8809
rect 214147 -8819 214533 -8753
rect 213533 -8860 213568 -8826
rect 213882 -8832 213893 -8819
rect 213816 -8874 213893 -8832
rect 213945 -8874 214533 -8819
rect 213816 -8877 214533 -8874
rect 213533 -8928 213568 -8894
rect 213736 -8942 213771 -8908
rect 213781 -8942 213782 -8900
rect 213617 -8991 213618 -8980
rect 213628 -9025 213663 -8991
rect 213736 -9042 213771 -9008
rect 213781 -9042 213782 -8997
rect 213629 -9078 213664 -9044
rect 213701 -9078 213736 -9044
rect 213773 -9078 213808 -9044
rect 212775 -9131 212810 -9097
rect 212871 -9131 212906 -9097
rect 212967 -9131 213002 -9097
rect 213063 -9131 213098 -9097
rect 213159 -9131 213194 -9097
rect 213816 -9114 213961 -8877
rect 214147 -8899 214533 -8877
rect 214071 -8985 214533 -8899
rect 214074 -8993 214275 -8985
rect 214090 -9003 214259 -8993
rect 213816 -9140 213991 -9114
rect 213323 -9174 213358 -9140
rect 213419 -9174 213454 -9140
rect 213515 -9174 213550 -9140
rect 213611 -9174 213646 -9140
rect 213707 -9174 213742 -9140
rect 213803 -9174 213991 -9140
rect 213816 -9200 213991 -9174
rect 214016 -9174 214117 -9050
rect 213894 -9870 213929 -9200
rect 214016 -9228 214019 -9174
rect 213701 -9936 213846 -9924
rect 213369 -9970 213846 -9936
rect 213701 -9971 213846 -9970
rect 213882 -9971 213929 -9870
rect 214028 -9971 214063 -9174
rect 214286 -9971 214321 -9062
rect 214420 -9971 214455 -8985
rect 3135 -10032 3802 -9971
rect 6479 -10032 7146 -9971
rect 9824 -10032 10490 -9971
rect 13168 -10032 13834 -9971
rect 16513 -10032 17178 -9971
rect 19857 -10032 20522 -9971
rect 23201 -10032 23866 -9971
rect 26545 -10032 27210 -9971
rect 29774 -9982 30554 -9971
rect 33118 -9982 33898 -9971
rect 36462 -9982 37242 -9971
rect 39806 -9982 40586 -9971
rect 43150 -9982 43930 -9971
rect 46494 -9982 47274 -9971
rect 49838 -9982 50618 -9971
rect 53182 -9982 53962 -9971
rect 56527 -9982 57306 -9971
rect 59871 -9982 60650 -9971
rect 63215 -9982 63994 -9971
rect 66559 -9982 67338 -9971
rect 69903 -9982 70682 -9971
rect 73247 -9982 74026 -9971
rect 76591 -9982 77370 -9971
rect 79935 -9982 80714 -9971
rect 83279 -9982 84058 -9971
rect 86623 -9982 87402 -9971
rect 89967 -9982 90746 -9971
rect 93311 -9982 94090 -9971
rect 96655 -9982 97434 -9971
rect 99999 -9982 100778 -9971
rect 103343 -9982 104122 -9971
rect 106687 -9982 107466 -9971
rect 110037 -9982 110810 -9971
rect 113381 -9982 114154 -9971
rect 116725 -9982 117498 -9971
rect 120069 -9982 120842 -9971
rect 123413 -9982 124186 -9971
rect 126757 -9982 127530 -9971
rect 130101 -9982 130874 -9971
rect 133445 -9982 134218 -9971
rect 136789 -9982 137562 -9971
rect 140133 -9982 140906 -9971
rect 143477 -9982 144250 -9971
rect 146821 -9982 147594 -9971
rect 150165 -9982 150938 -9971
rect 153509 -9982 154282 -9971
rect 156853 -9982 157626 -9971
rect 160197 -9982 160970 -9971
rect 163541 -9982 164314 -9971
rect 166885 -9982 167658 -9971
rect 170229 -9982 171002 -9971
rect 173573 -9982 174346 -9971
rect 176917 -9982 177690 -9971
rect 180261 -9982 181034 -9971
rect 183605 -9982 184378 -9971
rect 186949 -9982 187722 -9971
rect 190293 -9982 191066 -9971
rect 193637 -9982 194410 -9971
rect 196981 -9982 197754 -9971
rect 200325 -9982 201098 -9971
rect 203669 -9982 204442 -9971
rect 207013 -9982 207786 -9971
rect 210357 -9982 211130 -9971
rect 213701 -9982 214474 -9971
rect 29860 -10007 30554 -9982
rect 33204 -10007 33898 -9982
rect 36548 -10007 37242 -9982
rect 39892 -10007 40586 -9982
rect 43236 -10007 43930 -9982
rect 46580 -10007 47274 -9982
rect 49924 -10007 50618 -9982
rect 53268 -10007 53962 -9982
rect 56613 -10007 57306 -9982
rect 59957 -10007 60650 -9982
rect 63301 -10007 63994 -9982
rect 66645 -10007 67338 -9982
rect 69989 -10007 70682 -9982
rect 73333 -10007 74026 -9982
rect 76677 -10007 77370 -9982
rect 80021 -10007 80714 -9982
rect 83365 -10007 84058 -9982
rect 86709 -10007 87402 -9982
rect 90053 -10007 90746 -9982
rect 93397 -10007 94090 -9982
rect 96741 -10007 97434 -9982
rect 100085 -10007 100778 -9982
rect 103429 -10007 104122 -9982
rect 106773 -10007 107466 -9982
rect 110123 -10007 110810 -9982
rect 113467 -10007 114154 -9982
rect 116811 -10007 117498 -9982
rect 120155 -10007 120842 -9982
rect 123499 -10007 124186 -9982
rect 126843 -10007 127530 -9982
rect 130187 -10007 130874 -9982
rect 133531 -10007 134218 -9982
rect 136875 -10007 137562 -9982
rect 140219 -10007 140906 -9982
rect 143563 -10007 144250 -9982
rect 146907 -10007 147594 -9982
rect 150251 -10007 150938 -9982
rect 153595 -10007 154282 -9982
rect 156939 -10007 157626 -9982
rect 160283 -10007 160970 -9982
rect 163627 -10007 164314 -9982
rect 166971 -10007 167658 -9982
rect 170315 -10007 171002 -9982
rect 173659 -10007 174346 -9982
rect 177003 -10007 177690 -9982
rect 180347 -10007 181034 -9982
rect 183691 -10007 184378 -9982
rect 187035 -10007 187722 -9982
rect 190379 -10007 191066 -9982
rect 193723 -10007 194410 -9982
rect 197067 -10007 197754 -9982
rect 200411 -10007 201098 -9982
rect 203755 -10007 204442 -9982
rect 207099 -10007 207786 -9982
rect 210443 -10007 211130 -9982
rect 213787 -10007 214474 -9982
rect 29890 -10032 30554 -10007
rect 33234 -10032 33898 -10007
rect 36578 -10032 37242 -10007
rect 39922 -10032 40586 -10007
rect 43266 -10032 43930 -10007
rect 46610 -10032 47274 -10007
rect 49954 -10032 50618 -10007
rect 53298 -10032 53962 -10007
rect 2591 -10194 2636 -10032
rect 3117 -10036 3802 -10032
rect 2787 -10108 2966 -10074
rect 3117 -10128 3861 -10036
rect 3870 -10118 4249 -10084
rect 2725 -10182 2770 -10151
rect 2771 -10182 2781 -10156
rect 2952 -10182 3040 -10155
rect 2713 -10194 3096 -10182
rect 2591 -10228 3096 -10194
rect 2557 -10240 2558 -10228
rect 2591 -10240 2636 -10228
rect 2713 -10229 3096 -10228
rect 3105 -10229 3861 -10128
rect 4331 -10180 4345 -10118
rect 2713 -10240 3861 -10229
rect 2525 -10506 2570 -10240
rect 2579 -10506 2636 -10240
rect 2725 -10301 2770 -10240
rect 2713 -10316 2770 -10301
rect 2771 -10316 2781 -10240
rect 2952 -10265 3861 -10240
rect 3970 -10256 4149 -10222
rect 2713 -10332 2772 -10316
rect 2888 -10332 2935 -10285
rect 2713 -10366 2935 -10332
rect 2646 -10506 2648 -10413
rect 2658 -10506 2670 -10409
rect 2691 -10413 2692 -10409
rect 2713 -10413 2771 -10366
rect 2983 -10385 3028 -10265
rect 2949 -10413 2950 -10409
rect 2691 -10415 2698 -10413
rect 2719 -10415 2770 -10413
rect 2949 -10414 2956 -10413
rect 2691 -10425 2692 -10415
rect 2687 -10506 2692 -10425
rect 2725 -10506 2770 -10415
rect 2905 -10425 2956 -10414
rect 2916 -10506 2956 -10425
rect 2977 -10506 3028 -10385
rect 3038 -10506 3040 -10265
rect 3050 -10342 3861 -10265
rect 4288 -10276 4297 -10220
rect 4300 -10276 4345 -10180
rect 3896 -10330 3905 -10294
rect 3908 -10330 3953 -10306
rect 3954 -10330 3964 -10295
rect 4155 -10306 4165 -10295
rect 4166 -10330 4211 -10306
rect 4214 -10330 4223 -10294
rect 3896 -10342 4223 -10330
rect 4234 -10341 4279 -10330
rect 3050 -10376 4223 -10342
rect 3050 -10388 3887 -10376
rect 3896 -10388 4223 -10376
rect 3050 -10448 3861 -10388
rect 3896 -10448 3905 -10388
rect 3908 -10448 3953 -10388
rect 3954 -10448 3964 -10388
rect 4071 -10448 4109 -10442
rect 4166 -10448 4211 -10388
rect 4212 -10448 4223 -10388
rect 4232 -10448 4279 -10341
rect 4288 -10395 4345 -10276
rect 4286 -10448 4345 -10395
rect 4365 -10245 4379 -10149
rect 4461 -10183 4840 -10149
rect 4365 -10407 4410 -10245
rect 4413 -10395 4422 -10285
rect 4561 -10321 4740 -10287
rect 4879 -10341 4888 -10285
rect 4891 -10341 4936 -10245
rect 4487 -10395 4496 -10359
rect 4499 -10395 4544 -10371
rect 4545 -10395 4555 -10360
rect 4746 -10371 4756 -10360
rect 4757 -10395 4802 -10371
rect 4805 -10395 4814 -10359
rect 4487 -10407 4814 -10395
rect 4365 -10441 4814 -10407
rect 4825 -10441 4870 -10395
rect 4365 -10448 4410 -10441
rect 3050 -10506 4482 -10448
rect 2525 -10543 4482 -10506
rect 4487 -10453 4814 -10441
rect 4487 -10514 4496 -10453
rect 4499 -10514 4544 -10453
rect 4487 -10529 4544 -10514
rect 4545 -10529 4555 -10453
rect 4487 -10543 4545 -10529
rect 4662 -10543 4700 -10507
rect 4757 -10543 4802 -10453
rect 4805 -10543 4814 -10453
rect 4824 -10543 4870 -10441
rect 4879 -10543 4936 -10341
rect 5935 -10506 5980 -10032
rect 6461 -10036 7146 -10032
rect 6131 -10108 6310 -10074
rect 6069 -10506 6114 -10167
rect 6115 -10506 6125 -10156
rect 6316 -10167 6326 -10156
rect 6327 -10506 6372 -10167
rect 6461 -10448 7205 -10036
rect 7214 -10118 7593 -10084
rect 7675 -10180 7689 -10118
rect 7314 -10256 7493 -10222
rect 7240 -10448 7249 -10294
rect 7252 -10448 7297 -10306
rect 7298 -10448 7308 -10295
rect 7499 -10306 7509 -10295
rect 7510 -10448 7555 -10306
rect 7558 -10448 7567 -10294
rect 7632 -10448 7641 -10220
rect 7644 -10448 7689 -10180
rect 7709 -10245 7723 -10149
rect 7805 -10183 8184 -10149
rect 7709 -10448 7754 -10245
rect 7757 -10448 7766 -10285
rect 7905 -10321 8084 -10287
rect 6461 -10506 7826 -10448
rect 5888 -10543 7826 -10506
rect 7831 -10543 7840 -10359
rect 7843 -10543 7888 -10371
rect 7889 -10543 7899 -10360
rect 8090 -10371 8100 -10360
rect 8101 -10543 8146 -10371
rect 8149 -10543 8158 -10359
rect 8223 -10543 8232 -10285
rect 8235 -10543 8280 -10245
rect 9280 -10506 9324 -10032
rect 9806 -10036 10490 -10032
rect 9476 -10108 9654 -10074
rect 9414 -10506 9458 -10167
rect 9460 -10506 9469 -10156
rect 9661 -10167 9670 -10156
rect 9672 -10506 9716 -10167
rect 9806 -10448 10549 -10036
rect 10559 -10118 10937 -10084
rect 11020 -10180 11033 -10118
rect 10659 -10256 10837 -10222
rect 10585 -10448 10593 -10294
rect 10597 -10448 10641 -10306
rect 10643 -10448 10652 -10295
rect 10844 -10306 10853 -10295
rect 10855 -10448 10899 -10306
rect 10903 -10448 10911 -10294
rect 10977 -10448 10985 -10220
rect 10989 -10448 11033 -10180
rect 11054 -10245 11067 -10149
rect 11150 -10183 11528 -10149
rect 11054 -10448 11098 -10245
rect 11102 -10448 11110 -10285
rect 11250 -10321 11428 -10287
rect 9806 -10506 11170 -10448
rect 9233 -10543 11170 -10506
rect 11176 -10543 11184 -10359
rect 11188 -10543 11232 -10371
rect 11234 -10543 11243 -10360
rect 11435 -10371 11444 -10360
rect 11446 -10543 11490 -10371
rect 11494 -10543 11502 -10359
rect 11568 -10543 11576 -10285
rect 11580 -10543 11624 -10245
rect 12624 -10506 12668 -10032
rect 13150 -10036 13834 -10032
rect 12820 -10108 12998 -10074
rect 12758 -10506 12802 -10167
rect 12804 -10506 12813 -10156
rect 13005 -10167 13014 -10156
rect 13016 -10506 13060 -10167
rect 13150 -10448 13893 -10036
rect 13903 -10118 14281 -10084
rect 14364 -10180 14377 -10118
rect 14003 -10256 14181 -10222
rect 13929 -10448 13937 -10294
rect 13941 -10448 13985 -10306
rect 13987 -10448 13996 -10295
rect 14188 -10306 14197 -10295
rect 14199 -10448 14243 -10306
rect 14247 -10448 14255 -10294
rect 14321 -10448 14329 -10220
rect 14333 -10448 14377 -10180
rect 14398 -10245 14411 -10149
rect 14494 -10183 14872 -10149
rect 14398 -10448 14442 -10245
rect 14446 -10448 14454 -10285
rect 14594 -10321 14772 -10287
rect 13150 -10506 14514 -10448
rect 12577 -10543 14514 -10506
rect 14520 -10543 14528 -10359
rect 14532 -10543 14576 -10371
rect 14578 -10543 14587 -10360
rect 14779 -10371 14788 -10360
rect 14790 -10543 14834 -10371
rect 14838 -10543 14846 -10359
rect 14912 -10543 14920 -10285
rect 14924 -10543 14968 -10245
rect 15969 -10506 16012 -10032
rect 16495 -10036 17178 -10032
rect 16165 -10108 16342 -10074
rect 16103 -10506 16146 -10167
rect 16149 -10506 16157 -10156
rect 16350 -10167 16358 -10156
rect 16361 -10506 16404 -10167
rect 16495 -10448 17237 -10036
rect 17248 -10118 17625 -10084
rect 17709 -10180 17721 -10118
rect 17348 -10256 17525 -10222
rect 17274 -10448 17281 -10294
rect 17286 -10448 17329 -10306
rect 17332 -10448 17340 -10295
rect 17533 -10306 17541 -10295
rect 17544 -10448 17587 -10306
rect 17592 -10448 17599 -10294
rect 17666 -10448 17673 -10220
rect 17678 -10448 17721 -10180
rect 17743 -10245 17755 -10149
rect 17839 -10183 18216 -10149
rect 17743 -10448 17786 -10245
rect 17791 -10448 17798 -10285
rect 17939 -10321 18116 -10287
rect 16495 -10506 17858 -10448
rect 15922 -10543 17858 -10506
rect 17865 -10543 17872 -10359
rect 17877 -10543 17920 -10371
rect 17923 -10543 17931 -10360
rect 18124 -10371 18132 -10360
rect 18135 -10543 18178 -10371
rect 18183 -10543 18190 -10359
rect 18257 -10543 18264 -10285
rect 18269 -10543 18312 -10245
rect 19313 -10506 19356 -10032
rect 19839 -10036 20522 -10032
rect 19509 -10108 19686 -10074
rect 19447 -10506 19490 -10167
rect 19493 -10506 19501 -10156
rect 19694 -10167 19702 -10156
rect 19705 -10506 19748 -10167
rect 19839 -10448 20581 -10036
rect 20592 -10118 20969 -10084
rect 21053 -10180 21065 -10118
rect 20692 -10256 20869 -10222
rect 20618 -10448 20625 -10294
rect 20630 -10448 20673 -10306
rect 20676 -10448 20684 -10295
rect 20877 -10306 20885 -10295
rect 20888 -10448 20931 -10306
rect 20936 -10448 20943 -10294
rect 21010 -10448 21017 -10220
rect 21022 -10448 21065 -10180
rect 21087 -10245 21099 -10149
rect 21183 -10183 21560 -10149
rect 21087 -10448 21130 -10245
rect 21135 -10448 21142 -10285
rect 21283 -10321 21460 -10287
rect 19839 -10506 21202 -10448
rect 19266 -10543 21202 -10506
rect 21209 -10543 21216 -10359
rect 21221 -10543 21264 -10371
rect 21267 -10543 21275 -10360
rect 21468 -10371 21476 -10360
rect 21479 -10543 21522 -10371
rect 21527 -10543 21534 -10359
rect 21601 -10543 21608 -10285
rect 21613 -10543 21656 -10245
rect 22657 -10506 22700 -10032
rect 23183 -10036 23866 -10032
rect 22853 -10108 23030 -10074
rect 22791 -10506 22834 -10167
rect 22837 -10506 22845 -10156
rect 23038 -10167 23046 -10156
rect 23049 -10506 23092 -10167
rect 23183 -10448 23925 -10036
rect 23936 -10118 24313 -10084
rect 24397 -10180 24409 -10118
rect 24036 -10256 24213 -10222
rect 23962 -10448 23969 -10294
rect 23974 -10448 24017 -10306
rect 24020 -10448 24028 -10295
rect 24221 -10306 24229 -10295
rect 24232 -10448 24275 -10306
rect 24280 -10448 24287 -10294
rect 24354 -10448 24361 -10220
rect 24366 -10448 24409 -10180
rect 24431 -10245 24443 -10149
rect 24527 -10183 24904 -10149
rect 24431 -10448 24474 -10245
rect 24479 -10448 24486 -10285
rect 24627 -10321 24804 -10287
rect 23183 -10506 24546 -10448
rect 22610 -10543 24546 -10506
rect 24553 -10543 24560 -10359
rect 24565 -10543 24608 -10371
rect 24611 -10543 24619 -10360
rect 24812 -10371 24820 -10360
rect 24823 -10543 24866 -10371
rect 24871 -10543 24878 -10359
rect 24945 -10543 24952 -10285
rect 24957 -10543 25000 -10245
rect 26001 -10506 26044 -10032
rect 26527 -10036 27210 -10032
rect 26197 -10108 26374 -10074
rect 26135 -10506 26178 -10167
rect 26181 -10506 26189 -10156
rect 26382 -10167 26390 -10156
rect 26393 -10506 26436 -10167
rect 26527 -10448 27269 -10036
rect 27280 -10118 27657 -10084
rect 27741 -10180 27753 -10118
rect 27380 -10256 27557 -10222
rect 27306 -10448 27313 -10294
rect 27318 -10448 27361 -10306
rect 27364 -10448 27372 -10295
rect 27565 -10306 27573 -10295
rect 27576 -10448 27619 -10306
rect 27624 -10448 27631 -10294
rect 27698 -10448 27705 -10220
rect 27710 -10448 27753 -10180
rect 27775 -10245 27787 -10149
rect 27871 -10183 28248 -10149
rect 27775 -10448 27818 -10245
rect 27823 -10448 27830 -10285
rect 27971 -10321 28148 -10287
rect 26527 -10506 27890 -10448
rect 25954 -10543 27890 -10506
rect 27897 -10543 27904 -10359
rect 27909 -10543 27952 -10371
rect 27955 -10543 27963 -10360
rect 28156 -10371 28164 -10360
rect 28167 -10543 28210 -10371
rect 28215 -10543 28222 -10359
rect 28289 -10543 28296 -10285
rect 28301 -10543 28344 -10245
rect 29346 -10506 29388 -10032
rect 29872 -10036 30554 -10032
rect 29542 -10108 29718 -10074
rect 29480 -10506 29522 -10167
rect 29526 -10506 29533 -10156
rect 29727 -10167 29734 -10156
rect 29738 -10506 29780 -10167
rect 29872 -10448 30613 -10036
rect 30625 -10118 31001 -10084
rect 31086 -10180 31097 -10118
rect 30725 -10256 30901 -10222
rect 30651 -10448 30657 -10294
rect 30663 -10448 30705 -10306
rect 30709 -10448 30716 -10295
rect 30910 -10306 30917 -10295
rect 30921 -10448 30963 -10306
rect 30969 -10448 30975 -10294
rect 31043 -10448 31049 -10220
rect 31055 -10448 31097 -10180
rect 31120 -10245 31131 -10149
rect 31216 -10183 31592 -10149
rect 31120 -10448 31162 -10245
rect 31168 -10448 31174 -10285
rect 31316 -10321 31492 -10287
rect 29872 -10506 31234 -10448
rect 29299 -10543 31234 -10506
rect 31242 -10543 31248 -10359
rect 31254 -10543 31296 -10371
rect 31300 -10543 31307 -10360
rect 31501 -10371 31508 -10360
rect 31512 -10543 31554 -10371
rect 31560 -10543 31566 -10359
rect 31634 -10543 31640 -10285
rect 31646 -10543 31688 -10245
rect 32690 -10506 32732 -10032
rect 33216 -10036 33898 -10032
rect 32886 -10108 33062 -10074
rect 32824 -10506 32866 -10167
rect 32870 -10506 32877 -10156
rect 33071 -10167 33078 -10156
rect 33082 -10506 33124 -10167
rect 33216 -10448 33957 -10036
rect 33969 -10118 34345 -10084
rect 34430 -10180 34441 -10118
rect 34069 -10256 34245 -10222
rect 33995 -10448 34001 -10294
rect 34007 -10448 34049 -10306
rect 34053 -10448 34060 -10295
rect 34254 -10306 34261 -10295
rect 34265 -10448 34307 -10306
rect 34313 -10448 34319 -10294
rect 34387 -10448 34393 -10220
rect 34399 -10448 34441 -10180
rect 34464 -10245 34475 -10149
rect 34560 -10183 34936 -10149
rect 34464 -10448 34506 -10245
rect 34512 -10448 34518 -10285
rect 34660 -10321 34836 -10287
rect 33216 -10506 34578 -10448
rect 32643 -10543 34578 -10506
rect 34586 -10543 34592 -10359
rect 34598 -10543 34640 -10371
rect 34644 -10543 34651 -10360
rect 34845 -10371 34852 -10360
rect 34856 -10543 34898 -10371
rect 34904 -10543 34910 -10359
rect 34978 -10543 34984 -10285
rect 34990 -10543 35032 -10245
rect 36034 -10506 36076 -10032
rect 36560 -10036 37242 -10032
rect 36230 -10108 36406 -10074
rect 36168 -10506 36210 -10167
rect 36214 -10506 36221 -10156
rect 36415 -10167 36422 -10156
rect 36426 -10506 36468 -10167
rect 36560 -10448 37301 -10036
rect 37313 -10118 37689 -10084
rect 37774 -10180 37785 -10118
rect 37413 -10256 37589 -10222
rect 37339 -10448 37345 -10294
rect 37351 -10448 37393 -10306
rect 37397 -10448 37404 -10295
rect 37598 -10306 37605 -10295
rect 37609 -10448 37651 -10306
rect 37657 -10448 37663 -10294
rect 37731 -10448 37737 -10220
rect 37743 -10448 37785 -10180
rect 37808 -10245 37819 -10149
rect 37904 -10183 38280 -10149
rect 37808 -10448 37850 -10245
rect 37856 -10448 37862 -10285
rect 38004 -10321 38180 -10287
rect 36560 -10506 37922 -10448
rect 35987 -10543 37922 -10506
rect 37930 -10543 37936 -10359
rect 37942 -10543 37984 -10371
rect 37988 -10543 37995 -10360
rect 38189 -10371 38196 -10360
rect 38200 -10543 38242 -10371
rect 38248 -10543 38254 -10359
rect 38322 -10543 38328 -10285
rect 38334 -10543 38376 -10245
rect 39378 -10506 39420 -10032
rect 39904 -10036 40586 -10032
rect 39574 -10108 39750 -10074
rect 39512 -10506 39554 -10167
rect 39558 -10506 39565 -10156
rect 39759 -10167 39766 -10156
rect 39770 -10506 39812 -10167
rect 39904 -10448 40645 -10036
rect 40657 -10118 41033 -10084
rect 41118 -10180 41129 -10118
rect 40757 -10256 40933 -10222
rect 40683 -10448 40689 -10294
rect 40695 -10448 40737 -10306
rect 40741 -10448 40748 -10295
rect 40942 -10306 40949 -10295
rect 40953 -10448 40995 -10306
rect 41001 -10448 41007 -10294
rect 41075 -10448 41081 -10220
rect 41087 -10448 41129 -10180
rect 41152 -10245 41163 -10149
rect 41248 -10183 41624 -10149
rect 41152 -10448 41194 -10245
rect 41200 -10448 41206 -10285
rect 41348 -10321 41524 -10287
rect 39904 -10506 41266 -10448
rect 39331 -10543 41266 -10506
rect 41274 -10543 41280 -10359
rect 41286 -10543 41328 -10371
rect 41332 -10543 41339 -10360
rect 41533 -10371 41540 -10360
rect 41544 -10543 41586 -10371
rect 41592 -10543 41598 -10359
rect 41666 -10543 41672 -10285
rect 41678 -10543 41720 -10245
rect 42722 -10506 42764 -10032
rect 43248 -10036 43930 -10032
rect 42918 -10108 43094 -10074
rect 42856 -10506 42898 -10167
rect 42902 -10506 42909 -10156
rect 43103 -10167 43110 -10156
rect 43114 -10506 43156 -10167
rect 43248 -10448 43989 -10036
rect 44001 -10118 44377 -10084
rect 44462 -10180 44473 -10118
rect 44101 -10256 44277 -10222
rect 44027 -10448 44033 -10294
rect 44039 -10448 44081 -10306
rect 44085 -10448 44092 -10295
rect 44286 -10306 44293 -10295
rect 44297 -10448 44339 -10306
rect 44345 -10448 44351 -10294
rect 44419 -10448 44425 -10220
rect 44431 -10448 44473 -10180
rect 44496 -10245 44507 -10149
rect 44592 -10183 44968 -10149
rect 44496 -10448 44538 -10245
rect 44544 -10448 44550 -10285
rect 44692 -10321 44868 -10287
rect 43248 -10506 44610 -10448
rect 42675 -10543 44610 -10506
rect 44618 -10543 44624 -10359
rect 44630 -10543 44672 -10371
rect 44676 -10543 44683 -10360
rect 44877 -10371 44884 -10360
rect 44888 -10543 44930 -10371
rect 44936 -10543 44942 -10359
rect 45010 -10543 45016 -10285
rect 45022 -10543 45064 -10245
rect 46066 -10506 46108 -10032
rect 46592 -10036 47274 -10032
rect 46262 -10108 46438 -10074
rect 46200 -10506 46242 -10167
rect 46246 -10506 46253 -10156
rect 46447 -10167 46454 -10156
rect 46458 -10506 46500 -10167
rect 46592 -10448 47333 -10036
rect 47345 -10118 47721 -10084
rect 47806 -10180 47817 -10118
rect 47445 -10256 47621 -10222
rect 47371 -10448 47377 -10294
rect 47383 -10448 47425 -10306
rect 47429 -10448 47436 -10295
rect 47630 -10306 47637 -10295
rect 47641 -10448 47683 -10306
rect 47689 -10448 47695 -10294
rect 47763 -10448 47769 -10220
rect 47775 -10448 47817 -10180
rect 47840 -10245 47851 -10149
rect 47936 -10183 48312 -10149
rect 47840 -10448 47882 -10245
rect 47888 -10448 47894 -10285
rect 48036 -10321 48212 -10287
rect 46592 -10506 47954 -10448
rect 46019 -10543 47954 -10506
rect 47962 -10543 47968 -10359
rect 47974 -10543 48016 -10371
rect 48020 -10543 48027 -10360
rect 48221 -10371 48228 -10360
rect 48232 -10543 48274 -10371
rect 48280 -10543 48286 -10359
rect 48354 -10543 48360 -10285
rect 48366 -10543 48408 -10245
rect 49410 -10506 49452 -10032
rect 49936 -10036 50618 -10032
rect 49606 -10108 49782 -10074
rect 49544 -10506 49586 -10167
rect 49590 -10506 49597 -10156
rect 49791 -10167 49798 -10156
rect 49802 -10506 49844 -10167
rect 49936 -10448 50677 -10036
rect 50689 -10118 51065 -10084
rect 51150 -10180 51161 -10118
rect 50789 -10256 50965 -10222
rect 50715 -10448 50721 -10294
rect 50727 -10448 50769 -10306
rect 50773 -10448 50780 -10295
rect 50974 -10306 50981 -10295
rect 50985 -10448 51027 -10306
rect 51033 -10448 51039 -10294
rect 51107 -10448 51113 -10220
rect 51119 -10448 51161 -10180
rect 51184 -10245 51195 -10149
rect 51280 -10183 51656 -10149
rect 51184 -10448 51226 -10245
rect 51232 -10448 51238 -10285
rect 51380 -10321 51556 -10287
rect 49936 -10506 51298 -10448
rect 49363 -10543 51298 -10506
rect 51306 -10543 51312 -10359
rect 51318 -10543 51360 -10371
rect 51364 -10543 51371 -10360
rect 51565 -10371 51572 -10360
rect 51576 -10543 51618 -10371
rect 51624 -10543 51630 -10359
rect 51698 -10543 51704 -10285
rect 51710 -10543 51752 -10245
rect 52754 -10506 52796 -10032
rect 53280 -10036 53962 -10032
rect 52950 -10108 53126 -10074
rect 52888 -10506 52930 -10167
rect 52934 -10506 52941 -10156
rect 53135 -10167 53142 -10156
rect 53146 -10506 53188 -10167
rect 53280 -10448 54021 -10036
rect 54033 -10118 54409 -10084
rect 54494 -10180 54505 -10118
rect 54133 -10256 54309 -10222
rect 54059 -10448 54065 -10294
rect 54071 -10448 54113 -10306
rect 54117 -10448 54124 -10295
rect 54318 -10306 54325 -10295
rect 54329 -10448 54371 -10306
rect 54377 -10448 54383 -10294
rect 54451 -10448 54457 -10220
rect 54463 -10448 54505 -10180
rect 54528 -10245 54539 -10149
rect 54624 -10183 55000 -10149
rect 54528 -10448 54570 -10245
rect 54576 -10448 54582 -10285
rect 54724 -10321 54900 -10287
rect 53280 -10506 54642 -10448
rect 52707 -10543 54642 -10506
rect 54650 -10543 54656 -10359
rect 54662 -10543 54704 -10371
rect 54708 -10543 54715 -10360
rect 54909 -10371 54916 -10360
rect 54920 -10543 54962 -10371
rect 54968 -10543 54974 -10359
rect 55042 -10543 55048 -10285
rect 55054 -10543 55096 -10245
rect 56099 -10506 56140 -10032
rect 56625 -10036 57306 -10007
rect 56295 -10108 56470 -10074
rect 56233 -10506 56274 -10167
rect 56279 -10506 56285 -10156
rect 56480 -10167 56486 -10156
rect 56491 -10506 56532 -10167
rect 56625 -10448 57365 -10036
rect 57378 -10118 57753 -10084
rect 57839 -10180 57849 -10118
rect 57478 -10256 57653 -10222
rect 57404 -10448 57409 -10294
rect 57416 -10448 57457 -10306
rect 57462 -10448 57468 -10295
rect 57663 -10306 57669 -10295
rect 57674 -10448 57715 -10306
rect 57722 -10448 57727 -10294
rect 57796 -10448 57801 -10220
rect 57808 -10448 57849 -10180
rect 57873 -10245 57883 -10149
rect 57969 -10183 58344 -10149
rect 57873 -10448 57914 -10245
rect 57921 -10448 57926 -10285
rect 58069 -10321 58244 -10287
rect 56625 -10506 57986 -10448
rect 56052 -10543 57986 -10506
rect 57995 -10543 58000 -10359
rect 58007 -10543 58048 -10371
rect 58053 -10543 58059 -10360
rect 58254 -10371 58260 -10360
rect 58265 -10543 58306 -10371
rect 58313 -10543 58318 -10359
rect 58387 -10543 58392 -10285
rect 58399 -10543 58440 -10245
rect 59443 -10506 59484 -10032
rect 59969 -10036 60650 -10007
rect 59639 -10108 59814 -10074
rect 59577 -10506 59618 -10167
rect 59623 -10506 59629 -10156
rect 59824 -10167 59830 -10156
rect 59835 -10506 59876 -10167
rect 59969 -10448 60709 -10036
rect 60722 -10118 61097 -10084
rect 61183 -10180 61193 -10118
rect 60822 -10256 60997 -10222
rect 60748 -10448 60753 -10294
rect 60760 -10448 60801 -10306
rect 60806 -10448 60812 -10295
rect 61007 -10306 61013 -10295
rect 61018 -10448 61059 -10306
rect 61066 -10448 61071 -10294
rect 61140 -10448 61145 -10220
rect 61152 -10448 61193 -10180
rect 61217 -10245 61227 -10149
rect 61313 -10183 61688 -10149
rect 61217 -10448 61258 -10245
rect 61265 -10448 61270 -10285
rect 61413 -10321 61588 -10287
rect 59969 -10506 61330 -10448
rect 59396 -10543 61330 -10506
rect 61339 -10543 61344 -10359
rect 61351 -10543 61392 -10371
rect 61397 -10543 61403 -10360
rect 61598 -10371 61604 -10360
rect 61609 -10543 61650 -10371
rect 61657 -10543 61662 -10359
rect 61731 -10543 61736 -10285
rect 61743 -10543 61784 -10245
rect 62787 -10506 62828 -10032
rect 63313 -10036 63994 -10007
rect 62983 -10108 63158 -10074
rect 62921 -10506 62962 -10167
rect 62967 -10506 62973 -10156
rect 63168 -10167 63174 -10156
rect 63179 -10506 63220 -10167
rect 63313 -10448 64053 -10036
rect 64066 -10118 64441 -10084
rect 64527 -10180 64537 -10118
rect 64166 -10256 64341 -10222
rect 64092 -10448 64097 -10294
rect 64104 -10448 64145 -10306
rect 64150 -10448 64156 -10295
rect 64351 -10306 64357 -10295
rect 64362 -10448 64403 -10306
rect 64410 -10448 64415 -10294
rect 64484 -10448 64489 -10220
rect 64496 -10448 64537 -10180
rect 64561 -10245 64571 -10149
rect 64657 -10183 65032 -10149
rect 64561 -10448 64602 -10245
rect 64609 -10448 64614 -10285
rect 64757 -10321 64932 -10287
rect 63313 -10506 64674 -10448
rect 62740 -10543 64674 -10506
rect 64683 -10543 64688 -10359
rect 64695 -10543 64736 -10371
rect 64741 -10543 64747 -10360
rect 64942 -10371 64948 -10360
rect 64953 -10543 64994 -10371
rect 65001 -10543 65006 -10359
rect 65075 -10543 65080 -10285
rect 65087 -10543 65128 -10245
rect 66131 -10506 66172 -10032
rect 66657 -10036 67338 -10007
rect 66327 -10108 66502 -10074
rect 66265 -10506 66306 -10167
rect 66311 -10506 66317 -10156
rect 66512 -10167 66518 -10156
rect 66523 -10506 66564 -10167
rect 66657 -10448 67397 -10036
rect 67410 -10118 67785 -10084
rect 67871 -10180 67881 -10118
rect 67510 -10256 67685 -10222
rect 67436 -10448 67441 -10294
rect 67448 -10448 67489 -10306
rect 67494 -10448 67500 -10295
rect 67695 -10306 67701 -10295
rect 67706 -10448 67747 -10306
rect 67754 -10448 67759 -10294
rect 67828 -10448 67833 -10220
rect 67840 -10448 67881 -10180
rect 67905 -10245 67915 -10149
rect 68001 -10183 68376 -10149
rect 67905 -10448 67946 -10245
rect 67953 -10448 67958 -10285
rect 68101 -10321 68276 -10287
rect 66657 -10506 68018 -10448
rect 66084 -10543 68018 -10506
rect 68027 -10543 68032 -10359
rect 68039 -10543 68080 -10371
rect 68085 -10543 68091 -10360
rect 68286 -10371 68292 -10360
rect 68297 -10543 68338 -10371
rect 68345 -10543 68350 -10359
rect 68419 -10543 68424 -10285
rect 68431 -10543 68472 -10245
rect 69475 -10506 69516 -10032
rect 70001 -10036 70682 -10007
rect 69671 -10108 69846 -10074
rect 69609 -10506 69650 -10167
rect 69655 -10506 69661 -10156
rect 69856 -10167 69862 -10156
rect 69867 -10506 69908 -10167
rect 70001 -10448 70741 -10036
rect 70754 -10118 71129 -10084
rect 71215 -10180 71225 -10118
rect 70854 -10256 71029 -10222
rect 70780 -10448 70785 -10294
rect 70792 -10448 70833 -10306
rect 70838 -10448 70844 -10295
rect 71039 -10306 71045 -10295
rect 71050 -10448 71091 -10306
rect 71098 -10448 71103 -10294
rect 71172 -10448 71177 -10220
rect 71184 -10448 71225 -10180
rect 71249 -10245 71259 -10149
rect 71345 -10183 71720 -10149
rect 71249 -10448 71290 -10245
rect 71297 -10448 71302 -10285
rect 71445 -10321 71620 -10287
rect 70001 -10506 71362 -10448
rect 69428 -10543 71362 -10506
rect 71371 -10543 71376 -10359
rect 71383 -10543 71424 -10371
rect 71429 -10543 71435 -10360
rect 71630 -10371 71636 -10360
rect 71641 -10543 71682 -10371
rect 71689 -10543 71694 -10359
rect 71763 -10543 71768 -10285
rect 71775 -10543 71816 -10245
rect 72819 -10506 72860 -10032
rect 73345 -10036 74026 -10007
rect 73015 -10108 73190 -10074
rect 72953 -10506 72994 -10167
rect 72999 -10506 73005 -10156
rect 73200 -10167 73206 -10156
rect 73211 -10506 73252 -10167
rect 73345 -10448 74085 -10036
rect 74098 -10118 74473 -10084
rect 74559 -10180 74569 -10118
rect 74198 -10256 74373 -10222
rect 74124 -10448 74129 -10294
rect 74136 -10448 74177 -10306
rect 74182 -10448 74188 -10295
rect 74383 -10306 74389 -10295
rect 74394 -10448 74435 -10306
rect 74442 -10448 74447 -10294
rect 74516 -10448 74521 -10220
rect 74528 -10448 74569 -10180
rect 74593 -10245 74603 -10149
rect 74689 -10183 75064 -10149
rect 74593 -10448 74634 -10245
rect 74641 -10448 74646 -10285
rect 74789 -10321 74964 -10287
rect 73345 -10506 74706 -10448
rect 72772 -10543 74706 -10506
rect 74715 -10543 74720 -10359
rect 74727 -10543 74768 -10371
rect 74773 -10543 74779 -10360
rect 74974 -10371 74980 -10360
rect 74985 -10543 75026 -10371
rect 75033 -10543 75038 -10359
rect 75107 -10543 75112 -10285
rect 75119 -10543 75160 -10245
rect 76163 -10506 76204 -10032
rect 76689 -10036 77370 -10007
rect 76359 -10108 76534 -10074
rect 76297 -10506 76338 -10167
rect 76343 -10506 76349 -10156
rect 76544 -10167 76550 -10156
rect 76555 -10506 76596 -10167
rect 76689 -10448 77429 -10036
rect 77442 -10118 77817 -10084
rect 77903 -10180 77913 -10118
rect 77542 -10256 77717 -10222
rect 77468 -10448 77473 -10294
rect 77480 -10448 77521 -10306
rect 77526 -10448 77532 -10295
rect 77727 -10306 77733 -10295
rect 77738 -10448 77779 -10306
rect 77786 -10448 77791 -10294
rect 77860 -10448 77865 -10220
rect 77872 -10448 77913 -10180
rect 77937 -10245 77947 -10149
rect 78033 -10183 78408 -10149
rect 77937 -10448 77978 -10245
rect 77985 -10448 77990 -10285
rect 78133 -10321 78308 -10287
rect 76689 -10506 78050 -10448
rect 76116 -10543 78050 -10506
rect 78059 -10543 78064 -10359
rect 78071 -10543 78112 -10371
rect 78117 -10543 78123 -10360
rect 78318 -10371 78324 -10360
rect 78329 -10543 78370 -10371
rect 78377 -10543 78382 -10359
rect 78451 -10543 78456 -10285
rect 78463 -10543 78504 -10245
rect 79507 -10506 79548 -10032
rect 80033 -10036 80714 -10007
rect 79703 -10108 79878 -10074
rect 79641 -10506 79682 -10167
rect 79687 -10506 79693 -10156
rect 79888 -10167 79894 -10156
rect 79899 -10506 79940 -10167
rect 80033 -10448 80773 -10036
rect 80786 -10118 81161 -10084
rect 81247 -10180 81257 -10118
rect 80886 -10256 81061 -10222
rect 80812 -10448 80817 -10294
rect 80824 -10448 80865 -10306
rect 80870 -10448 80876 -10295
rect 81071 -10306 81077 -10295
rect 81082 -10448 81123 -10306
rect 81130 -10448 81135 -10294
rect 81204 -10448 81209 -10220
rect 81216 -10448 81257 -10180
rect 81281 -10245 81291 -10149
rect 81377 -10183 81752 -10149
rect 81281 -10448 81322 -10245
rect 81329 -10448 81334 -10285
rect 81477 -10321 81652 -10287
rect 80033 -10506 81394 -10448
rect 79460 -10543 81394 -10506
rect 81403 -10543 81408 -10359
rect 81415 -10543 81456 -10371
rect 81461 -10543 81467 -10360
rect 81662 -10371 81668 -10360
rect 81673 -10543 81714 -10371
rect 81721 -10543 81726 -10359
rect 81795 -10543 81800 -10285
rect 81807 -10543 81848 -10245
rect 82851 -10506 82892 -10032
rect 83377 -10036 84058 -10007
rect 83047 -10108 83222 -10074
rect 82985 -10506 83026 -10167
rect 83031 -10506 83037 -10156
rect 83232 -10167 83238 -10156
rect 83243 -10506 83284 -10167
rect 83377 -10448 84117 -10036
rect 84130 -10118 84505 -10084
rect 84591 -10180 84601 -10118
rect 84230 -10256 84405 -10222
rect 84156 -10448 84161 -10294
rect 84168 -10448 84209 -10306
rect 84214 -10448 84220 -10295
rect 84415 -10306 84421 -10295
rect 84426 -10448 84467 -10306
rect 84474 -10448 84479 -10294
rect 84548 -10448 84553 -10220
rect 84560 -10448 84601 -10180
rect 84625 -10245 84635 -10149
rect 84721 -10183 85096 -10149
rect 84625 -10448 84666 -10245
rect 84673 -10448 84678 -10285
rect 84821 -10321 84996 -10287
rect 83377 -10506 84738 -10448
rect 82804 -10543 84738 -10506
rect 84747 -10543 84752 -10359
rect 84759 -10543 84800 -10371
rect 84805 -10543 84811 -10360
rect 85006 -10371 85012 -10360
rect 85017 -10543 85058 -10371
rect 85065 -10543 85070 -10359
rect 85139 -10543 85144 -10285
rect 85151 -10543 85192 -10245
rect 86195 -10506 86236 -10032
rect 86721 -10036 87402 -10007
rect 86391 -10108 86566 -10074
rect 86329 -10506 86370 -10167
rect 86375 -10506 86381 -10156
rect 86576 -10167 86582 -10156
rect 86587 -10506 86628 -10167
rect 86721 -10448 87461 -10036
rect 87474 -10118 87849 -10084
rect 87935 -10180 87945 -10118
rect 87574 -10256 87749 -10222
rect 87500 -10448 87505 -10294
rect 87512 -10448 87553 -10306
rect 87558 -10448 87564 -10295
rect 87759 -10306 87765 -10295
rect 87770 -10448 87811 -10306
rect 87818 -10448 87823 -10294
rect 87892 -10448 87897 -10220
rect 87904 -10448 87945 -10180
rect 87969 -10245 87979 -10149
rect 88065 -10183 88440 -10149
rect 87969 -10448 88010 -10245
rect 88017 -10448 88022 -10285
rect 88165 -10321 88340 -10287
rect 86721 -10506 88082 -10448
rect 86148 -10543 88082 -10506
rect 88091 -10543 88096 -10359
rect 88103 -10543 88144 -10371
rect 88149 -10543 88155 -10360
rect 88350 -10371 88356 -10360
rect 88361 -10543 88402 -10371
rect 88409 -10543 88414 -10359
rect 88483 -10543 88488 -10285
rect 88495 -10543 88536 -10245
rect 89539 -10506 89580 -10032
rect 90065 -10036 90746 -10007
rect 89735 -10108 89910 -10074
rect 89673 -10506 89714 -10167
rect 89719 -10506 89725 -10156
rect 89920 -10167 89926 -10156
rect 89931 -10506 89972 -10167
rect 90065 -10448 90805 -10036
rect 90818 -10118 91193 -10084
rect 91279 -10180 91289 -10118
rect 90918 -10256 91093 -10222
rect 90844 -10448 90849 -10294
rect 90856 -10448 90897 -10306
rect 90902 -10448 90908 -10295
rect 91103 -10306 91109 -10295
rect 91114 -10448 91155 -10306
rect 91162 -10448 91167 -10294
rect 91236 -10448 91241 -10220
rect 91248 -10448 91289 -10180
rect 91313 -10245 91323 -10149
rect 91409 -10183 91784 -10149
rect 91313 -10448 91354 -10245
rect 91361 -10448 91366 -10285
rect 91509 -10321 91684 -10287
rect 90065 -10506 91426 -10448
rect 89492 -10543 91426 -10506
rect 91435 -10543 91440 -10359
rect 91447 -10543 91488 -10371
rect 91493 -10543 91499 -10360
rect 91694 -10371 91700 -10360
rect 91705 -10543 91746 -10371
rect 91753 -10543 91758 -10359
rect 91827 -10543 91832 -10285
rect 91839 -10543 91880 -10245
rect 92883 -10506 92924 -10032
rect 93409 -10036 94090 -10007
rect 93079 -10108 93254 -10074
rect 93017 -10506 93058 -10167
rect 93063 -10506 93069 -10156
rect 93264 -10167 93270 -10156
rect 93275 -10506 93316 -10167
rect 93409 -10448 94149 -10036
rect 94162 -10118 94537 -10084
rect 94623 -10180 94633 -10118
rect 94262 -10256 94437 -10222
rect 94188 -10448 94193 -10294
rect 94200 -10448 94241 -10306
rect 94246 -10448 94252 -10295
rect 94447 -10306 94453 -10295
rect 94458 -10448 94499 -10306
rect 94506 -10448 94511 -10294
rect 94580 -10448 94585 -10220
rect 94592 -10448 94633 -10180
rect 94657 -10245 94667 -10149
rect 94753 -10183 95128 -10149
rect 94657 -10448 94698 -10245
rect 94705 -10448 94710 -10285
rect 94853 -10321 95028 -10287
rect 93409 -10506 94770 -10448
rect 92836 -10543 94770 -10506
rect 94779 -10543 94784 -10359
rect 94791 -10543 94832 -10371
rect 94837 -10543 94843 -10360
rect 95038 -10371 95044 -10360
rect 95049 -10543 95090 -10371
rect 95097 -10543 95102 -10359
rect 95171 -10543 95176 -10285
rect 95183 -10543 95224 -10245
rect 96227 -10506 96268 -10032
rect 96753 -10036 97434 -10007
rect 96423 -10108 96598 -10074
rect 96361 -10506 96402 -10167
rect 96407 -10506 96413 -10156
rect 96608 -10167 96614 -10156
rect 96619 -10506 96660 -10167
rect 96753 -10448 97493 -10036
rect 97506 -10118 97881 -10084
rect 97967 -10180 97977 -10118
rect 97606 -10256 97781 -10222
rect 97532 -10448 97537 -10294
rect 97544 -10448 97585 -10306
rect 97590 -10448 97596 -10295
rect 97791 -10306 97797 -10295
rect 97802 -10448 97843 -10306
rect 97850 -10448 97855 -10294
rect 97924 -10448 97929 -10220
rect 97936 -10448 97977 -10180
rect 98001 -10245 98011 -10149
rect 98097 -10183 98472 -10149
rect 98001 -10448 98042 -10245
rect 98049 -10448 98054 -10285
rect 98197 -10321 98372 -10287
rect 96753 -10506 98114 -10448
rect 96180 -10543 98114 -10506
rect 98123 -10543 98128 -10359
rect 98135 -10543 98176 -10371
rect 98181 -10543 98187 -10360
rect 98382 -10371 98388 -10360
rect 98393 -10543 98434 -10371
rect 98441 -10543 98446 -10359
rect 98515 -10543 98520 -10285
rect 98527 -10543 98568 -10245
rect 99571 -10506 99612 -10032
rect 100097 -10036 100778 -10007
rect 99767 -10108 99942 -10074
rect 99705 -10506 99746 -10167
rect 99751 -10506 99757 -10156
rect 99952 -10167 99958 -10156
rect 99963 -10506 100004 -10167
rect 100097 -10448 100837 -10036
rect 100850 -10118 101225 -10084
rect 101311 -10180 101321 -10118
rect 100950 -10256 101125 -10222
rect 100876 -10448 100881 -10294
rect 100888 -10448 100929 -10306
rect 100934 -10448 100940 -10295
rect 101135 -10306 101141 -10295
rect 101146 -10448 101187 -10306
rect 101194 -10448 101199 -10294
rect 101268 -10448 101273 -10220
rect 101280 -10448 101321 -10180
rect 101345 -10245 101355 -10149
rect 101441 -10183 101816 -10149
rect 101345 -10448 101386 -10245
rect 101393 -10448 101398 -10285
rect 101541 -10321 101716 -10287
rect 100097 -10506 101458 -10448
rect 99524 -10543 101458 -10506
rect 101467 -10543 101472 -10359
rect 101479 -10543 101520 -10371
rect 101525 -10543 101531 -10360
rect 101726 -10371 101732 -10360
rect 101737 -10543 101778 -10371
rect 101785 -10543 101790 -10359
rect 101859 -10543 101864 -10285
rect 101871 -10543 101912 -10245
rect 102915 -10506 102956 -10032
rect 103441 -10036 104122 -10007
rect 103111 -10108 103286 -10074
rect 103049 -10506 103090 -10167
rect 103095 -10506 103101 -10156
rect 103296 -10167 103302 -10156
rect 103307 -10506 103348 -10167
rect 103441 -10448 104181 -10036
rect 104194 -10118 104569 -10084
rect 104655 -10180 104665 -10118
rect 104294 -10256 104469 -10222
rect 104220 -10448 104225 -10294
rect 104232 -10448 104273 -10306
rect 104278 -10448 104284 -10295
rect 104479 -10306 104485 -10295
rect 104490 -10448 104531 -10306
rect 104538 -10448 104543 -10294
rect 104612 -10448 104617 -10220
rect 104624 -10448 104665 -10180
rect 104689 -10245 104699 -10149
rect 104785 -10183 105160 -10149
rect 104689 -10448 104730 -10245
rect 104737 -10448 104742 -10285
rect 104885 -10321 105060 -10287
rect 103441 -10506 104802 -10448
rect 102868 -10543 104802 -10506
rect 104811 -10543 104816 -10359
rect 104823 -10543 104864 -10371
rect 104869 -10543 104875 -10360
rect 105070 -10371 105076 -10360
rect 105081 -10543 105122 -10371
rect 105129 -10543 105134 -10359
rect 105203 -10543 105208 -10285
rect 105215 -10543 105256 -10245
rect 106259 -10506 106300 -10032
rect 106785 -10036 107466 -10007
rect 106455 -10108 106630 -10074
rect 106393 -10506 106434 -10167
rect 106439 -10506 106445 -10156
rect 106640 -10167 106646 -10156
rect 106651 -10506 106692 -10167
rect 106785 -10448 107525 -10036
rect 107538 -10118 107913 -10084
rect 107999 -10180 108009 -10118
rect 107638 -10256 107813 -10222
rect 107564 -10448 107569 -10294
rect 107576 -10448 107617 -10306
rect 107622 -10448 107628 -10295
rect 107823 -10306 107829 -10295
rect 107834 -10448 107875 -10306
rect 107882 -10448 107887 -10294
rect 107956 -10448 107961 -10220
rect 107968 -10448 108009 -10180
rect 108033 -10245 108043 -10149
rect 108129 -10183 108504 -10149
rect 108033 -10448 108074 -10245
rect 108081 -10448 108086 -10285
rect 108229 -10321 108404 -10287
rect 106785 -10506 108146 -10448
rect 106212 -10543 108146 -10506
rect 108155 -10543 108160 -10359
rect 108167 -10543 108208 -10371
rect 108213 -10543 108219 -10360
rect 108414 -10371 108420 -10360
rect 108425 -10543 108466 -10371
rect 108473 -10543 108478 -10359
rect 108547 -10543 108552 -10285
rect 108559 -10543 108600 -10245
rect 109609 -10506 109644 -10032
rect 110135 -10036 110810 -10007
rect 109805 -10108 109974 -10074
rect 109743 -10506 109778 -10167
rect 110001 -10506 110036 -10167
rect 110135 -10448 110869 -10036
rect 110888 -10118 111257 -10084
rect 110988 -10256 111157 -10222
rect 110926 -10448 110961 -10306
rect 111184 -10448 111219 -10306
rect 111317 -10448 111365 -10083
rect 111371 -10448 111419 -10137
rect 111479 -10183 111848 -10149
rect 111579 -10321 111748 -10287
rect 110135 -10506 111490 -10448
rect 109562 -10543 111490 -10506
rect 111517 -10543 111552 -10371
rect 111775 -10543 111810 -10371
rect 111909 -10543 111944 -10245
rect 112953 -10506 112988 -10032
rect 113479 -10036 114154 -10007
rect 113149 -10108 113318 -10074
rect 113087 -10506 113122 -10167
rect 113345 -10506 113380 -10167
rect 113479 -10448 114213 -10036
rect 114232 -10118 114601 -10084
rect 114332 -10256 114501 -10222
rect 114270 -10448 114305 -10306
rect 114528 -10448 114563 -10306
rect 114661 -10448 114709 -10083
rect 114715 -10448 114763 -10137
rect 114823 -10183 115192 -10149
rect 114923 -10321 115092 -10287
rect 113479 -10506 114834 -10448
rect 112906 -10543 114834 -10506
rect 114861 -10543 114896 -10371
rect 115119 -10543 115154 -10371
rect 115253 -10543 115288 -10245
rect 116297 -10506 116332 -10032
rect 116823 -10036 117498 -10007
rect 116493 -10108 116662 -10074
rect 116431 -10506 116466 -10167
rect 116689 -10506 116724 -10167
rect 116823 -10448 117557 -10036
rect 117576 -10118 117945 -10084
rect 117676 -10256 117845 -10222
rect 117614 -10448 117649 -10306
rect 117872 -10448 117907 -10306
rect 118005 -10448 118053 -10083
rect 118059 -10448 118107 -10137
rect 118167 -10183 118536 -10149
rect 118267 -10321 118436 -10287
rect 116823 -10506 118178 -10448
rect 116250 -10543 118178 -10506
rect 118205 -10543 118240 -10371
rect 118463 -10543 118498 -10371
rect 118597 -10543 118632 -10245
rect 119641 -10506 119676 -10032
rect 120167 -10036 120842 -10007
rect 119837 -10108 120006 -10074
rect 119775 -10506 119810 -10167
rect 120033 -10506 120068 -10167
rect 120167 -10448 120901 -10036
rect 120920 -10118 121289 -10084
rect 121020 -10256 121189 -10222
rect 120958 -10448 120993 -10306
rect 121216 -10448 121251 -10306
rect 121349 -10448 121397 -10083
rect 121403 -10448 121451 -10137
rect 121511 -10183 121880 -10149
rect 121611 -10321 121780 -10287
rect 120167 -10506 121522 -10448
rect 119594 -10543 121522 -10506
rect 121549 -10543 121584 -10371
rect 121807 -10543 121842 -10371
rect 121941 -10543 121976 -10245
rect 122985 -10506 123020 -10032
rect 123511 -10036 124186 -10007
rect 123181 -10108 123350 -10074
rect 123119 -10506 123154 -10167
rect 123377 -10506 123412 -10167
rect 123511 -10448 124245 -10036
rect 124264 -10118 124633 -10084
rect 124364 -10256 124533 -10222
rect 124302 -10448 124337 -10306
rect 124560 -10448 124595 -10306
rect 124693 -10448 124741 -10083
rect 124747 -10448 124795 -10137
rect 124855 -10183 125224 -10149
rect 124955 -10321 125124 -10287
rect 123511 -10506 124866 -10448
rect 122938 -10543 124866 -10506
rect 124893 -10543 124928 -10371
rect 125151 -10543 125186 -10371
rect 125285 -10543 125320 -10245
rect 126329 -10506 126364 -10032
rect 126855 -10036 127530 -10007
rect 126525 -10108 126694 -10074
rect 126463 -10506 126498 -10167
rect 126721 -10506 126756 -10167
rect 126855 -10448 127589 -10036
rect 127608 -10118 127977 -10084
rect 127708 -10256 127877 -10222
rect 127646 -10448 127681 -10306
rect 127904 -10448 127939 -10306
rect 128037 -10448 128085 -10083
rect 128091 -10448 128139 -10137
rect 128199 -10183 128568 -10149
rect 128299 -10321 128468 -10287
rect 126855 -10506 128210 -10448
rect 126282 -10543 128210 -10506
rect 128237 -10543 128272 -10371
rect 128495 -10543 128530 -10371
rect 128629 -10543 128664 -10245
rect 129673 -10506 129708 -10032
rect 130199 -10036 130874 -10007
rect 129869 -10108 130038 -10074
rect 129807 -10506 129842 -10167
rect 130065 -10506 130100 -10167
rect 130199 -10448 130933 -10036
rect 130952 -10118 131321 -10084
rect 131052 -10256 131221 -10222
rect 130990 -10448 131025 -10306
rect 131248 -10448 131283 -10306
rect 131381 -10448 131429 -10083
rect 131435 -10448 131483 -10137
rect 131543 -10183 131912 -10149
rect 131643 -10321 131812 -10287
rect 130199 -10506 131554 -10448
rect 129626 -10543 131554 -10506
rect 131581 -10543 131616 -10371
rect 131839 -10543 131874 -10371
rect 131973 -10543 132008 -10245
rect 133017 -10506 133052 -10032
rect 133543 -10036 134218 -10007
rect 133213 -10108 133382 -10074
rect 133151 -10506 133186 -10167
rect 133409 -10506 133444 -10167
rect 133543 -10448 134277 -10036
rect 134296 -10118 134665 -10084
rect 134396 -10256 134565 -10222
rect 134334 -10448 134369 -10306
rect 134592 -10448 134627 -10306
rect 134725 -10448 134773 -10083
rect 134779 -10448 134827 -10137
rect 134887 -10183 135256 -10149
rect 134987 -10321 135156 -10287
rect 133543 -10506 134898 -10448
rect 132970 -10543 134898 -10506
rect 134925 -10543 134960 -10371
rect 135183 -10543 135218 -10371
rect 135317 -10543 135352 -10245
rect 136361 -10506 136396 -10032
rect 136887 -10036 137562 -10007
rect 136557 -10108 136726 -10074
rect 136495 -10506 136530 -10167
rect 136753 -10506 136788 -10167
rect 136887 -10448 137621 -10036
rect 137640 -10118 138009 -10084
rect 137740 -10256 137909 -10222
rect 137678 -10448 137713 -10306
rect 137936 -10448 137971 -10306
rect 138069 -10448 138117 -10083
rect 138123 -10448 138171 -10137
rect 138231 -10183 138600 -10149
rect 138331 -10321 138500 -10287
rect 136887 -10506 138242 -10448
rect 136314 -10543 138242 -10506
rect 138269 -10543 138304 -10371
rect 138527 -10543 138562 -10371
rect 138661 -10543 138696 -10245
rect 139705 -10506 139740 -10032
rect 140231 -10036 140906 -10007
rect 139901 -10108 140070 -10074
rect 139839 -10506 139874 -10167
rect 140097 -10506 140132 -10167
rect 140231 -10448 140965 -10036
rect 140984 -10118 141353 -10084
rect 141084 -10256 141253 -10222
rect 141022 -10448 141057 -10306
rect 141280 -10448 141315 -10306
rect 141413 -10448 141461 -10083
rect 141467 -10448 141515 -10137
rect 141575 -10183 141944 -10149
rect 141675 -10321 141844 -10287
rect 140231 -10506 141586 -10448
rect 139658 -10543 141586 -10506
rect 141613 -10543 141648 -10371
rect 141871 -10543 141906 -10371
rect 142005 -10543 142040 -10245
rect 143049 -10506 143084 -10032
rect 143575 -10036 144250 -10007
rect 143245 -10108 143414 -10074
rect 143183 -10506 143218 -10167
rect 143441 -10506 143476 -10167
rect 143575 -10448 144309 -10036
rect 144328 -10118 144697 -10084
rect 144428 -10256 144597 -10222
rect 144366 -10448 144401 -10306
rect 144624 -10448 144659 -10306
rect 144757 -10448 144805 -10083
rect 144811 -10448 144859 -10137
rect 144919 -10183 145288 -10149
rect 145019 -10321 145188 -10287
rect 143575 -10506 144930 -10448
rect 143002 -10543 144930 -10506
rect 144957 -10543 144992 -10371
rect 145215 -10543 145250 -10371
rect 145349 -10543 145384 -10245
rect 146393 -10506 146428 -10032
rect 146919 -10036 147594 -10007
rect 146589 -10108 146758 -10074
rect 146527 -10506 146562 -10167
rect 146785 -10506 146820 -10167
rect 146919 -10448 147653 -10036
rect 147672 -10118 148041 -10084
rect 147772 -10256 147941 -10222
rect 147710 -10448 147745 -10306
rect 147968 -10448 148003 -10306
rect 148101 -10448 148149 -10083
rect 148155 -10448 148203 -10137
rect 148263 -10183 148632 -10149
rect 148363 -10321 148532 -10287
rect 146919 -10506 148274 -10448
rect 146346 -10543 148274 -10506
rect 148301 -10543 148336 -10371
rect 148559 -10543 148594 -10371
rect 148693 -10543 148728 -10245
rect 149737 -10506 149772 -10032
rect 150263 -10036 150938 -10007
rect 149933 -10108 150102 -10074
rect 149871 -10506 149906 -10167
rect 150129 -10506 150164 -10167
rect 150263 -10448 150997 -10036
rect 151016 -10118 151385 -10084
rect 151116 -10256 151285 -10222
rect 151054 -10448 151089 -10306
rect 151312 -10448 151347 -10306
rect 151445 -10448 151493 -10083
rect 151499 -10448 151547 -10137
rect 151607 -10183 151976 -10149
rect 151707 -10321 151876 -10287
rect 150263 -10506 151618 -10448
rect 149690 -10543 151618 -10506
rect 151645 -10543 151680 -10371
rect 151903 -10543 151938 -10371
rect 152037 -10543 152072 -10245
rect 153081 -10506 153116 -10032
rect 153607 -10036 154282 -10007
rect 153277 -10108 153446 -10074
rect 153215 -10506 153250 -10167
rect 153473 -10506 153508 -10167
rect 153607 -10448 154341 -10036
rect 154360 -10118 154729 -10084
rect 154460 -10256 154629 -10222
rect 154398 -10448 154433 -10306
rect 154656 -10448 154691 -10306
rect 154789 -10448 154837 -10083
rect 154843 -10448 154891 -10137
rect 154951 -10183 155320 -10149
rect 155051 -10321 155220 -10287
rect 153607 -10506 154962 -10448
rect 153034 -10543 154962 -10506
rect 154989 -10543 155024 -10371
rect 155247 -10543 155282 -10371
rect 155381 -10543 155416 -10245
rect 156425 -10506 156460 -10032
rect 156951 -10036 157626 -10007
rect 156621 -10108 156790 -10074
rect 156559 -10506 156594 -10167
rect 156817 -10506 156852 -10167
rect 156951 -10448 157685 -10036
rect 157704 -10118 158073 -10084
rect 157804 -10256 157973 -10222
rect 157742 -10448 157777 -10306
rect 158000 -10448 158035 -10306
rect 158133 -10448 158181 -10083
rect 158187 -10448 158235 -10137
rect 158295 -10183 158664 -10149
rect 158395 -10321 158564 -10287
rect 156951 -10506 158306 -10448
rect 156378 -10543 158306 -10506
rect 158333 -10543 158368 -10371
rect 158591 -10543 158626 -10371
rect 158725 -10543 158760 -10245
rect 159769 -10506 159804 -10032
rect 160295 -10036 160970 -10007
rect 159965 -10108 160134 -10074
rect 159903 -10506 159938 -10167
rect 160161 -10506 160196 -10167
rect 160295 -10448 161029 -10036
rect 161048 -10118 161417 -10084
rect 161148 -10256 161317 -10222
rect 161086 -10448 161121 -10306
rect 161344 -10448 161379 -10306
rect 161477 -10448 161525 -10083
rect 161531 -10448 161579 -10137
rect 161639 -10183 162008 -10149
rect 161739 -10321 161908 -10287
rect 160295 -10506 161650 -10448
rect 159722 -10543 161650 -10506
rect 161677 -10543 161712 -10371
rect 161935 -10543 161970 -10371
rect 162069 -10543 162104 -10245
rect 163113 -10506 163148 -10032
rect 163639 -10036 164314 -10007
rect 163309 -10108 163478 -10074
rect 163247 -10506 163282 -10167
rect 163505 -10506 163540 -10167
rect 163639 -10448 164373 -10036
rect 164392 -10118 164761 -10084
rect 164492 -10256 164661 -10222
rect 164430 -10448 164465 -10306
rect 164688 -10448 164723 -10306
rect 164821 -10448 164869 -10083
rect 164875 -10448 164923 -10137
rect 164983 -10183 165352 -10149
rect 165083 -10321 165252 -10287
rect 163639 -10506 164994 -10448
rect 163066 -10543 164994 -10506
rect 165021 -10543 165056 -10371
rect 165279 -10543 165314 -10371
rect 165413 -10543 165448 -10245
rect 166457 -10506 166492 -10032
rect 166983 -10036 167658 -10007
rect 166653 -10108 166822 -10074
rect 166591 -10506 166626 -10167
rect 166849 -10506 166884 -10167
rect 166983 -10448 167717 -10036
rect 167736 -10118 168105 -10084
rect 167836 -10256 168005 -10222
rect 167774 -10448 167809 -10306
rect 168032 -10448 168067 -10306
rect 168165 -10448 168213 -10083
rect 168219 -10448 168267 -10137
rect 168327 -10183 168696 -10149
rect 168427 -10321 168596 -10287
rect 166983 -10506 168338 -10448
rect 166410 -10543 168338 -10506
rect 168365 -10543 168400 -10371
rect 168623 -10543 168658 -10371
rect 168757 -10543 168792 -10245
rect 169801 -10506 169836 -10032
rect 170327 -10036 171002 -10007
rect 169997 -10108 170166 -10074
rect 169935 -10506 169970 -10167
rect 170193 -10506 170228 -10167
rect 170327 -10448 171061 -10036
rect 171080 -10118 171449 -10084
rect 171180 -10256 171349 -10222
rect 171118 -10448 171153 -10306
rect 171376 -10448 171411 -10306
rect 171509 -10448 171557 -10083
rect 171563 -10448 171611 -10137
rect 171671 -10183 172040 -10149
rect 171771 -10321 171940 -10287
rect 170327 -10506 171682 -10448
rect 169754 -10543 171682 -10506
rect 171709 -10543 171744 -10371
rect 171967 -10543 172002 -10371
rect 172101 -10543 172136 -10245
rect 173145 -10506 173180 -10032
rect 173671 -10036 174346 -10007
rect 173341 -10108 173510 -10074
rect 173279 -10506 173314 -10167
rect 173537 -10506 173572 -10167
rect 173671 -10448 174405 -10036
rect 174424 -10118 174793 -10084
rect 174524 -10256 174693 -10222
rect 174462 -10448 174497 -10306
rect 174720 -10448 174755 -10306
rect 174853 -10448 174901 -10083
rect 174907 -10448 174955 -10137
rect 175015 -10183 175384 -10149
rect 175115 -10321 175284 -10287
rect 173671 -10506 175026 -10448
rect 173098 -10543 175026 -10506
rect 175053 -10543 175088 -10371
rect 175311 -10543 175346 -10371
rect 175445 -10543 175480 -10245
rect 176489 -10506 176524 -10032
rect 177015 -10036 177690 -10007
rect 176685 -10108 176854 -10074
rect 176623 -10506 176658 -10167
rect 176881 -10506 176916 -10167
rect 177015 -10448 177749 -10036
rect 177768 -10118 178137 -10084
rect 177868 -10256 178037 -10222
rect 177806 -10448 177841 -10306
rect 178064 -10448 178099 -10306
rect 178197 -10448 178245 -10083
rect 178251 -10448 178299 -10137
rect 178359 -10183 178728 -10149
rect 178459 -10321 178628 -10287
rect 177015 -10506 178370 -10448
rect 176442 -10543 178370 -10506
rect 178397 -10543 178432 -10371
rect 178655 -10543 178690 -10371
rect 178789 -10543 178824 -10245
rect 179833 -10506 179868 -10032
rect 180359 -10036 181034 -10007
rect 180029 -10108 180198 -10074
rect 179967 -10506 180002 -10167
rect 180225 -10506 180260 -10167
rect 180359 -10448 181093 -10036
rect 181112 -10118 181481 -10084
rect 181212 -10256 181381 -10222
rect 181150 -10448 181185 -10306
rect 181408 -10448 181443 -10306
rect 181541 -10448 181589 -10083
rect 181595 -10448 181643 -10137
rect 181703 -10183 182072 -10149
rect 181803 -10321 181972 -10287
rect 180359 -10506 181714 -10448
rect 179786 -10543 181714 -10506
rect 181741 -10543 181776 -10371
rect 181999 -10543 182034 -10371
rect 182133 -10543 182168 -10245
rect 183177 -10506 183212 -10032
rect 183703 -10036 184378 -10007
rect 183373 -10108 183542 -10074
rect 183311 -10506 183346 -10167
rect 183569 -10506 183604 -10167
rect 183703 -10448 184437 -10036
rect 184456 -10118 184825 -10084
rect 184556 -10256 184725 -10222
rect 184494 -10448 184529 -10306
rect 184752 -10448 184787 -10306
rect 184885 -10448 184933 -10083
rect 184939 -10448 184987 -10137
rect 185047 -10183 185416 -10149
rect 185147 -10321 185316 -10287
rect 183703 -10506 185058 -10448
rect 183130 -10543 185058 -10506
rect 185085 -10543 185120 -10371
rect 185343 -10543 185378 -10371
rect 185477 -10543 185512 -10245
rect 186521 -10506 186556 -10032
rect 187047 -10036 187722 -10007
rect 186717 -10108 186886 -10074
rect 186655 -10506 186690 -10167
rect 186913 -10506 186948 -10167
rect 187047 -10448 187781 -10036
rect 187800 -10118 188169 -10084
rect 187900 -10256 188069 -10222
rect 187838 -10448 187873 -10306
rect 188096 -10448 188131 -10306
rect 188229 -10448 188277 -10083
rect 188283 -10448 188331 -10137
rect 188391 -10183 188760 -10149
rect 188491 -10321 188660 -10287
rect 187047 -10506 188402 -10448
rect 186474 -10543 188402 -10506
rect 188429 -10543 188464 -10371
rect 188687 -10543 188722 -10371
rect 188821 -10543 188856 -10245
rect 189865 -10506 189900 -10032
rect 190391 -10036 191066 -10007
rect 190061 -10108 190230 -10074
rect 189999 -10506 190034 -10167
rect 190257 -10506 190292 -10167
rect 190391 -10448 191125 -10036
rect 191144 -10118 191513 -10084
rect 191244 -10256 191413 -10222
rect 191182 -10448 191217 -10306
rect 191440 -10448 191475 -10306
rect 191573 -10448 191621 -10083
rect 191627 -10448 191675 -10137
rect 191735 -10183 192104 -10149
rect 191835 -10321 192004 -10287
rect 190391 -10506 191746 -10448
rect 189818 -10543 191746 -10506
rect 191773 -10543 191808 -10371
rect 192031 -10543 192066 -10371
rect 192165 -10543 192200 -10245
rect 193209 -10506 193244 -10032
rect 193735 -10036 194410 -10007
rect 193405 -10108 193574 -10074
rect 193343 -10506 193378 -10167
rect 193601 -10506 193636 -10167
rect 193735 -10448 194469 -10036
rect 194488 -10118 194857 -10084
rect 194588 -10256 194757 -10222
rect 194526 -10448 194561 -10306
rect 194784 -10448 194819 -10306
rect 194917 -10448 194965 -10083
rect 194971 -10448 195019 -10137
rect 195079 -10183 195448 -10149
rect 195179 -10321 195348 -10287
rect 193735 -10506 195090 -10448
rect 193162 -10543 195090 -10506
rect 195117 -10543 195152 -10371
rect 195375 -10543 195410 -10371
rect 195509 -10543 195544 -10245
rect 196553 -10506 196588 -10032
rect 197079 -10036 197754 -10007
rect 196749 -10108 196918 -10074
rect 196687 -10506 196722 -10167
rect 196945 -10506 196980 -10167
rect 197079 -10448 197813 -10036
rect 197832 -10118 198201 -10084
rect 197932 -10256 198101 -10222
rect 197870 -10448 197905 -10306
rect 198128 -10448 198163 -10306
rect 198261 -10448 198309 -10083
rect 198315 -10448 198363 -10137
rect 198423 -10183 198792 -10149
rect 198523 -10321 198692 -10287
rect 197079 -10506 198434 -10448
rect 196506 -10543 198434 -10506
rect 198461 -10543 198496 -10371
rect 198719 -10543 198754 -10371
rect 198853 -10543 198888 -10245
rect 199897 -10506 199932 -10032
rect 200423 -10036 201098 -10007
rect 200093 -10108 200262 -10074
rect 200031 -10506 200066 -10167
rect 200289 -10506 200324 -10167
rect 200423 -10448 201157 -10036
rect 201176 -10118 201545 -10084
rect 201276 -10256 201445 -10222
rect 201214 -10448 201249 -10306
rect 201472 -10448 201507 -10306
rect 201605 -10448 201653 -10083
rect 201659 -10448 201707 -10137
rect 201767 -10183 202136 -10149
rect 201867 -10321 202036 -10287
rect 200423 -10506 201778 -10448
rect 199850 -10543 201778 -10506
rect 201805 -10543 201840 -10371
rect 202063 -10543 202098 -10371
rect 202197 -10543 202232 -10245
rect 203241 -10506 203276 -10032
rect 203767 -10036 204442 -10007
rect 203437 -10108 203606 -10074
rect 203375 -10506 203410 -10167
rect 203633 -10506 203668 -10167
rect 203767 -10448 204501 -10036
rect 204520 -10118 204889 -10084
rect 204620 -10256 204789 -10222
rect 204558 -10448 204593 -10306
rect 204816 -10448 204851 -10306
rect 204949 -10448 204997 -10083
rect 205003 -10448 205051 -10137
rect 205111 -10183 205480 -10149
rect 205211 -10321 205380 -10287
rect 203767 -10506 205122 -10448
rect 203194 -10543 205122 -10506
rect 205149 -10543 205184 -10371
rect 205407 -10543 205442 -10371
rect 205541 -10543 205576 -10245
rect 206585 -10506 206620 -10032
rect 207111 -10036 207786 -10007
rect 206781 -10108 206950 -10074
rect 206719 -10506 206754 -10167
rect 206977 -10506 207012 -10167
rect 207111 -10448 207845 -10036
rect 207864 -10118 208233 -10084
rect 207964 -10256 208133 -10222
rect 207902 -10448 207937 -10306
rect 208160 -10448 208195 -10306
rect 208293 -10448 208341 -10083
rect 208347 -10448 208395 -10137
rect 208455 -10183 208824 -10149
rect 208555 -10321 208724 -10287
rect 207111 -10506 208466 -10448
rect 206538 -10543 208466 -10506
rect 208493 -10543 208528 -10371
rect 208751 -10543 208786 -10371
rect 208885 -10543 208920 -10245
rect 209929 -10506 209964 -10032
rect 210455 -10036 211130 -10007
rect 210125 -10108 210294 -10074
rect 210063 -10506 210098 -10167
rect 210321 -10506 210356 -10167
rect 210455 -10448 211189 -10036
rect 211208 -10118 211577 -10084
rect 211308 -10256 211477 -10222
rect 211246 -10448 211281 -10306
rect 211504 -10448 211539 -10306
rect 211637 -10448 211685 -10083
rect 211691 -10448 211739 -10137
rect 211799 -10183 212168 -10149
rect 211899 -10321 212068 -10287
rect 210455 -10506 211810 -10448
rect 209882 -10543 211810 -10506
rect 211837 -10543 211872 -10371
rect 212095 -10543 212130 -10371
rect 212229 -10543 212264 -10245
rect 213273 -10506 213308 -10032
rect 213799 -10036 214474 -10007
rect 213469 -10108 213638 -10074
rect 213407 -10506 213442 -10167
rect 213665 -10506 213700 -10167
rect 213799 -10448 214533 -10036
rect 214552 -10118 214921 -10084
rect 214652 -10256 214821 -10222
rect 214590 -10448 214625 -10306
rect 214848 -10448 214883 -10306
rect 214981 -10448 215029 -10083
rect 215035 -10448 215083 -10137
rect 215143 -10183 215512 -10149
rect 215243 -10321 215412 -10287
rect 213799 -10506 215154 -10448
rect 213226 -10543 215154 -10506
rect 215181 -10543 215216 -10371
rect 215439 -10543 215474 -10371
rect 215573 -10543 215608 -10245
rect 2525 -10667 4984 -10543
rect 5888 -10667 8328 -10543
rect 9233 -10667 11672 -10543
rect 12577 -10667 15016 -10543
rect 15922 -10667 18360 -10543
rect 19266 -10667 21704 -10543
rect 22610 -10667 25048 -10543
rect 25954 -10667 28392 -10543
rect 29299 -10667 31736 -10543
rect 32643 -10667 35080 -10543
rect 35987 -10667 38424 -10543
rect 39331 -10667 41768 -10543
rect 42675 -10667 45112 -10543
rect 46019 -10667 48456 -10543
rect 49363 -10667 51800 -10543
rect 52707 -10667 55144 -10543
rect 56052 -10667 58488 -10543
rect 59396 -10667 61832 -10543
rect 62740 -10667 65176 -10543
rect 66084 -10667 68520 -10543
rect 69428 -10667 71864 -10543
rect 72772 -10667 75208 -10543
rect 76116 -10667 78552 -10543
rect 79460 -10667 81896 -10543
rect 82804 -10667 85240 -10543
rect 86148 -10667 88584 -10543
rect 89492 -10667 91928 -10543
rect 92836 -10667 95272 -10543
rect 96180 -10667 98616 -10543
rect 99524 -10667 101960 -10543
rect 102868 -10667 105304 -10543
rect 106212 -10667 108648 -10543
rect 109562 -10667 111992 -10543
rect 112906 -10667 115336 -10543
rect 116250 -10667 118680 -10543
rect 119594 -10667 122024 -10543
rect 122938 -10667 125368 -10543
rect 126282 -10667 128712 -10543
rect 129626 -10667 132056 -10543
rect 132970 -10667 135400 -10543
rect 136314 -10667 138744 -10543
rect 139658 -10667 142088 -10543
rect 143002 -10667 145432 -10543
rect 146346 -10667 148776 -10543
rect 149690 -10667 152120 -10543
rect 153034 -10667 155464 -10543
rect 156378 -10667 158808 -10543
rect 159722 -10667 162152 -10543
rect 163066 -10667 165496 -10543
rect 166410 -10667 168840 -10543
rect 169754 -10667 172184 -10543
rect 173098 -10667 175528 -10543
rect 176442 -10667 178872 -10543
rect 179786 -10667 182216 -10543
rect 183130 -10667 185560 -10543
rect 186474 -10667 188904 -10543
rect 189818 -10667 192248 -10543
rect 193162 -10667 195592 -10543
rect 196506 -10667 198936 -10543
rect 199850 -10667 202280 -10543
rect 203194 -10667 205624 -10543
rect 206538 -10667 208968 -10543
rect 209882 -10667 212312 -10543
rect 213226 -10667 215656 -10543
rect 2525 -10764 5037 -10667
rect 2477 -10867 5037 -10764
rect 2477 -11763 5025 -10867
rect 5888 -11622 8381 -10667
rect 9233 -11622 11725 -10667
rect 12577 -11622 15069 -10667
rect 15922 -11622 18413 -10667
rect 19266 -11622 21757 -10667
rect 22610 -11622 25101 -10667
rect 25954 -11622 28445 -10667
rect 29299 -11622 31789 -10667
rect 32643 -11622 35133 -10667
rect 35987 -11622 38477 -10667
rect 39331 -11622 41821 -10667
rect 42675 -11622 45165 -10667
rect 46019 -11622 48509 -10667
rect 49363 -11622 51853 -10667
rect 52707 -11622 55197 -10667
rect 56052 -11622 58541 -10667
rect 59396 -11622 61885 -10667
rect 62740 -11622 65229 -10667
rect 66084 -11622 68573 -10667
rect 69428 -11622 71917 -10667
rect 72772 -11622 75261 -10667
rect 76116 -11622 78605 -10667
rect 79460 -11622 81949 -10667
rect 82804 -11622 85293 -10667
rect 86148 -11622 88637 -10667
rect 89492 -11622 91981 -10667
rect 92836 -11622 95325 -10667
rect 96180 -11622 98669 -10667
rect 99524 -11622 102013 -10667
rect 102868 -11622 105357 -10667
rect 106212 -11622 108701 -10667
rect 109562 -11622 112045 -10667
rect 112906 -11622 115389 -10667
rect 116250 -11622 118733 -10667
rect 119594 -11622 122077 -10667
rect 122938 -11622 125421 -10667
rect 126282 -11622 128765 -10667
rect 129626 -11622 132109 -10667
rect 132970 -11622 135453 -10667
rect 136314 -11622 138797 -10667
rect 139658 -11622 142141 -10667
rect 143002 -11622 145485 -10667
rect 146346 -11622 148829 -10667
rect 149690 -11622 152173 -10667
rect 153034 -11622 155517 -10667
rect 156378 -11622 158861 -10667
rect 159722 -11622 162205 -10667
rect 163066 -11622 165549 -10667
rect 166410 -11622 168893 -10667
rect 169754 -11622 172237 -10667
rect 173098 -11622 175581 -10667
rect 176442 -11622 178925 -10667
rect 179786 -11622 182269 -10667
rect 183130 -11622 185613 -10667
rect 186474 -11622 188957 -10667
rect 189818 -11622 192301 -10667
rect 193162 -11622 195645 -10667
rect 196506 -11622 198989 -10667
rect 199850 -11622 202333 -10667
rect 203194 -11622 205677 -10667
rect 206538 -11622 209021 -10667
rect 209882 -11622 212365 -10667
rect 213226 -11622 215709 -10667
rect 216571 -11622 217034 -10506
rect 6479 -11687 8381 -11622
rect 9824 -11687 11725 -11622
rect 13168 -11687 15069 -11622
rect 16513 -11687 18413 -11622
rect 19857 -11687 21757 -11622
rect 23201 -11687 25101 -11622
rect 26545 -11687 28445 -11622
rect 29890 -11687 31789 -11622
rect 33234 -11687 35133 -11622
rect 36578 -11687 38477 -11622
rect 39922 -11687 41821 -11622
rect 43266 -11687 45165 -11622
rect 46610 -11687 48509 -11622
rect 49954 -11687 51853 -11622
rect 53298 -11687 55197 -11622
rect 56643 -11687 58541 -11622
rect 59987 -11687 61885 -11622
rect 63331 -11687 65229 -11622
rect 66675 -11687 68573 -11622
rect 70019 -11687 71917 -11622
rect 73363 -11687 75261 -11622
rect 76707 -11687 78605 -11622
rect 80051 -11687 81949 -11622
rect 83395 -11687 85293 -11622
rect 86739 -11687 88637 -11622
rect 90083 -11687 91981 -11622
rect 93427 -11687 95325 -11622
rect 96771 -11687 98669 -11622
rect 100115 -11687 102013 -11622
rect 103459 -11687 105357 -11622
rect 106803 -11687 108701 -11622
rect 110153 -11687 112045 -11622
rect 113497 -11687 115389 -11622
rect 116841 -11687 118733 -11622
rect 120185 -11687 122077 -11622
rect 123529 -11687 125421 -11622
rect 126873 -11687 128765 -11622
rect 130217 -11687 132109 -11622
rect 133561 -11687 135453 -11622
rect 136905 -11687 138797 -11622
rect 140249 -11687 142141 -11622
rect 143593 -11687 145485 -11622
rect 146937 -11687 148829 -11622
rect 150281 -11687 152173 -11622
rect 153625 -11687 155517 -11622
rect 156969 -11687 158861 -11622
rect 160313 -11687 162205 -11622
rect 163657 -11687 165549 -11622
rect 167001 -11687 168893 -11622
rect 170345 -11687 172237 -11622
rect 173689 -11687 175581 -11622
rect 177033 -11687 178925 -11622
rect 180377 -11687 182269 -11622
rect 183721 -11687 185613 -11622
rect 187065 -11687 188957 -11622
rect 190409 -11687 192301 -11622
rect 193753 -11687 195645 -11622
rect 197097 -11687 198989 -11622
rect 200441 -11687 202333 -11622
rect 203785 -11687 205677 -11622
rect 207129 -11687 209021 -11622
rect 210473 -11687 212365 -11622
rect 213817 -11687 215709 -11622
rect 7070 -11747 8381 -11687
rect 10415 -11747 11725 -11687
rect 13759 -11747 15069 -11687
rect 17104 -11747 18413 -11687
rect 20448 -11747 21757 -11687
rect 23792 -11747 25101 -11687
rect 27136 -11747 28445 -11687
rect 30481 -11747 31789 -11687
rect 33825 -11747 35133 -11687
rect 37169 -11747 38477 -11687
rect 40513 -11747 41821 -11687
rect 43857 -11747 45165 -11687
rect 47201 -11747 48509 -11687
rect 50545 -11747 51853 -11687
rect 53889 -11747 55197 -11687
rect 57234 -11747 58541 -11687
rect 60578 -11747 61885 -11687
rect 63922 -11747 65229 -11687
rect 67266 -11747 68573 -11687
rect 70610 -11747 71917 -11687
rect 73954 -11747 75261 -11687
rect 77298 -11747 78605 -11687
rect 80642 -11747 81949 -11687
rect 83986 -11747 85293 -11687
rect 87330 -11747 88637 -11687
rect 90674 -11747 91981 -11687
rect 94018 -11747 95325 -11687
rect 97362 -11747 98669 -11687
rect 100706 -11747 102013 -11687
rect 104050 -11747 105357 -11687
rect 107394 -11747 108701 -11687
rect 110744 -11747 112045 -11687
rect 114088 -11747 115389 -11687
rect 117432 -11747 118733 -11687
rect 120776 -11747 122077 -11687
rect 124120 -11747 125421 -11687
rect 127464 -11747 128765 -11687
rect 130808 -11747 132109 -11687
rect 134152 -11747 135453 -11687
rect 137496 -11747 138797 -11687
rect 140840 -11747 142141 -11687
rect 144184 -11747 145485 -11687
rect 147528 -11747 148829 -11687
rect 150872 -11747 152173 -11687
rect 154216 -11747 155517 -11687
rect 157560 -11747 158861 -11687
rect 160904 -11747 162205 -11687
rect 164248 -11747 165549 -11687
rect 167592 -11747 168893 -11687
rect 170936 -11747 172237 -11687
rect 174280 -11747 175581 -11687
rect 177624 -11747 178925 -11687
rect 180968 -11747 182269 -11687
rect 184312 -11747 185613 -11687
rect 187656 -11747 188957 -11687
rect 191000 -11747 192301 -11687
rect 194344 -11747 195645 -11687
rect 197688 -11747 198989 -11687
rect 201032 -11747 202333 -11687
rect 204376 -11747 205677 -11687
rect 207720 -11747 209021 -11687
rect 211064 -11747 212365 -11687
rect 214408 -11747 215709 -11687
rect 7099 -11752 8381 -11747
rect 10444 -11752 11725 -11747
rect 13788 -11752 15069 -11747
rect 17133 -11752 18413 -11747
rect 20477 -11752 21757 -11747
rect 23821 -11752 25101 -11747
rect 27165 -11752 28445 -11747
rect 30510 -11752 31789 -11747
rect 33854 -11752 35133 -11747
rect 37198 -11752 38477 -11747
rect 40542 -11752 41821 -11747
rect 43886 -11752 45165 -11747
rect 47230 -11752 48509 -11747
rect 50574 -11752 51853 -11747
rect 53918 -11752 55197 -11747
rect 57263 -11752 58541 -11747
rect 60607 -11752 61885 -11747
rect 63951 -11752 65229 -11747
rect 67295 -11752 68573 -11747
rect 70639 -11752 71917 -11747
rect 73983 -11752 75261 -11747
rect 77327 -11752 78605 -11747
rect 80671 -11752 81949 -11747
rect 84015 -11752 85293 -11747
rect 87359 -11752 88637 -11747
rect 90703 -11752 91981 -11747
rect 94047 -11752 95325 -11747
rect 97391 -11752 98669 -11747
rect 100735 -11752 102013 -11747
rect 104079 -11752 105357 -11747
rect 107423 -11752 108701 -11747
rect 110773 -11752 112045 -11747
rect 114117 -11752 115389 -11747
rect 117461 -11752 118733 -11747
rect 120805 -11752 122077 -11747
rect 124149 -11752 125421 -11747
rect 127493 -11752 128765 -11747
rect 130837 -11752 132109 -11747
rect 134181 -11752 135453 -11747
rect 137525 -11752 138797 -11747
rect 140869 -11752 142141 -11747
rect 144213 -11752 145485 -11747
rect 147557 -11752 148829 -11747
rect 150901 -11752 152173 -11747
rect 154245 -11752 155517 -11747
rect 157589 -11752 158861 -11747
rect 160933 -11752 162205 -11747
rect 164277 -11752 165549 -11747
rect 167621 -11752 168893 -11747
rect 170965 -11752 172237 -11747
rect 174309 -11752 175581 -11747
rect 177653 -11752 178925 -11747
rect 180997 -11752 182269 -11747
rect 184341 -11752 185613 -11747
rect 187685 -11752 188957 -11747
rect 191029 -11752 192301 -11747
rect 194373 -11752 195645 -11747
rect 197717 -11752 198989 -11747
rect 201061 -11752 202333 -11747
rect 204405 -11752 205677 -11747
rect 207749 -11752 209021 -11747
rect 211093 -11752 212365 -11747
rect 214437 -11752 215709 -11747
rect 2477 -11781 5013 -11763
rect 7234 -11770 8381 -11752
rect 10578 -11770 11725 -11752
rect 13922 -11770 15069 -11752
rect 17266 -11770 18413 -11752
rect 20610 -11770 21757 -11752
rect 23954 -11770 25101 -11752
rect 27298 -11770 28445 -11752
rect 30642 -11770 31789 -11752
rect 33986 -11770 35133 -11752
rect 37330 -11770 38477 -11752
rect 40674 -11770 41821 -11752
rect 44018 -11770 45165 -11752
rect 47362 -11770 48509 -11752
rect 50706 -11770 51853 -11752
rect 54050 -11770 55197 -11752
rect 57394 -11770 58541 -11752
rect 60738 -11770 61885 -11752
rect 64082 -11770 65229 -11752
rect 67426 -11770 68573 -11752
rect 70770 -11770 71917 -11752
rect 74114 -11770 75261 -11752
rect 77458 -11770 78605 -11752
rect 80802 -11770 81949 -11752
rect 84146 -11770 85293 -11752
rect 87490 -11770 88637 -11752
rect 90834 -11770 91981 -11752
rect 94178 -11770 95325 -11752
rect 97522 -11770 98669 -11752
rect 100866 -11770 102013 -11752
rect 104210 -11770 105357 -11752
rect 107554 -11770 108701 -11752
rect 110898 -11770 112045 -11752
rect 114242 -11770 115389 -11752
rect 117586 -11770 118733 -11752
rect 120930 -11770 122077 -11752
rect 124274 -11770 125421 -11752
rect 127618 -11770 128765 -11752
rect 130962 -11770 132109 -11752
rect 134306 -11770 135453 -11752
rect 137650 -11770 138797 -11752
rect 140994 -11770 142141 -11752
rect 144338 -11770 145485 -11752
rect 147682 -11770 148829 -11752
rect 151026 -11770 152173 -11752
rect 154370 -11770 155517 -11752
rect 157714 -11770 158861 -11752
rect 161058 -11770 162205 -11752
rect 164402 -11770 165549 -11752
rect 167746 -11770 168893 -11752
rect 171090 -11770 172237 -11752
rect 174434 -11770 175581 -11752
rect 177778 -11770 178925 -11752
rect 181122 -11770 182269 -11752
rect 184466 -11770 185613 -11752
rect 187810 -11770 188957 -11752
rect 191154 -11770 192301 -11752
rect 194498 -11770 195645 -11752
rect 197842 -11770 198989 -11752
rect 201186 -11770 202333 -11752
rect 204530 -11770 205677 -11752
rect 207874 -11770 209021 -11752
rect 211218 -11770 212365 -11752
rect 214562 -11770 215709 -11752
rect 7661 -11781 8381 -11770
rect 11006 -11781 11725 -11770
rect 14350 -11781 15069 -11770
rect 17695 -11781 18413 -11770
rect 21039 -11781 21757 -11770
rect 24383 -11781 25101 -11770
rect 27727 -11781 28445 -11770
rect 31072 -11781 31789 -11770
rect 34416 -11781 35133 -11770
rect 37760 -11781 38477 -11770
rect 41104 -11781 41821 -11770
rect 44448 -11781 45165 -11770
rect 47792 -11781 48509 -11770
rect 51136 -11781 51853 -11770
rect 54480 -11781 55197 -11770
rect 57825 -11781 58541 -11770
rect 61169 -11781 61885 -11770
rect 64513 -11781 65229 -11770
rect 67857 -11781 68573 -11770
rect 71201 -11781 71917 -11770
rect 74545 -11781 75261 -11770
rect 77889 -11781 78605 -11770
rect 81233 -11781 81949 -11770
rect 84577 -11781 85293 -11770
rect 87921 -11781 88637 -11770
rect 91265 -11781 91981 -11770
rect 94609 -11781 95325 -11770
rect 97953 -11781 98669 -11770
rect 101297 -11781 102013 -11770
rect 104641 -11781 105357 -11770
rect 107985 -11781 108701 -11770
rect 111335 -11781 112045 -11770
rect 114679 -11781 115389 -11770
rect 118023 -11781 118733 -11770
rect 121367 -11781 122077 -11770
rect 124711 -11781 125421 -11770
rect 128055 -11781 128765 -11770
rect 131399 -11781 132109 -11770
rect 134743 -11781 135453 -11770
rect 138087 -11781 138797 -11770
rect 141431 -11781 142141 -11770
rect 144775 -11781 145485 -11770
rect 148119 -11781 148829 -11770
rect 151463 -11781 152173 -11770
rect 154807 -11781 155517 -11770
rect 158151 -11781 158861 -11770
rect 161495 -11781 162205 -11770
rect 164839 -11781 165549 -11770
rect 168183 -11781 168893 -11770
rect 171527 -11781 172237 -11770
rect 174871 -11781 175581 -11770
rect 178215 -11781 178925 -11770
rect 181559 -11781 182269 -11770
rect 184903 -11781 185613 -11770
rect 188247 -11781 188957 -11770
rect 191591 -11781 192301 -11770
rect 194935 -11781 195645 -11770
rect 198279 -11781 198989 -11770
rect 201623 -11781 202333 -11770
rect 204967 -11781 205677 -11770
rect 208311 -11781 209021 -11770
rect 211655 -11781 212365 -11770
rect 214999 -11781 215709 -11770
rect 2477 -11813 5022 -11781
rect 2477 -11817 4984 -11813
rect 7661 -11817 8346 -11781
rect 11006 -11817 11690 -11781
rect 14350 -11817 15034 -11781
rect 17695 -11817 18378 -11781
rect 21039 -11817 21722 -11781
rect 24383 -11817 25066 -11781
rect 27727 -11817 28410 -11781
rect 31072 -11817 31754 -11781
rect 34416 -11817 35098 -11781
rect 37760 -11817 38442 -11781
rect 41104 -11817 41786 -11781
rect 44448 -11817 45130 -11781
rect 47792 -11817 48474 -11781
rect 51136 -11817 51818 -11781
rect 54480 -11817 55162 -11781
rect 57825 -11817 58506 -11781
rect 61169 -11817 61850 -11781
rect 64513 -11817 65194 -11781
rect 67857 -11817 68538 -11781
rect 71201 -11817 71882 -11781
rect 74545 -11817 75226 -11781
rect 77889 -11817 78570 -11781
rect 81233 -11817 81914 -11781
rect 84577 -11817 85258 -11781
rect 87921 -11817 88602 -11781
rect 91265 -11817 91946 -11781
rect 94609 -11817 95290 -11781
rect 97953 -11817 98634 -11781
rect 101297 -11817 101978 -11781
rect 104641 -11817 105322 -11781
rect 107985 -11817 108666 -11781
rect 111335 -11817 112010 -11781
rect 114679 -11817 115354 -11781
rect 118023 -11817 118698 -11781
rect 121367 -11817 122042 -11781
rect 124711 -11817 125386 -11781
rect 128055 -11817 128730 -11781
rect 131399 -11817 132074 -11781
rect 134743 -11817 135418 -11781
rect 138087 -11817 138762 -11781
rect 141431 -11817 142106 -11781
rect 144775 -11817 145450 -11781
rect 148119 -11817 148794 -11781
rect 151463 -11817 152138 -11781
rect 154807 -11817 155482 -11781
rect 158151 -11817 158826 -11781
rect 161495 -11817 162170 -11781
rect 164839 -11817 165514 -11781
rect 168183 -11817 168858 -11781
rect 171527 -11817 172202 -11781
rect 174871 -11817 175546 -11781
rect 178215 -11817 178890 -11781
rect 181559 -11817 182234 -11781
rect 184903 -11817 185578 -11781
rect 188247 -11817 188922 -11781
rect 191591 -11817 192266 -11781
rect 194935 -11817 195610 -11781
rect 198279 -11817 198954 -11781
rect 201623 -11817 202298 -11781
rect 204967 -11817 205642 -11781
rect 208311 -11817 208986 -11781
rect 211655 -11817 212330 -11781
rect 214999 -11817 215674 -11781
rect 2477 -11825 4906 -11817
rect 4913 -11825 4947 -11817
rect 4980 -11825 4981 -11817
rect 2477 -11859 4947 -11825
rect 7855 -11835 8346 -11817
rect 11199 -11835 11690 -11817
rect 14543 -11835 15034 -11817
rect 17887 -11835 18378 -11817
rect 21231 -11835 21722 -11817
rect 24575 -11835 25066 -11817
rect 27919 -11835 28410 -11817
rect 31263 -11835 31754 -11817
rect 34607 -11835 35098 -11817
rect 37951 -11835 38442 -11817
rect 41295 -11835 41786 -11817
rect 44639 -11835 45130 -11817
rect 47983 -11835 48474 -11817
rect 51327 -11835 51818 -11817
rect 54671 -11835 55162 -11817
rect 58015 -11835 58506 -11817
rect 61359 -11835 61850 -11817
rect 64703 -11835 65194 -11817
rect 68047 -11835 68538 -11817
rect 71391 -11835 71882 -11817
rect 74735 -11835 75226 -11817
rect 78079 -11835 78570 -11817
rect 81423 -11835 81914 -11817
rect 84767 -11835 85258 -11817
rect 88111 -11835 88602 -11817
rect 91455 -11835 91946 -11817
rect 94799 -11835 95290 -11817
rect 98143 -11835 98634 -11817
rect 101487 -11835 101978 -11817
rect 104831 -11835 105322 -11817
rect 108175 -11835 108666 -11817
rect 111519 -11835 112010 -11817
rect 114863 -11835 115354 -11817
rect 118207 -11835 118698 -11817
rect 121551 -11835 122042 -11817
rect 124895 -11835 125386 -11817
rect 128239 -11835 128730 -11817
rect 131583 -11835 132074 -11817
rect 134927 -11835 135418 -11817
rect 138271 -11835 138762 -11817
rect 141615 -11835 142106 -11817
rect 144959 -11835 145450 -11817
rect 148303 -11835 148794 -11817
rect 151647 -11835 152138 -11817
rect 154991 -11835 155482 -11817
rect 158335 -11835 158826 -11817
rect 161679 -11835 162170 -11817
rect 165023 -11835 165514 -11817
rect 168367 -11835 168858 -11817
rect 171711 -11835 172202 -11817
rect 175055 -11835 175546 -11817
rect 178399 -11835 178890 -11817
rect 181743 -11835 182234 -11817
rect 185087 -11835 185578 -11817
rect 188431 -11835 188922 -11817
rect 191775 -11835 192266 -11817
rect 195119 -11835 195610 -11817
rect 198463 -11835 198954 -11817
rect 201807 -11835 202298 -11817
rect 205151 -11835 205642 -11817
rect 208495 -11835 208986 -11817
rect 211839 -11835 212330 -11817
rect 215183 -11835 215674 -11817
rect 7894 -11859 8273 -11835
rect 11239 -11859 11617 -11835
rect 14583 -11859 14961 -11835
rect 17928 -11859 18305 -11835
rect 21272 -11859 21649 -11835
rect 24616 -11859 24993 -11835
rect 27960 -11859 28337 -11835
rect 31305 -11859 31681 -11835
rect 34649 -11859 35025 -11835
rect 37993 -11859 38369 -11835
rect 41337 -11859 41713 -11835
rect 44681 -11859 45057 -11835
rect 48025 -11859 48401 -11835
rect 51369 -11859 51745 -11835
rect 54713 -11859 55089 -11835
rect 58058 -11859 58433 -11835
rect 61402 -11859 61777 -11835
rect 64746 -11859 65121 -11835
rect 68090 -11859 68465 -11835
rect 71434 -11859 71809 -11835
rect 74778 -11859 75153 -11835
rect 78122 -11859 78497 -11835
rect 81466 -11859 81841 -11835
rect 84810 -11859 85185 -11835
rect 88154 -11859 88529 -11835
rect 91498 -11859 91873 -11835
rect 94842 -11859 95217 -11835
rect 98186 -11859 98561 -11835
rect 101530 -11859 101905 -11835
rect 104874 -11859 105249 -11835
rect 108218 -11859 108593 -11835
rect 111568 -11859 111937 -11835
rect 114912 -11859 115281 -11835
rect 118256 -11859 118625 -11835
rect 121600 -11859 121969 -11835
rect 124944 -11859 125313 -11835
rect 128288 -11859 128657 -11835
rect 131632 -11859 132001 -11835
rect 134976 -11859 135345 -11835
rect 138320 -11859 138689 -11835
rect 141664 -11859 142033 -11835
rect 145008 -11859 145377 -11835
rect 148352 -11859 148721 -11835
rect 151696 -11859 152065 -11835
rect 155040 -11859 155409 -11835
rect 158384 -11859 158753 -11835
rect 161728 -11859 162097 -11835
rect 165072 -11859 165441 -11835
rect 168416 -11859 168785 -11835
rect 171760 -11859 172129 -11835
rect 175104 -11859 175473 -11835
rect 178448 -11859 178817 -11835
rect 181792 -11859 182161 -11835
rect 185136 -11859 185505 -11835
rect 188480 -11859 188849 -11835
rect 191824 -11859 192193 -11835
rect 195168 -11859 195537 -11835
rect 198512 -11859 198881 -11835
rect 201856 -11859 202225 -11835
rect 205200 -11859 205569 -11835
rect 208544 -11859 208913 -11835
rect 211888 -11859 212257 -11835
rect 215232 -11859 215601 -11835
rect 2477 -11871 4906 -11859
rect 4913 -11871 4947 -11859
rect 2477 -11880 4959 -11871
rect 3068 -11945 4959 -11880
rect 3659 -12005 4959 -11945
rect 3688 -12010 4959 -12005
rect 3812 -12028 4959 -12010
rect 4250 -12039 4959 -12028
rect 4250 -12075 4924 -12039
rect 4433 -12093 4924 -12075
<< error_ps >>
rect 217161 -9114 217305 -8874
rect 217491 -8899 217877 -8753
rect 217415 -8985 217877 -8899
rect 217161 -9200 217335 -9114
rect 217162 -10036 217818 -9971
rect 217162 -10448 217877 -10036
rect 217162 -10506 218294 -10448
rect 217034 -11622 218294 -10506
rect 217162 -11687 218294 -11622
rect 217753 -11747 218294 -11687
rect 217782 -11752 218294 -11747
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
use icell1scs  x1
timestamp 1717439242
transform 1 0 3 0 1 -5600
box -66 -6595 5022 200
use icell2scs  x2
timestamp 1717439242
transform 1 0 4 0 1 -5600
box 0 -6337 8432 458
use icell4scs  x3
timestamp 1717439242
transform 1 0 5 0 1 -5600
box 0 -6337 15120 458
use mosgsconnected  x4
timestamp 1717439242
transform 1 0 16 0 1 -5600
box -95 -495 621 2499
use p_ibias_mirror  x5
timestamp 1717439242
transform 1 0 17 0 1 -5600
box -95 -2270 7078 1109
use lvhvbuff  x6
timestamp 1717439242
transform 1 0 0 0 1 -5600
box -66 -1729 4518 200
use lvhvbuff  x7
timestamp 1717439242
transform 1 0 1 0 1 -5600
box -66 -1729 4518 200
use lvhvbuff  x8
timestamp 1717439242
transform 1 0 2 0 1 -5600
box -66 -1729 4518 200
use icell8scs  x9
timestamp 1717439242
transform 1 0 6 0 1 -5600
box 0 -6337 28496 458
use icell16scs  x10
timestamp 1717439242
transform 1 0 7 0 1 -5600
box 0 -6337 55248 458
use icell32scs  x11
timestamp 1717439242
transform 1 0 8 0 1 -5600
box 0 -6337 108752 458
use lvhvbuff  x12
timestamp 1717439242
transform 1 0 9 0 1 -5600
box -66 -1729 4518 200
use lvhvbuff  x13
timestamp 1717439242
transform 1 0 10 0 1 -5600
box -66 -1729 4518 200
use lvhvbuff  x14
timestamp 1717439242
transform 1 0 11 0 1 -5600
box -66 -1729 4518 200
use lvhvbuff  x15
timestamp 1717439242
transform 1 0 12 0 1 -5600
box -66 -1729 4518 200
use lvhvbuff  x16
timestamp 1717439242
transform 1 0 13 0 1 -5600
box -66 -1729 4518 200
use icell64scs  x17
timestamp 1717439242
transform 1 0 14 0 1 -5600
box 0 -6337 215760 458
use icell128scs  x18
timestamp 1717439242
transform 1 0 15 0 1 -5600
box 0 -6337 429776 458
use n_ibias_mirror  x19
timestamp 1717439242
transform 1 0 18 0 1 -5600
box -65 -1985 4815 721
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 avdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 dvdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 iout
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 din0
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 idir_sel
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 din1
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 avss
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 din2
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 din3
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 iref
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 din4
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 din5
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 din6
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 din7
port 14 nsew
<< end >>
