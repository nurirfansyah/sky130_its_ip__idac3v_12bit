magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 3986 655814 4368 655848
rect 3890 348809 3938 655752
rect 4086 655676 4268 655710
rect 4070 655617 4072 655628
rect 4271 655617 4284 655628
rect 4024 653241 4072 655617
rect 4282 653241 4330 655617
rect 4086 653148 4268 653182
rect 4086 653040 4268 653074
rect 4070 652981 4072 652992
rect 4271 652981 4284 652992
rect 4024 650605 4072 652981
rect 4282 650605 4330 652981
rect 4086 650512 4268 650546
rect 4086 650404 4268 650438
rect 4070 650345 4072 650356
rect 4271 650345 4284 650356
rect 4024 647969 4072 650345
rect 4282 647969 4330 650345
rect 4086 647876 4268 647910
rect 4086 647768 4268 647802
rect 4070 647709 4072 647720
rect 4271 647709 4284 647720
rect 4024 645333 4072 647709
rect 4282 645333 4330 647709
rect 4086 645240 4268 645274
rect 4086 645132 4268 645166
rect 4070 645073 4072 645084
rect 4271 645073 4284 645084
rect 4024 642697 4072 645073
rect 4282 642697 4330 645073
rect 4086 642604 4268 642638
rect 4086 642496 4268 642530
rect 4070 642437 4072 642448
rect 4271 642437 4284 642448
rect 4024 640061 4072 642437
rect 4282 640061 4330 642437
rect 4086 639968 4268 640002
rect 4086 639860 4268 639894
rect 4070 639801 4072 639812
rect 4271 639801 4284 639812
rect 4024 637425 4072 639801
rect 4282 637425 4330 639801
rect 4086 637332 4268 637366
rect 4086 637224 4268 637258
rect 4070 637165 4072 637176
rect 4271 637165 4284 637176
rect 4024 634789 4072 637165
rect 4282 634789 4330 637165
rect 4086 634696 4268 634730
rect 4086 634588 4268 634622
rect 4070 634529 4072 634540
rect 4271 634529 4284 634540
rect 4024 632153 4072 634529
rect 4282 632153 4330 634529
rect 4086 632060 4268 632094
rect 4086 631952 4268 631986
rect 4070 631893 4072 631904
rect 4271 631893 4284 631904
rect 4024 629517 4072 631893
rect 4282 629517 4330 631893
rect 4086 629424 4268 629458
rect 4086 629316 4268 629350
rect 4070 629257 4072 629268
rect 4271 629257 4284 629268
rect 4024 626881 4072 629257
rect 4282 626881 4330 629257
rect 4086 626788 4268 626822
rect 4086 626680 4268 626714
rect 4070 626621 4072 626632
rect 4271 626621 4284 626632
rect 4024 624245 4072 626621
rect 4282 624245 4330 626621
rect 4086 624152 4268 624186
rect 4086 624044 4268 624078
rect 4070 623985 4072 623996
rect 4271 623985 4284 623996
rect 4024 621609 4072 623985
rect 4282 621609 4330 623985
rect 4086 621516 4268 621550
rect 4086 621408 4268 621442
rect 4070 621349 4072 621360
rect 4271 621349 4284 621360
rect 4024 618973 4072 621349
rect 4282 618973 4330 621349
rect 4086 618880 4268 618914
rect 4086 618772 4268 618806
rect 4070 618713 4072 618724
rect 4271 618713 4284 618724
rect 4024 616337 4072 618713
rect 4282 616337 4330 618713
rect 4086 616244 4268 616278
rect 4086 616136 4268 616170
rect 4070 616077 4072 616088
rect 4271 616077 4284 616088
rect 4024 613701 4072 616077
rect 4282 613701 4330 616077
rect 4086 613608 4268 613642
rect 4086 613500 4268 613534
rect 4070 613441 4072 613452
rect 4271 613441 4284 613452
rect 4024 611065 4072 613441
rect 4282 611065 4330 613441
rect 4086 610972 4268 611006
rect 4086 610864 4268 610898
rect 4070 610805 4072 610816
rect 4271 610805 4284 610816
rect 4024 608429 4072 610805
rect 4282 608429 4330 610805
rect 4086 608336 4268 608370
rect 4086 608228 4268 608262
rect 4070 608169 4072 608180
rect 4271 608169 4284 608180
rect 4024 605793 4072 608169
rect 4282 605793 4330 608169
rect 4086 605700 4268 605734
rect 4086 605592 4268 605626
rect 4070 605533 4072 605544
rect 4271 605533 4284 605544
rect 4024 603157 4072 605533
rect 4282 603157 4330 605533
rect 4086 603064 4268 603098
rect 4086 602956 4268 602990
rect 4070 602897 4072 602908
rect 4271 602897 4284 602908
rect 4024 600521 4072 602897
rect 4282 600521 4330 602897
rect 4086 600428 4268 600462
rect 4086 600320 4268 600354
rect 4070 600261 4072 600272
rect 4271 600261 4284 600272
rect 4024 597885 4072 600261
rect 4282 597885 4330 600261
rect 4086 597792 4268 597826
rect 4086 597684 4268 597718
rect 4070 597625 4072 597636
rect 4271 597625 4284 597636
rect 4024 595249 4072 597625
rect 4282 595249 4330 597625
rect 4086 595156 4268 595190
rect 4086 595048 4268 595082
rect 4070 594989 4072 595000
rect 4271 594989 4284 595000
rect 4024 592613 4072 594989
rect 4282 592613 4330 594989
rect 4086 592520 4268 592554
rect 4086 592412 4268 592446
rect 4070 592353 4072 592364
rect 4271 592353 4284 592364
rect 4024 589977 4072 592353
rect 4282 589977 4330 592353
rect 4086 589884 4268 589918
rect 4086 589776 4268 589810
rect 4070 589717 4072 589728
rect 4271 589717 4284 589728
rect 4024 587341 4072 589717
rect 4282 587341 4330 589717
rect 4086 587248 4268 587282
rect 4086 587140 4268 587174
rect 4070 587081 4072 587092
rect 4271 587081 4284 587092
rect 4024 584705 4072 587081
rect 4282 584705 4330 587081
rect 4086 584612 4268 584646
rect 4086 584504 4268 584538
rect 4070 584445 4072 584456
rect 4271 584445 4284 584456
rect 4024 582069 4072 584445
rect 4282 582069 4330 584445
rect 4086 581976 4268 582010
rect 4086 581868 4268 581902
rect 4070 581809 4072 581820
rect 4271 581809 4284 581820
rect 4024 579433 4072 581809
rect 4282 579433 4330 581809
rect 4086 579340 4268 579374
rect 4086 579232 4268 579266
rect 4070 579173 4072 579184
rect 4271 579173 4284 579184
rect 4024 576797 4072 579173
rect 4282 576797 4330 579173
rect 4086 576704 4268 576738
rect 4086 576596 4268 576630
rect 4070 576537 4072 576548
rect 4271 576537 4284 576548
rect 4024 574161 4072 576537
rect 4282 574161 4330 576537
rect 4086 574068 4268 574102
rect 4086 573960 4268 573994
rect 4070 573901 4072 573912
rect 4271 573901 4284 573912
rect 4024 571525 4072 573901
rect 4282 571525 4330 573901
rect 4086 571432 4268 571466
rect 4086 571324 4268 571358
rect 4070 571265 4072 571276
rect 4271 571265 4284 571276
rect 4024 568889 4072 571265
rect 4282 568889 4330 571265
rect 4086 568796 4268 568830
rect 4086 568688 4268 568722
rect 4070 568629 4072 568640
rect 4271 568629 4284 568640
rect 4024 566253 4072 568629
rect 4282 566253 4330 568629
rect 4086 566160 4268 566194
rect 4086 566052 4268 566086
rect 4070 565993 4072 566004
rect 4271 565993 4284 566004
rect 4024 563617 4072 565993
rect 4282 563617 4330 565993
rect 4086 563524 4268 563558
rect 4086 563416 4268 563450
rect 4070 563357 4072 563368
rect 4271 563357 4284 563368
rect 4024 560981 4072 563357
rect 4282 560981 4330 563357
rect 4086 560888 4268 560922
rect 4086 560780 4268 560814
rect 4070 560721 4072 560732
rect 4271 560721 4284 560732
rect 4024 558345 4072 560721
rect 4282 558345 4330 560721
rect 4086 558252 4268 558286
rect 4086 558144 4268 558178
rect 4070 558085 4072 558096
rect 4271 558085 4284 558096
rect 4024 555709 4072 558085
rect 4282 555709 4330 558085
rect 4086 555616 4268 555650
rect 4086 555508 4268 555542
rect 4070 555449 4072 555460
rect 4271 555449 4284 555460
rect 4024 553073 4072 555449
rect 4282 553073 4330 555449
rect 4086 552980 4268 553014
rect 4086 552872 4268 552906
rect 4070 552813 4072 552824
rect 4271 552813 4284 552824
rect 4024 550437 4072 552813
rect 4282 550437 4330 552813
rect 4086 550344 4268 550378
rect 4086 550236 4268 550270
rect 4070 550177 4072 550188
rect 4271 550177 4284 550188
rect 4024 547801 4072 550177
rect 4282 547801 4330 550177
rect 4086 547708 4268 547742
rect 4086 547600 4268 547634
rect 4070 547541 4072 547552
rect 4271 547541 4284 547552
rect 4024 545165 4072 547541
rect 4282 545165 4330 547541
rect 4086 545072 4268 545106
rect 4086 544964 4268 544998
rect 4070 544905 4072 544916
rect 4271 544905 4284 544916
rect 4024 542529 4072 544905
rect 4282 542529 4330 544905
rect 4086 542436 4268 542470
rect 4086 542328 4268 542362
rect 4070 542269 4072 542280
rect 4271 542269 4284 542280
rect 4024 539893 4072 542269
rect 4282 539893 4330 542269
rect 4086 539800 4268 539834
rect 4086 539692 4268 539726
rect 4070 539633 4072 539644
rect 4271 539633 4284 539644
rect 4024 537257 4072 539633
rect 4282 537257 4330 539633
rect 4086 537164 4268 537198
rect 4086 537056 4268 537090
rect 4070 536997 4072 537008
rect 4271 536997 4284 537008
rect 4024 534621 4072 536997
rect 4282 534621 4330 536997
rect 4086 534528 4268 534562
rect 4086 534420 4268 534454
rect 4070 534361 4072 534372
rect 4271 534361 4284 534372
rect 4024 531985 4072 534361
rect 4282 531985 4330 534361
rect 4086 531892 4268 531926
rect 4086 531784 4268 531818
rect 4070 531725 4072 531736
rect 4271 531725 4284 531736
rect 4024 529349 4072 531725
rect 4282 529349 4330 531725
rect 4086 529256 4268 529290
rect 4086 529148 4268 529182
rect 4070 529089 4072 529100
rect 4271 529089 4284 529100
rect 4024 526713 4072 529089
rect 4282 526713 4330 529089
rect 4086 526620 4268 526654
rect 4086 526512 4268 526546
rect 4070 526453 4072 526464
rect 4271 526453 4284 526464
rect 4024 524077 4072 526453
rect 4282 524077 4330 526453
rect 4086 523984 4268 524018
rect 4086 523876 4268 523910
rect 4070 523817 4072 523828
rect 4271 523817 4284 523828
rect 4024 521441 4072 523817
rect 4282 521441 4330 523817
rect 4086 521348 4268 521382
rect 4086 521240 4268 521274
rect 4070 521181 4072 521192
rect 4271 521181 4284 521192
rect 4024 518805 4072 521181
rect 4282 518805 4330 521181
rect 4086 518712 4268 518746
rect 4086 518604 4268 518638
rect 4070 518545 4072 518556
rect 4271 518545 4284 518556
rect 4024 516169 4072 518545
rect 4282 516169 4330 518545
rect 4086 516076 4268 516110
rect 4086 515968 4268 516002
rect 4070 515909 4072 515920
rect 4271 515909 4284 515920
rect 4024 513533 4072 515909
rect 4282 513533 4330 515909
rect 4086 513440 4268 513474
rect 4086 513332 4268 513366
rect 4070 513273 4072 513284
rect 4271 513273 4284 513284
rect 4024 510897 4072 513273
rect 4282 510897 4330 513273
rect 4086 510804 4268 510838
rect 4086 510696 4268 510730
rect 4070 510637 4072 510648
rect 4271 510637 4284 510648
rect 4024 508261 4072 510637
rect 4282 508261 4330 510637
rect 4086 508168 4268 508202
rect 4086 508060 4268 508094
rect 4070 508001 4072 508012
rect 4271 508001 4284 508012
rect 4024 505625 4072 508001
rect 4282 505625 4330 508001
rect 4086 505532 4268 505566
rect 4086 505424 4268 505458
rect 4070 505365 4072 505376
rect 4271 505365 4284 505376
rect 4024 502989 4072 505365
rect 4282 502989 4330 505365
rect 4086 502896 4268 502930
rect 4086 502788 4268 502822
rect 4070 502729 4072 502740
rect 4271 502729 4284 502740
rect 4024 500353 4072 502729
rect 4282 500353 4330 502729
rect 4086 500260 4268 500294
rect 4086 500152 4268 500186
rect 4070 500093 4072 500104
rect 4271 500093 4284 500104
rect 4024 497717 4072 500093
rect 4282 497717 4330 500093
rect 4086 497624 4268 497658
rect 4086 497516 4268 497550
rect 4070 497457 4072 497468
rect 4271 497457 4284 497468
rect 4024 495081 4072 497457
rect 4282 495081 4330 497457
rect 4086 494988 4268 495022
rect 4086 494880 4268 494914
rect 4070 494821 4072 494832
rect 4271 494821 4284 494832
rect 4024 492445 4072 494821
rect 4282 492445 4330 494821
rect 4086 492352 4268 492386
rect 4086 492244 4268 492278
rect 4070 492185 4072 492196
rect 4271 492185 4284 492196
rect 4024 489809 4072 492185
rect 4282 489809 4330 492185
rect 4086 489716 4268 489750
rect 4086 489608 4268 489642
rect 4070 489549 4072 489560
rect 4271 489549 4284 489560
rect 4024 487173 4072 489549
rect 4282 487173 4330 489549
rect 4086 487080 4268 487114
rect 4086 486972 4268 487006
rect 4070 486913 4072 486924
rect 4271 486913 4284 486924
rect 4024 484537 4072 486913
rect 4282 484537 4330 486913
rect 4086 484444 4268 484478
rect 4086 484336 4268 484370
rect 4070 484277 4072 484288
rect 4271 484277 4284 484288
rect 4024 481901 4072 484277
rect 4282 481901 4330 484277
rect 4086 481808 4268 481842
rect 4086 481700 4268 481734
rect 4070 481641 4072 481652
rect 4271 481641 4284 481652
rect 4024 479265 4072 481641
rect 4282 479265 4330 481641
rect 4086 479172 4268 479206
rect 4086 479064 4268 479098
rect 4070 479005 4072 479016
rect 4271 479005 4284 479016
rect 4024 476629 4072 479005
rect 4282 476629 4330 479005
rect 4086 476536 4268 476570
rect 4086 476428 4268 476462
rect 4070 476369 4072 476380
rect 4271 476369 4284 476380
rect 4024 473993 4072 476369
rect 4282 473993 4330 476369
rect 4086 473900 4268 473934
rect 4086 473792 4268 473826
rect 4070 473733 4072 473744
rect 4271 473733 4284 473744
rect 4024 471357 4072 473733
rect 4282 471357 4330 473733
rect 4086 471264 4268 471298
rect 4086 471156 4268 471190
rect 4070 471097 4072 471108
rect 4271 471097 4284 471108
rect 4024 468721 4072 471097
rect 4282 468721 4330 471097
rect 4086 468628 4268 468662
rect 4086 468520 4268 468554
rect 4070 468461 4072 468472
rect 4271 468461 4284 468472
rect 4024 466085 4072 468461
rect 4282 466085 4330 468461
rect 4086 465992 4268 466026
rect 4086 465884 4268 465918
rect 4070 465825 4072 465836
rect 4271 465825 4284 465836
rect 4024 463449 4072 465825
rect 4282 463449 4330 465825
rect 4086 463356 4268 463390
rect 4086 463248 4268 463282
rect 4070 463189 4072 463200
rect 4271 463189 4284 463200
rect 4024 460813 4072 463189
rect 4282 460813 4330 463189
rect 4086 460720 4268 460754
rect 4086 460612 4268 460646
rect 4070 460553 4072 460564
rect 4271 460553 4284 460564
rect 4024 458177 4072 460553
rect 4282 458177 4330 460553
rect 4086 458084 4268 458118
rect 4086 457976 4268 458010
rect 4070 457917 4072 457928
rect 4271 457917 4284 457928
rect 4024 455541 4072 457917
rect 4282 455541 4330 457917
rect 4086 455448 4268 455482
rect 4086 455340 4268 455374
rect 4070 455281 4072 455292
rect 4271 455281 4284 455292
rect 4024 452905 4072 455281
rect 4282 452905 4330 455281
rect 4086 452812 4268 452846
rect 4086 452704 4268 452738
rect 4070 452645 4072 452656
rect 4271 452645 4284 452656
rect 4024 450269 4072 452645
rect 4282 450269 4330 452645
rect 4086 450176 4268 450210
rect 4086 450068 4268 450102
rect 4070 450009 4072 450020
rect 4271 450009 4284 450020
rect 4024 447633 4072 450009
rect 4282 447633 4330 450009
rect 4086 447540 4268 447574
rect 4086 447432 4268 447466
rect 4070 447373 4072 447384
rect 4271 447373 4284 447384
rect 4024 444997 4072 447373
rect 4282 444997 4330 447373
rect 4086 444904 4268 444938
rect 4086 444796 4268 444830
rect 4070 444737 4072 444748
rect 4271 444737 4284 444748
rect 4024 442361 4072 444737
rect 4282 442361 4330 444737
rect 4086 442268 4268 442302
rect 4086 442160 4268 442194
rect 4070 442101 4072 442112
rect 4271 442101 4284 442112
rect 4024 439725 4072 442101
rect 4282 439725 4330 442101
rect 4086 439632 4268 439666
rect 4086 439524 4268 439558
rect 4070 439465 4072 439476
rect 4271 439465 4284 439476
rect 4024 437089 4072 439465
rect 4282 437089 4330 439465
rect 4086 436996 4268 437030
rect 4086 436888 4268 436922
rect 4070 436829 4072 436840
rect 4271 436829 4284 436840
rect 4024 434453 4072 436829
rect 4282 434453 4330 436829
rect 4086 434360 4268 434394
rect 4086 434252 4268 434286
rect 4070 434193 4072 434204
rect 4271 434193 4284 434204
rect 4024 431817 4072 434193
rect 4282 431817 4330 434193
rect 4086 431724 4268 431758
rect 4086 431616 4268 431650
rect 4070 431557 4072 431568
rect 4271 431557 4284 431568
rect 4024 429181 4072 431557
rect 4282 429181 4330 431557
rect 4086 429088 4268 429122
rect 4086 428980 4268 429014
rect 4070 428921 4072 428932
rect 4271 428921 4284 428932
rect 4024 426545 4072 428921
rect 4282 426545 4330 428921
rect 4086 426452 4268 426486
rect 4086 426344 4268 426378
rect 4070 426285 4072 426296
rect 4271 426285 4284 426296
rect 4024 423909 4072 426285
rect 4282 423909 4330 426285
rect 4086 423816 4268 423850
rect 4086 423708 4268 423742
rect 4070 423649 4072 423660
rect 4271 423649 4284 423660
rect 4024 421273 4072 423649
rect 4282 421273 4330 423649
rect 4086 421180 4268 421214
rect 4086 421072 4268 421106
rect 4070 421013 4072 421024
rect 4271 421013 4284 421024
rect 4024 418637 4072 421013
rect 4282 418637 4330 421013
rect 4086 418544 4268 418578
rect 4086 418436 4268 418470
rect 4070 418377 4072 418388
rect 4271 418377 4284 418388
rect 4024 416001 4072 418377
rect 4282 416001 4330 418377
rect 4086 415908 4268 415942
rect 4086 415800 4268 415834
rect 4070 415741 4072 415752
rect 4271 415741 4284 415752
rect 4024 413365 4072 415741
rect 4282 413365 4330 415741
rect 4086 413272 4268 413306
rect 4086 413164 4268 413198
rect 4070 413105 4072 413116
rect 4271 413105 4284 413116
rect 4024 410729 4072 413105
rect 4282 410729 4330 413105
rect 4086 410636 4268 410670
rect 4086 410528 4268 410562
rect 4070 410469 4072 410480
rect 4271 410469 4284 410480
rect 4024 408093 4072 410469
rect 4282 408093 4330 410469
rect 4086 408000 4268 408034
rect 4086 407892 4268 407926
rect 4070 407833 4072 407844
rect 4271 407833 4284 407844
rect 4024 405457 4072 407833
rect 4282 405457 4330 407833
rect 4086 405364 4268 405398
rect 4086 405256 4268 405290
rect 4070 405197 4072 405208
rect 4271 405197 4284 405208
rect 4024 402821 4072 405197
rect 4282 402821 4330 405197
rect 4086 402728 4268 402762
rect 4086 402620 4268 402654
rect 4070 402561 4072 402572
rect 4271 402561 4284 402572
rect 4024 400185 4072 402561
rect 4282 400185 4330 402561
rect 4086 400092 4268 400126
rect 4086 399984 4268 400018
rect 4070 399925 4072 399936
rect 4271 399925 4284 399936
rect 4024 397549 4072 399925
rect 4282 397549 4330 399925
rect 4086 397456 4268 397490
rect 4086 397348 4268 397382
rect 4070 397289 4072 397300
rect 4271 397289 4284 397300
rect 4024 394913 4072 397289
rect 4282 394913 4330 397289
rect 4086 394820 4268 394854
rect 4086 394712 4268 394746
rect 4070 394653 4072 394664
rect 4271 394653 4284 394664
rect 4024 392277 4072 394653
rect 4282 392277 4330 394653
rect 4086 392184 4268 392218
rect 4086 392076 4268 392110
rect 4070 392017 4072 392028
rect 4271 392017 4284 392028
rect 4024 389641 4072 392017
rect 4282 389641 4330 392017
rect 4086 389548 4268 389582
rect 4086 389440 4268 389474
rect 4070 389381 4072 389392
rect 4271 389381 4284 389392
rect 4024 387005 4072 389381
rect 4282 387005 4330 389381
rect 4086 386912 4268 386946
rect 4086 386804 4268 386838
rect 4070 386745 4072 386756
rect 4271 386745 4284 386756
rect 4024 384369 4072 386745
rect 4282 384369 4330 386745
rect 4086 384276 4268 384310
rect 4086 384168 4268 384202
rect 4070 384109 4072 384120
rect 4271 384109 4284 384120
rect 4024 381733 4072 384109
rect 4282 381733 4330 384109
rect 4086 381640 4268 381674
rect 4086 381532 4268 381566
rect 4070 381473 4072 381484
rect 4271 381473 4284 381484
rect 4024 379097 4072 381473
rect 4282 379097 4330 381473
rect 4086 379004 4268 379038
rect 4086 378896 4268 378930
rect 4070 378837 4072 378848
rect 4271 378837 4284 378848
rect 4024 376461 4072 378837
rect 4282 376461 4330 378837
rect 4086 376368 4268 376402
rect 4086 376260 4268 376294
rect 4070 376201 4072 376212
rect 4271 376201 4284 376212
rect 4024 373825 4072 376201
rect 4282 373825 4330 376201
rect 4086 373732 4268 373766
rect 4086 373624 4268 373658
rect 4070 373565 4072 373576
rect 4271 373565 4284 373576
rect 4024 371189 4072 373565
rect 4282 371189 4330 373565
rect 4086 371096 4268 371130
rect 4086 370988 4268 371022
rect 4070 370929 4072 370940
rect 4271 370929 4284 370940
rect 4024 368553 4072 370929
rect 4282 368553 4330 370929
rect 4086 368460 4268 368494
rect 4086 368352 4268 368386
rect 4070 368293 4072 368304
rect 4271 368293 4284 368304
rect 4024 365917 4072 368293
rect 4282 365917 4330 368293
rect 4086 365824 4268 365858
rect 4086 365716 4268 365750
rect 4070 365657 4072 365668
rect 4271 365657 4284 365668
rect 4024 363281 4072 365657
rect 4282 363281 4330 365657
rect 4086 363188 4268 363222
rect 4086 363080 4268 363114
rect 4070 363021 4072 363032
rect 4271 363021 4284 363032
rect 4024 360645 4072 363021
rect 4282 360645 4330 363021
rect 4086 360552 4268 360586
rect 4086 360444 4268 360478
rect 4070 360385 4072 360396
rect 4271 360385 4284 360396
rect 4024 358009 4072 360385
rect 4282 358009 4330 360385
rect 4086 357916 4268 357950
rect 4086 357808 4268 357842
rect 4070 357749 4072 357760
rect 4271 357749 4284 357760
rect 4024 355373 4072 357749
rect 4282 355373 4330 357749
rect 4086 355280 4268 355314
rect 4086 355172 4268 355206
rect 4070 355113 4072 355124
rect 4271 355113 4284 355124
rect 4024 352737 4072 355113
rect 4282 352737 4330 355113
rect 4086 352644 4268 352678
rect 4086 352536 4268 352570
rect 4070 352477 4072 352488
rect 4271 352477 4284 352488
rect 4024 350101 4072 352477
rect 4282 350101 4330 352477
rect 4086 350008 4268 350042
rect 4086 349900 4268 349934
rect 4070 349841 4072 349852
rect 4271 349841 4284 349852
rect 3365 348709 3747 348743
rect 3824 348647 3855 348755
rect 3269 190583 3317 348647
rect 3465 348571 3647 348605
rect 3449 348512 3451 348523
rect 3650 348512 3663 348523
rect 3403 347336 3451 348512
rect 3661 347336 3709 348512
rect 3465 347243 3647 347277
rect 3465 347135 3647 347169
rect 3449 347076 3451 347087
rect 3650 347076 3663 347087
rect 3403 345900 3451 347076
rect 3661 345900 3709 347076
rect 3465 345807 3647 345841
rect 3465 345699 3647 345733
rect 3449 345640 3451 345651
rect 3650 345640 3663 345651
rect 3403 344464 3451 345640
rect 3661 344464 3709 345640
rect 3465 344371 3647 344405
rect 3465 344263 3647 344297
rect 3449 344204 3451 344215
rect 3650 344204 3663 344215
rect 3403 343028 3451 344204
rect 3661 343028 3709 344204
rect 3795 344118 3855 348647
rect 3878 344118 3938 348809
rect 4024 347465 4072 349841
rect 4282 347465 4330 349841
rect 4086 347372 4268 347406
rect 4086 347264 4268 347298
rect 4070 347205 4072 347216
rect 4271 347205 4284 347216
rect 4024 344829 4072 347205
rect 4282 344829 4330 347205
rect 4086 344736 4268 344770
rect 4086 344628 4268 344662
rect 4070 344569 4072 344580
rect 4271 344569 4284 344580
rect 4024 344118 4072 344569
rect 4282 344118 4330 344569
rect 4416 344118 4464 655752
rect 3795 344053 4481 344118
rect 3465 342935 3647 342969
rect 3465 342827 3647 342861
rect 3449 342768 3451 342779
rect 3650 342768 3663 342779
rect 3403 341592 3451 342768
rect 3661 341592 3709 342768
rect 3465 341499 3647 341533
rect 3465 341391 3647 341425
rect 3449 341332 3451 341343
rect 3650 341332 3663 341343
rect 3403 340156 3451 341332
rect 3661 340156 3709 341332
rect 3465 340063 3647 340097
rect 3465 339955 3647 339989
rect 3449 339896 3451 339907
rect 3650 339896 3663 339907
rect 3403 338720 3451 339896
rect 3661 338720 3709 339896
rect 3465 338627 3647 338661
rect 3465 338519 3647 338553
rect 3449 338460 3451 338471
rect 3650 338460 3663 338471
rect 3403 337284 3451 338460
rect 3661 337284 3709 338460
rect 3465 337191 3647 337225
rect 3465 337083 3647 337117
rect 3449 337024 3451 337035
rect 3650 337024 3663 337035
rect 3403 335848 3451 337024
rect 3661 335848 3709 337024
rect 3465 335755 3647 335789
rect 3465 335647 3647 335681
rect 3449 335588 3451 335599
rect 3650 335588 3663 335599
rect 3403 334412 3451 335588
rect 3661 334412 3709 335588
rect 3465 334319 3647 334353
rect 3465 334211 3647 334245
rect 3449 334152 3451 334163
rect 3650 334152 3663 334163
rect 3403 332976 3451 334152
rect 3661 332976 3709 334152
rect 3465 332883 3647 332917
rect 3465 332775 3647 332809
rect 3449 332716 3451 332727
rect 3650 332716 3663 332727
rect 3403 331540 3451 332716
rect 3661 331540 3709 332716
rect 3465 331447 3647 331481
rect 3465 331339 3647 331373
rect 3449 331280 3451 331291
rect 3650 331280 3663 331291
rect 3403 330104 3451 331280
rect 3661 330104 3709 331280
rect 3465 330011 3647 330045
rect 3465 329903 3647 329937
rect 3449 329844 3451 329855
rect 3650 329844 3663 329855
rect 3403 328668 3451 329844
rect 3661 328668 3709 329844
rect 3465 328575 3647 328609
rect 3465 328467 3647 328501
rect 3449 328408 3451 328419
rect 3650 328408 3663 328419
rect 3403 327232 3451 328408
rect 3661 327232 3709 328408
rect 3465 327139 3647 327173
rect 3465 327031 3647 327065
rect 3449 326972 3451 326983
rect 3650 326972 3663 326983
rect 3403 325796 3451 326972
rect 3661 325796 3709 326972
rect 3465 325703 3647 325737
rect 3465 325595 3647 325629
rect 3449 325536 3451 325547
rect 3650 325536 3663 325547
rect 3403 324360 3451 325536
rect 3661 324360 3709 325536
rect 3465 324267 3647 324301
rect 3465 324159 3647 324193
rect 3449 324100 3451 324111
rect 3650 324100 3663 324111
rect 3403 322924 3451 324100
rect 3661 322924 3709 324100
rect 3465 322831 3647 322865
rect 3465 322723 3647 322757
rect 3449 322664 3451 322675
rect 3650 322664 3663 322675
rect 3403 321488 3451 322664
rect 3661 321488 3709 322664
rect 3465 321395 3647 321429
rect 3465 321287 3647 321321
rect 3449 321228 3451 321239
rect 3650 321228 3663 321239
rect 3403 320052 3451 321228
rect 3661 320052 3709 321228
rect 3465 319959 3647 319993
rect 3465 319851 3647 319885
rect 3449 319792 3451 319803
rect 3650 319792 3663 319803
rect 3403 318616 3451 319792
rect 3661 318616 3709 319792
rect 3465 318523 3647 318557
rect 3465 318415 3647 318449
rect 3449 318356 3451 318367
rect 3650 318356 3663 318367
rect 3403 317180 3451 318356
rect 3661 317180 3709 318356
rect 3465 317087 3647 317121
rect 3465 316979 3647 317013
rect 3449 316920 3451 316931
rect 3650 316920 3663 316931
rect 3403 315744 3451 316920
rect 3661 315744 3709 316920
rect 3465 315651 3647 315685
rect 3465 315543 3647 315577
rect 3449 315484 3451 315495
rect 3650 315484 3663 315495
rect 3403 314308 3451 315484
rect 3661 314308 3709 315484
rect 3465 314215 3647 314249
rect 3465 314107 3647 314141
rect 3449 314048 3451 314059
rect 3650 314048 3663 314059
rect 3403 312872 3451 314048
rect 3661 312872 3709 314048
rect 3465 312779 3647 312813
rect 3465 312671 3647 312705
rect 3449 312612 3451 312623
rect 3650 312612 3663 312623
rect 3403 311436 3451 312612
rect 3661 311436 3709 312612
rect 3465 311343 3647 311377
rect 3465 311235 3647 311269
rect 3449 311176 3451 311187
rect 3650 311176 3663 311187
rect 3403 310000 3451 311176
rect 3661 310000 3709 311176
rect 3465 309907 3647 309941
rect 3465 309799 3647 309833
rect 3449 309740 3451 309751
rect 3650 309740 3663 309751
rect 3403 308564 3451 309740
rect 3661 308564 3709 309740
rect 3465 308471 3647 308505
rect 3465 308363 3647 308397
rect 3449 308304 3451 308315
rect 3650 308304 3663 308315
rect 3403 307128 3451 308304
rect 3661 307128 3709 308304
rect 3465 307035 3647 307069
rect 3465 306927 3647 306961
rect 3449 306868 3451 306879
rect 3650 306868 3663 306879
rect 3403 305692 3451 306868
rect 3661 305692 3709 306868
rect 3465 305599 3647 305633
rect 3465 305491 3647 305525
rect 3449 305432 3451 305443
rect 3650 305432 3663 305443
rect 3403 304256 3451 305432
rect 3661 304256 3709 305432
rect 3465 304163 3647 304197
rect 3465 304055 3647 304089
rect 3449 303996 3451 304007
rect 3650 303996 3663 304007
rect 3403 302820 3451 303996
rect 3661 302820 3709 303996
rect 3465 302727 3647 302761
rect 3465 302619 3647 302653
rect 3449 302560 3451 302571
rect 3650 302560 3663 302571
rect 3403 301384 3451 302560
rect 3661 301384 3709 302560
rect 3465 301291 3647 301325
rect 3465 301183 3647 301217
rect 3449 301124 3451 301135
rect 3650 301124 3663 301135
rect 3403 299948 3451 301124
rect 3661 299948 3709 301124
rect 3465 299855 3647 299889
rect 3465 299747 3647 299781
rect 3449 299688 3451 299699
rect 3650 299688 3663 299699
rect 3403 298512 3451 299688
rect 3661 298512 3709 299688
rect 3465 298419 3647 298453
rect 3465 298311 3647 298345
rect 3449 298252 3451 298263
rect 3650 298252 3663 298263
rect 3403 297076 3451 298252
rect 3661 297076 3709 298252
rect 3465 296983 3647 297017
rect 3465 296875 3647 296909
rect 3449 296816 3451 296827
rect 3650 296816 3663 296827
rect 3403 295640 3451 296816
rect 3661 295640 3709 296816
rect 3465 295547 3647 295581
rect 3465 295439 3647 295473
rect 3449 295380 3451 295391
rect 3650 295380 3663 295391
rect 3403 294204 3451 295380
rect 3661 294204 3709 295380
rect 3465 294111 3647 294145
rect 3465 294003 3647 294037
rect 3449 293944 3451 293955
rect 3650 293944 3663 293955
rect 3403 292768 3451 293944
rect 3661 292768 3709 293944
rect 3465 292675 3647 292709
rect 3465 292567 3647 292601
rect 3449 292508 3451 292519
rect 3650 292508 3663 292519
rect 3403 291332 3451 292508
rect 3661 291332 3709 292508
rect 3465 291239 3647 291273
rect 3465 291131 3647 291165
rect 3449 291072 3451 291083
rect 3650 291072 3663 291083
rect 3403 289896 3451 291072
rect 3661 289896 3709 291072
rect 3465 289803 3647 289837
rect 3465 289695 3647 289729
rect 3449 289636 3451 289647
rect 3650 289636 3663 289647
rect 3403 288460 3451 289636
rect 3661 288460 3709 289636
rect 3465 288367 3647 288401
rect 3465 288259 3647 288293
rect 3449 288200 3451 288211
rect 3650 288200 3663 288211
rect 3403 287024 3451 288200
rect 3661 287024 3709 288200
rect 3465 286931 3647 286965
rect 3465 286823 3647 286857
rect 3449 286764 3451 286775
rect 3650 286764 3663 286775
rect 3403 285588 3451 286764
rect 3661 285588 3709 286764
rect 3465 285495 3647 285529
rect 3465 285387 3647 285421
rect 3449 285328 3451 285339
rect 3650 285328 3663 285339
rect 3403 284152 3451 285328
rect 3661 284152 3709 285328
rect 3465 284059 3647 284093
rect 3465 283951 3647 283985
rect 3449 283892 3451 283903
rect 3650 283892 3663 283903
rect 3403 282716 3451 283892
rect 3661 282716 3709 283892
rect 3465 282623 3647 282657
rect 3465 282515 3647 282549
rect 3449 282456 3451 282467
rect 3650 282456 3663 282467
rect 3403 281280 3451 282456
rect 3661 281280 3709 282456
rect 3465 281187 3647 281221
rect 3465 281079 3647 281113
rect 3449 281020 3451 281031
rect 3650 281020 3663 281031
rect 3403 279844 3451 281020
rect 3661 279844 3709 281020
rect 3465 279751 3647 279785
rect 3465 279643 3647 279677
rect 3449 279584 3451 279595
rect 3650 279584 3663 279595
rect 3403 278408 3451 279584
rect 3661 278408 3709 279584
rect 3465 278315 3647 278349
rect 3465 278207 3647 278241
rect 3449 278148 3451 278159
rect 3650 278148 3663 278159
rect 3403 276972 3451 278148
rect 3661 276972 3709 278148
rect 3465 276879 3647 276913
rect 3465 276771 3647 276805
rect 3449 276712 3451 276723
rect 3650 276712 3663 276723
rect 3403 275536 3451 276712
rect 3661 275536 3709 276712
rect 3465 275443 3647 275477
rect 3465 275335 3647 275369
rect 3449 275276 3451 275287
rect 3650 275276 3663 275287
rect 3403 274100 3451 275276
rect 3661 274100 3709 275276
rect 3465 274007 3647 274041
rect 3465 273899 3647 273933
rect 3449 273840 3451 273851
rect 3650 273840 3663 273851
rect 3403 272664 3451 273840
rect 3661 272664 3709 273840
rect 3465 272571 3647 272605
rect 3465 272463 3647 272497
rect 3449 272404 3451 272415
rect 3650 272404 3663 272415
rect 3403 271228 3451 272404
rect 3661 271228 3709 272404
rect 3465 271135 3647 271169
rect 3465 271027 3647 271061
rect 3449 270968 3451 270979
rect 3650 270968 3663 270979
rect 3403 269792 3451 270968
rect 3661 269792 3709 270968
rect 3465 269699 3647 269733
rect 3465 269591 3647 269625
rect 3449 269532 3451 269543
rect 3650 269532 3663 269543
rect 3403 268356 3451 269532
rect 3661 268356 3709 269532
rect 3465 268263 3647 268297
rect 3465 268155 3647 268189
rect 3449 268096 3451 268107
rect 3650 268096 3663 268107
rect 3403 266920 3451 268096
rect 3661 266920 3709 268096
rect 3465 266827 3647 266861
rect 3465 266719 3647 266753
rect 3449 266660 3451 266671
rect 3650 266660 3663 266671
rect 3403 265484 3451 266660
rect 3661 265484 3709 266660
rect 3465 265391 3647 265425
rect 3465 265283 3647 265317
rect 3449 265224 3451 265235
rect 3650 265224 3663 265235
rect 3403 264048 3451 265224
rect 3661 264048 3709 265224
rect 3465 263955 3647 263989
rect 3465 263847 3647 263881
rect 3449 263788 3451 263799
rect 3650 263788 3663 263799
rect 3403 262612 3451 263788
rect 3661 262612 3709 263788
rect 3465 262519 3647 262553
rect 3465 262411 3647 262445
rect 3449 262352 3451 262363
rect 3650 262352 3663 262363
rect 3403 261176 3451 262352
rect 3661 261176 3709 262352
rect 3465 261083 3647 261117
rect 3465 260975 3647 261009
rect 3449 260916 3451 260927
rect 3650 260916 3663 260927
rect 3403 259740 3451 260916
rect 3661 259740 3709 260916
rect 3465 259647 3647 259681
rect 3465 259539 3647 259573
rect 3449 259480 3451 259491
rect 3650 259480 3663 259491
rect 3403 258304 3451 259480
rect 3661 258304 3709 259480
rect 3465 258211 3647 258245
rect 3465 258103 3647 258137
rect 3449 258044 3451 258055
rect 3650 258044 3663 258055
rect 3403 256868 3451 258044
rect 3661 256868 3709 258044
rect 3465 256775 3647 256809
rect 3465 256667 3647 256701
rect 3449 256608 3451 256619
rect 3650 256608 3663 256619
rect 3403 255432 3451 256608
rect 3661 255432 3709 256608
rect 3465 255339 3647 255373
rect 3465 255231 3647 255265
rect 3449 255172 3451 255183
rect 3650 255172 3663 255183
rect 3403 253996 3451 255172
rect 3661 253996 3709 255172
rect 3465 253903 3647 253937
rect 3465 253795 3647 253829
rect 3449 253736 3451 253747
rect 3650 253736 3663 253747
rect 3403 252560 3451 253736
rect 3661 252560 3709 253736
rect 3465 252467 3647 252501
rect 3465 252359 3647 252393
rect 3449 252300 3451 252311
rect 3650 252300 3663 252311
rect 3403 251124 3451 252300
rect 3661 251124 3709 252300
rect 3465 251031 3647 251065
rect 3465 250923 3647 250957
rect 3449 250864 3451 250875
rect 3650 250864 3663 250875
rect 3403 249688 3451 250864
rect 3661 249688 3709 250864
rect 3465 249595 3647 249629
rect 3465 249487 3647 249521
rect 3449 249428 3451 249439
rect 3650 249428 3663 249439
rect 3403 248252 3451 249428
rect 3661 248252 3709 249428
rect 3465 248159 3647 248193
rect 3465 248051 3647 248085
rect 3449 247992 3451 248003
rect 3650 247992 3663 248003
rect 3403 246816 3451 247992
rect 3661 246816 3709 247992
rect 3465 246723 3647 246757
rect 3465 246615 3647 246649
rect 3449 246556 3451 246567
rect 3650 246556 3663 246567
rect 3403 245380 3451 246556
rect 3661 245380 3709 246556
rect 3795 246231 4542 344053
rect 4546 343971 4928 344005
rect 5007 343909 5024 343971
rect 4976 343869 5024 343909
rect 4646 343833 4828 343867
rect 4572 343783 4584 343795
rect 4630 343783 4632 343794
rect 4831 343783 4844 343794
rect 4890 343783 4902 343795
rect 4572 342607 4632 343783
rect 4842 342607 4902 343783
rect 4572 342595 4584 342607
rect 4890 342595 4902 342607
rect 4646 342523 4828 342557
rect 4964 342521 5024 343869
rect 4976 342451 5024 342521
rect 4646 342415 4828 342449
rect 4572 342365 4584 342377
rect 4630 342365 4632 342376
rect 4831 342365 4844 342376
rect 4890 342365 4902 342377
rect 4572 341189 4632 342365
rect 4842 341189 4902 342365
rect 4572 341177 4584 341189
rect 4890 341177 4902 341189
rect 4646 341105 4828 341139
rect 4964 341103 5024 342451
rect 4976 341033 5024 341103
rect 4646 340997 4828 341031
rect 4572 340947 4584 340959
rect 4630 340947 4632 340958
rect 4831 340947 4844 340958
rect 4890 340947 4902 340959
rect 4572 339771 4632 340947
rect 4842 339771 4902 340947
rect 4572 339759 4584 339771
rect 4890 339759 4902 339771
rect 4646 339687 4828 339721
rect 4964 339685 5024 341033
rect 4976 339615 5024 339685
rect 4646 339579 4828 339613
rect 4572 339529 4584 339541
rect 4630 339529 4632 339540
rect 4831 339529 4844 339540
rect 4890 339529 4902 339541
rect 4572 338353 4632 339529
rect 4842 338353 4902 339529
rect 4572 338341 4584 338353
rect 4890 338341 4902 338353
rect 4646 338269 4828 338303
rect 4964 338267 5024 339615
rect 4976 338197 5024 338267
rect 4646 338161 4828 338195
rect 4572 338111 4584 338123
rect 4630 338111 4632 338122
rect 4831 338111 4844 338122
rect 4890 338111 4902 338123
rect 4572 336935 4632 338111
rect 4842 336935 4902 338111
rect 4572 336923 4584 336935
rect 4890 336923 4902 336935
rect 4646 336851 4828 336885
rect 4964 336849 5024 338197
rect 4976 336779 5024 336849
rect 4646 336743 4828 336777
rect 4572 336693 4584 336705
rect 4630 336693 4632 336704
rect 4831 336693 4844 336704
rect 4890 336693 4902 336705
rect 4572 335517 4632 336693
rect 4842 335517 4902 336693
rect 4572 335505 4584 335517
rect 4890 335505 4902 335517
rect 4646 335433 4828 335467
rect 4964 335431 5024 336779
rect 4976 335361 5024 335431
rect 4646 335325 4828 335359
rect 4572 335275 4584 335287
rect 4630 335275 4632 335286
rect 4831 335275 4844 335286
rect 4890 335275 4902 335287
rect 4572 334099 4632 335275
rect 4842 334099 4902 335275
rect 4572 334087 4584 334099
rect 4890 334087 4902 334099
rect 4646 334015 4828 334049
rect 4964 334013 5024 335361
rect 4976 333943 5024 334013
rect 4646 333907 4828 333941
rect 4572 333857 4584 333869
rect 4630 333857 4632 333868
rect 4831 333857 4844 333868
rect 4890 333857 4902 333869
rect 4572 332681 4632 333857
rect 4842 332681 4902 333857
rect 4572 332669 4584 332681
rect 4890 332669 4902 332681
rect 4646 332597 4828 332631
rect 4964 332595 5024 333943
rect 4976 332525 5024 332595
rect 4646 332489 4828 332523
rect 4572 332439 4584 332451
rect 4630 332439 4632 332450
rect 4831 332439 4844 332450
rect 4890 332439 4902 332451
rect 4572 331263 4632 332439
rect 4842 331263 4902 332439
rect 4572 331251 4584 331263
rect 4890 331251 4902 331263
rect 4646 331179 4828 331213
rect 4964 331177 5024 332525
rect 4976 331107 5024 331177
rect 4646 331071 4828 331105
rect 4572 331021 4584 331033
rect 4630 331021 4632 331032
rect 4831 331021 4844 331032
rect 4890 331021 4902 331033
rect 4572 329845 4632 331021
rect 4842 329845 4902 331021
rect 4572 329833 4584 329845
rect 4890 329833 4902 329845
rect 4646 329761 4828 329795
rect 4964 329759 5024 331107
rect 4976 329689 5024 329759
rect 4646 329653 4828 329687
rect 4572 329603 4584 329615
rect 4630 329603 4632 329614
rect 4831 329603 4844 329614
rect 4890 329603 4902 329615
rect 4572 328427 4632 329603
rect 4842 328427 4902 329603
rect 4572 328415 4584 328427
rect 4890 328415 4902 328427
rect 4646 328343 4828 328377
rect 4964 328341 5024 329689
rect 4976 328271 5024 328341
rect 4646 328235 4828 328269
rect 4572 328185 4584 328197
rect 4630 328185 4632 328196
rect 4831 328185 4844 328196
rect 4890 328185 4902 328197
rect 4572 327009 4632 328185
rect 4842 327009 4902 328185
rect 4572 326997 4584 327009
rect 4890 326997 4902 327009
rect 4646 326925 4828 326959
rect 4964 326923 5024 328271
rect 4976 326853 5024 326923
rect 4646 326817 4828 326851
rect 4572 326767 4584 326779
rect 4630 326767 4632 326778
rect 4831 326767 4844 326778
rect 4890 326767 4902 326779
rect 4572 325591 4632 326767
rect 4842 325591 4902 326767
rect 4572 325579 4584 325591
rect 4890 325579 4902 325591
rect 4646 325507 4828 325541
rect 4964 325505 5024 326853
rect 4976 325435 5024 325505
rect 4646 325399 4828 325433
rect 4572 325349 4584 325361
rect 4630 325349 4632 325360
rect 4831 325349 4844 325360
rect 4890 325349 4902 325361
rect 4572 324173 4632 325349
rect 4842 324173 4902 325349
rect 4572 324161 4584 324173
rect 4890 324161 4902 324173
rect 4646 324089 4828 324123
rect 4964 324087 5024 325435
rect 4976 324017 5024 324087
rect 4646 323981 4828 324015
rect 4572 323931 4584 323943
rect 4630 323931 4632 323942
rect 4831 323931 4844 323942
rect 4890 323931 4902 323943
rect 4572 322755 4632 323931
rect 4842 322755 4902 323931
rect 4572 322743 4584 322755
rect 4890 322743 4902 322755
rect 4646 322671 4828 322705
rect 4964 322669 5024 324017
rect 4976 322599 5024 322669
rect 4646 322563 4828 322597
rect 4572 322513 4584 322525
rect 4630 322513 4632 322524
rect 4831 322513 4844 322524
rect 4890 322513 4902 322525
rect 4572 321337 4632 322513
rect 4842 321337 4902 322513
rect 4572 321325 4584 321337
rect 4890 321325 4902 321337
rect 4646 321253 4828 321287
rect 4964 321251 5024 322599
rect 4976 321181 5024 321251
rect 4646 321145 4828 321179
rect 4572 321095 4584 321107
rect 4630 321095 4632 321106
rect 4831 321095 4844 321106
rect 4890 321095 4902 321107
rect 4572 319919 4632 321095
rect 4842 319919 4902 321095
rect 4572 319907 4584 319919
rect 4890 319907 4902 319919
rect 4646 319835 4828 319869
rect 4964 319833 5024 321181
rect 4976 319763 5024 319833
rect 4646 319727 4828 319761
rect 4572 319677 4584 319689
rect 4630 319677 4632 319688
rect 4831 319677 4844 319688
rect 4890 319677 4902 319689
rect 4572 318501 4632 319677
rect 4842 318501 4902 319677
rect 4572 318489 4584 318501
rect 4890 318489 4902 318501
rect 4646 318417 4828 318451
rect 4964 318415 5024 319763
rect 4976 318345 5024 318415
rect 4646 318309 4828 318343
rect 4572 318259 4584 318271
rect 4630 318259 4632 318270
rect 4831 318259 4844 318270
rect 4890 318259 4902 318271
rect 4572 317083 4632 318259
rect 4842 317083 4902 318259
rect 4572 317071 4584 317083
rect 4890 317071 4902 317083
rect 4646 316999 4828 317033
rect 4964 316997 5024 318345
rect 4976 316927 5024 316997
rect 4646 316891 4828 316925
rect 4572 316841 4584 316853
rect 4630 316841 4632 316852
rect 4831 316841 4844 316852
rect 4890 316841 4902 316853
rect 4572 315665 4632 316841
rect 4842 315665 4902 316841
rect 4572 315653 4584 315665
rect 4890 315653 4902 315665
rect 4646 315581 4828 315615
rect 4964 315579 5024 316927
rect 4976 315509 5024 315579
rect 4646 315473 4828 315507
rect 4572 315423 4584 315435
rect 4630 315423 4632 315434
rect 4831 315423 4844 315434
rect 4890 315423 4902 315435
rect 4572 314247 4632 315423
rect 4842 314247 4902 315423
rect 4572 314235 4584 314247
rect 4890 314235 4902 314247
rect 4646 314163 4828 314197
rect 4964 314161 5024 315509
rect 4976 314091 5024 314161
rect 4646 314055 4828 314089
rect 4572 314005 4584 314017
rect 4630 314005 4632 314016
rect 4831 314005 4844 314016
rect 4890 314005 4902 314017
rect 4572 312829 4632 314005
rect 4842 312829 4902 314005
rect 4572 312817 4584 312829
rect 4890 312817 4902 312829
rect 4646 312745 4828 312779
rect 4964 312743 5024 314091
rect 4976 312673 5024 312743
rect 4646 312637 4828 312671
rect 4572 312587 4584 312599
rect 4630 312587 4632 312598
rect 4831 312587 4844 312598
rect 4890 312587 4902 312599
rect 4572 311411 4632 312587
rect 4842 311411 4902 312587
rect 4572 311399 4584 311411
rect 4890 311399 4902 311411
rect 4646 311327 4828 311361
rect 4964 311325 5024 312673
rect 4976 311255 5024 311325
rect 4646 311219 4828 311253
rect 4572 311169 4584 311181
rect 4630 311169 4632 311180
rect 4831 311169 4844 311180
rect 4890 311169 4902 311181
rect 4572 309993 4632 311169
rect 4842 309993 4902 311169
rect 4572 309981 4584 309993
rect 4890 309981 4902 309993
rect 4646 309909 4828 309943
rect 4964 309907 5024 311255
rect 4976 309837 5024 309907
rect 4646 309801 4828 309835
rect 4572 309751 4584 309763
rect 4630 309751 4632 309762
rect 4831 309751 4844 309762
rect 4890 309751 4902 309763
rect 4572 308575 4632 309751
rect 4842 308575 4902 309751
rect 4572 308563 4584 308575
rect 4890 308563 4902 308575
rect 4646 308491 4828 308525
rect 4964 308489 5024 309837
rect 4976 308419 5024 308489
rect 4646 308383 4828 308417
rect 4572 308333 4584 308345
rect 4630 308333 4632 308344
rect 4831 308333 4844 308344
rect 4890 308333 4902 308345
rect 4572 307157 4632 308333
rect 4842 307157 4902 308333
rect 4572 307145 4584 307157
rect 4890 307145 4902 307157
rect 4646 307073 4828 307107
rect 4964 307071 5024 308419
rect 4976 307001 5024 307071
rect 4646 306965 4828 306999
rect 4572 306915 4584 306927
rect 4630 306915 4632 306926
rect 4831 306915 4844 306926
rect 4890 306915 4902 306927
rect 4572 305739 4632 306915
rect 4842 305739 4902 306915
rect 4572 305727 4584 305739
rect 4890 305727 4902 305739
rect 4646 305655 4828 305689
rect 4964 305653 5024 307001
rect 4976 305583 5024 305653
rect 4646 305547 4828 305581
rect 4572 305497 4584 305509
rect 4630 305497 4632 305508
rect 4831 305497 4844 305508
rect 4890 305497 4902 305509
rect 4572 304321 4632 305497
rect 4842 304321 4902 305497
rect 4572 304309 4584 304321
rect 4890 304309 4902 304321
rect 4646 304237 4828 304271
rect 4964 304235 5024 305583
rect 4976 304165 5024 304235
rect 4646 304129 4828 304163
rect 4572 304079 4584 304091
rect 4630 304079 4632 304090
rect 4831 304079 4844 304090
rect 4890 304079 4902 304091
rect 4572 302903 4632 304079
rect 4842 302903 4902 304079
rect 4572 302891 4584 302903
rect 4890 302891 4902 302903
rect 4646 302819 4828 302853
rect 4964 302817 5024 304165
rect 4976 302747 5024 302817
rect 4646 302711 4828 302745
rect 4572 302661 4584 302673
rect 4630 302661 4632 302672
rect 4831 302661 4844 302672
rect 4890 302661 4902 302673
rect 4572 301485 4632 302661
rect 4842 301485 4902 302661
rect 4572 301473 4584 301485
rect 4890 301473 4902 301485
rect 4646 301401 4828 301435
rect 4964 301399 5024 302747
rect 4976 301329 5024 301399
rect 4646 301293 4828 301327
rect 4572 301243 4584 301255
rect 4630 301243 4632 301254
rect 4831 301243 4844 301254
rect 4890 301243 4902 301255
rect 4572 300067 4632 301243
rect 4842 300067 4902 301243
rect 4572 300055 4584 300067
rect 4890 300055 4902 300067
rect 4646 299983 4828 300017
rect 4964 299981 5024 301329
rect 4976 299911 5024 299981
rect 4646 299875 4828 299909
rect 4572 299825 4584 299837
rect 4630 299825 4632 299836
rect 4831 299825 4844 299836
rect 4890 299825 4902 299837
rect 4572 298649 4632 299825
rect 4842 298649 4902 299825
rect 4572 298637 4584 298649
rect 4890 298637 4902 298649
rect 4646 298565 4828 298599
rect 4964 298563 5024 299911
rect 4976 298493 5024 298563
rect 4646 298457 4828 298491
rect 4572 298407 4584 298419
rect 4630 298407 4632 298418
rect 4831 298407 4844 298418
rect 4890 298407 4902 298419
rect 4572 297231 4632 298407
rect 4842 297231 4902 298407
rect 4572 297219 4584 297231
rect 4890 297219 4902 297231
rect 4646 297147 4828 297181
rect 4964 297145 5024 298493
rect 4976 297075 5024 297145
rect 4646 297039 4828 297073
rect 4572 296989 4584 297001
rect 4630 296989 4632 297000
rect 4831 296989 4844 297000
rect 4890 296989 4902 297001
rect 4572 295813 4632 296989
rect 4842 295813 4902 296989
rect 4572 295801 4584 295813
rect 4890 295801 4902 295813
rect 4646 295729 4828 295763
rect 4964 295727 5024 297075
rect 4976 295657 5024 295727
rect 4646 295621 4828 295655
rect 4572 295571 4584 295583
rect 4630 295571 4632 295582
rect 4831 295571 4844 295582
rect 4890 295571 4902 295583
rect 4572 294395 4632 295571
rect 4842 294395 4902 295571
rect 4572 294383 4584 294395
rect 4890 294383 4902 294395
rect 4646 294311 4828 294345
rect 4964 294309 5024 295657
rect 4976 294239 5024 294309
rect 4646 294203 4828 294237
rect 4572 294153 4584 294165
rect 4630 294153 4632 294164
rect 4831 294153 4844 294164
rect 4890 294153 4902 294165
rect 4572 292977 4632 294153
rect 4842 292977 4902 294153
rect 4572 292965 4584 292977
rect 4890 292965 4902 292977
rect 4646 292893 4828 292927
rect 4964 292891 5024 294239
rect 4976 292821 5024 292891
rect 4646 292785 4828 292819
rect 4572 292735 4584 292747
rect 4630 292735 4632 292746
rect 4831 292735 4844 292746
rect 4890 292735 4902 292747
rect 4572 291559 4632 292735
rect 4842 291559 4902 292735
rect 4572 291547 4584 291559
rect 4890 291547 4902 291559
rect 4646 291475 4828 291509
rect 4964 291473 5024 292821
rect 4976 291403 5024 291473
rect 4646 291367 4828 291401
rect 4572 291317 4584 291329
rect 4630 291317 4632 291328
rect 4831 291317 4844 291328
rect 4890 291317 4902 291329
rect 4572 290141 4632 291317
rect 4842 290141 4902 291317
rect 4572 290129 4584 290141
rect 4890 290129 4902 290141
rect 4646 290057 4828 290091
rect 4964 290055 5024 291403
rect 4976 289985 5024 290055
rect 4646 289949 4828 289983
rect 4572 289899 4584 289911
rect 4630 289899 4632 289910
rect 4831 289899 4844 289910
rect 4890 289899 4902 289911
rect 4572 288723 4632 289899
rect 4842 288723 4902 289899
rect 4572 288711 4584 288723
rect 4890 288711 4902 288723
rect 4646 288639 4828 288673
rect 4964 288637 5024 289985
rect 4976 288567 5024 288637
rect 4646 288531 4828 288565
rect 4572 288481 4584 288493
rect 4630 288481 4632 288492
rect 4831 288481 4844 288492
rect 4890 288481 4902 288493
rect 4572 287305 4632 288481
rect 4842 287305 4902 288481
rect 4572 287293 4584 287305
rect 4890 287293 4902 287305
rect 4646 287221 4828 287255
rect 4964 287219 5024 288567
rect 4976 287149 5024 287219
rect 4646 287113 4828 287147
rect 4572 287063 4584 287075
rect 4630 287063 4632 287074
rect 4831 287063 4844 287074
rect 4890 287063 4902 287075
rect 4572 285887 4632 287063
rect 4842 285887 4902 287063
rect 4572 285875 4584 285887
rect 4890 285875 4902 285887
rect 4646 285803 4828 285837
rect 4964 285801 5024 287149
rect 4976 285731 5024 285801
rect 4646 285695 4828 285729
rect 4572 285645 4584 285657
rect 4630 285645 4632 285656
rect 4831 285645 4844 285656
rect 4890 285645 4902 285657
rect 4572 284469 4632 285645
rect 4842 284469 4902 285645
rect 4572 284457 4584 284469
rect 4890 284457 4902 284469
rect 4646 284385 4828 284419
rect 4964 284383 5024 285731
rect 4976 284313 5024 284383
rect 4646 284277 4828 284311
rect 4572 284227 4584 284239
rect 4630 284227 4632 284238
rect 4831 284227 4844 284238
rect 4890 284227 4902 284239
rect 4572 283051 4632 284227
rect 4842 283051 4902 284227
rect 4572 283039 4584 283051
rect 4890 283039 4902 283051
rect 4646 282967 4828 283001
rect 4964 282965 5024 284313
rect 4976 282895 5024 282965
rect 4646 282859 4828 282893
rect 4572 282809 4584 282821
rect 4630 282809 4632 282820
rect 4831 282809 4844 282820
rect 4890 282809 4902 282821
rect 4572 281633 4632 282809
rect 4842 281633 4902 282809
rect 4572 281621 4584 281633
rect 4890 281621 4902 281633
rect 4646 281549 4828 281583
rect 4964 281547 5024 282895
rect 4976 281477 5024 281547
rect 4646 281441 4828 281475
rect 4572 281391 4584 281403
rect 4630 281391 4632 281402
rect 4831 281391 4844 281402
rect 4890 281391 4902 281403
rect 4572 280215 4632 281391
rect 4842 280215 4902 281391
rect 4572 280203 4584 280215
rect 4890 280203 4902 280215
rect 4646 280131 4828 280165
rect 4964 280129 5024 281477
rect 4976 280059 5024 280129
rect 4646 280023 4828 280057
rect 4572 279973 4584 279985
rect 4630 279973 4632 279984
rect 4831 279973 4844 279984
rect 4890 279973 4902 279985
rect 4572 278797 4632 279973
rect 4842 278797 4902 279973
rect 4572 278785 4584 278797
rect 4890 278785 4902 278797
rect 4646 278713 4828 278747
rect 4964 278711 5024 280059
rect 4976 278641 5024 278711
rect 4646 278605 4828 278639
rect 4572 278555 4584 278567
rect 4630 278555 4632 278566
rect 4831 278555 4844 278566
rect 4890 278555 4902 278567
rect 4572 277379 4632 278555
rect 4842 277379 4902 278555
rect 4572 277367 4584 277379
rect 4890 277367 4902 277379
rect 4646 277295 4828 277329
rect 4964 277293 5024 278641
rect 4976 277223 5024 277293
rect 4646 277187 4828 277221
rect 4572 277137 4584 277149
rect 4630 277137 4632 277148
rect 4831 277137 4844 277148
rect 4890 277137 4902 277149
rect 4572 275961 4632 277137
rect 4842 275961 4902 277137
rect 4572 275949 4584 275961
rect 4890 275949 4902 275961
rect 4646 275877 4828 275911
rect 4964 275875 5024 277223
rect 4976 275805 5024 275875
rect 4646 275769 4828 275803
rect 4572 275719 4584 275731
rect 4630 275719 4632 275730
rect 4831 275719 4844 275730
rect 4890 275719 4902 275731
rect 4572 274543 4632 275719
rect 4842 274543 4902 275719
rect 4572 274531 4584 274543
rect 4890 274531 4902 274543
rect 4646 274459 4828 274493
rect 4964 274457 5024 275805
rect 4976 274387 5024 274457
rect 4646 274351 4828 274385
rect 4572 274301 4584 274313
rect 4630 274301 4632 274312
rect 4831 274301 4844 274312
rect 4890 274301 4902 274313
rect 4572 273125 4632 274301
rect 4842 273125 4902 274301
rect 4572 273113 4584 273125
rect 4890 273113 4902 273125
rect 4646 273041 4828 273075
rect 4964 273039 5024 274387
rect 4976 272969 5024 273039
rect 4646 272933 4828 272967
rect 4572 272883 4584 272895
rect 4630 272883 4632 272894
rect 4831 272883 4844 272894
rect 4890 272883 4902 272895
rect 4572 271707 4632 272883
rect 4842 271707 4902 272883
rect 4572 271695 4584 271707
rect 4890 271695 4902 271707
rect 4646 271623 4828 271657
rect 4964 271621 5024 272969
rect 4976 271551 5024 271621
rect 4646 271515 4828 271549
rect 4572 271465 4584 271477
rect 4630 271465 4632 271476
rect 4831 271465 4844 271476
rect 4890 271465 4902 271477
rect 4572 270289 4632 271465
rect 4842 270289 4902 271465
rect 4572 270277 4584 270289
rect 4890 270277 4902 270289
rect 4646 270205 4828 270239
rect 4964 270203 5024 271551
rect 4976 270133 5024 270203
rect 4646 270097 4828 270131
rect 4572 270047 4584 270059
rect 4630 270047 4632 270058
rect 4831 270047 4844 270058
rect 4890 270047 4902 270059
rect 4572 268871 4632 270047
rect 4842 268871 4902 270047
rect 4572 268859 4584 268871
rect 4890 268859 4902 268871
rect 4646 268787 4828 268821
rect 4964 268785 5024 270133
rect 4976 268715 5024 268785
rect 4646 268679 4828 268713
rect 4572 268629 4584 268641
rect 4630 268629 4632 268640
rect 4831 268629 4844 268640
rect 4890 268629 4902 268641
rect 4572 267453 4632 268629
rect 4842 267453 4902 268629
rect 4572 267441 4584 267453
rect 4890 267441 4902 267453
rect 4646 267369 4828 267403
rect 4964 267367 5024 268715
rect 4976 267297 5024 267367
rect 4646 267261 4828 267295
rect 4572 267211 4584 267223
rect 4630 267211 4632 267222
rect 4831 267211 4844 267222
rect 4890 267211 4902 267223
rect 4572 266035 4632 267211
rect 4842 266035 4902 267211
rect 4572 266023 4584 266035
rect 4890 266023 4902 266035
rect 4646 265951 4828 265985
rect 4964 265949 5024 267297
rect 4976 265879 5024 265949
rect 4646 265843 4828 265877
rect 4572 265793 4584 265805
rect 4630 265793 4632 265804
rect 4831 265793 4844 265804
rect 4890 265793 4902 265805
rect 4572 264617 4632 265793
rect 4842 264617 4902 265793
rect 4572 264605 4584 264617
rect 4890 264605 4902 264617
rect 4646 264533 4828 264567
rect 4964 264531 5024 265879
rect 4976 264461 5024 264531
rect 4646 264425 4828 264459
rect 4572 264375 4584 264387
rect 4630 264375 4632 264386
rect 4831 264375 4844 264386
rect 4890 264375 4902 264387
rect 4572 263199 4632 264375
rect 4842 263199 4902 264375
rect 4572 263187 4584 263199
rect 4890 263187 4902 263199
rect 4646 263115 4828 263149
rect 4964 263113 5024 264461
rect 4976 263043 5024 263113
rect 4646 263007 4828 263041
rect 4572 262957 4584 262969
rect 4630 262957 4632 262968
rect 4831 262957 4844 262968
rect 4890 262957 4902 262969
rect 4572 261781 4632 262957
rect 4842 261781 4902 262957
rect 4572 261769 4584 261781
rect 4890 261769 4902 261781
rect 4646 261697 4828 261731
rect 4964 261695 5024 263043
rect 4976 261625 5024 261695
rect 4646 261589 4828 261623
rect 4572 261539 4584 261551
rect 4630 261539 4632 261550
rect 4831 261539 4844 261550
rect 4890 261539 4902 261551
rect 4572 260363 4632 261539
rect 4842 260363 4902 261539
rect 4572 260351 4584 260363
rect 4890 260351 4902 260363
rect 4646 260279 4828 260313
rect 4964 260277 5024 261625
rect 4976 260207 5024 260277
rect 4646 260171 4828 260205
rect 4572 260121 4584 260133
rect 4630 260121 4632 260132
rect 4831 260121 4844 260132
rect 4890 260121 4902 260133
rect 4572 258945 4632 260121
rect 4842 258945 4902 260121
rect 4572 258933 4584 258945
rect 4890 258933 4902 258945
rect 4646 258861 4828 258895
rect 4964 258859 5024 260207
rect 4976 258789 5024 258859
rect 4646 258753 4828 258787
rect 4572 258703 4584 258715
rect 4630 258703 4632 258714
rect 4831 258703 4844 258714
rect 4890 258703 4902 258715
rect 4572 257527 4632 258703
rect 4842 257527 4902 258703
rect 4572 257515 4584 257527
rect 4890 257515 4902 257527
rect 4646 257443 4828 257477
rect 4964 257441 5024 258789
rect 4976 257371 5024 257441
rect 4646 257335 4828 257369
rect 4572 257285 4584 257297
rect 4630 257285 4632 257296
rect 4831 257285 4844 257296
rect 4890 257285 4902 257297
rect 4572 256109 4632 257285
rect 4842 256109 4902 257285
rect 4572 256097 4584 256109
rect 4890 256097 4902 256109
rect 4646 256025 4828 256059
rect 4964 256023 5024 257371
rect 4976 255953 5024 256023
rect 4646 255917 4828 255951
rect 4572 255867 4584 255879
rect 4630 255867 4632 255878
rect 4831 255867 4844 255878
rect 4890 255867 4902 255879
rect 4572 254691 4632 255867
rect 4842 254691 4902 255867
rect 4572 254679 4584 254691
rect 4890 254679 4902 254691
rect 4646 254607 4828 254641
rect 4964 254605 5024 255953
rect 4976 254535 5024 254605
rect 4646 254499 4828 254533
rect 4572 254449 4584 254461
rect 4630 254449 4632 254460
rect 4831 254449 4844 254460
rect 4890 254449 4902 254461
rect 4572 253273 4632 254449
rect 4842 253273 4902 254449
rect 4572 253261 4584 253273
rect 4890 253261 4902 253273
rect 4646 253189 4828 253223
rect 4964 253187 5024 254535
rect 4976 253117 5024 253187
rect 4646 253081 4828 253115
rect 4572 253031 4584 253043
rect 4630 253031 4632 253042
rect 4831 253031 4844 253042
rect 4890 253031 4902 253043
rect 4572 251855 4632 253031
rect 4842 251855 4902 253031
rect 4572 251843 4584 251855
rect 4890 251843 4902 251855
rect 4646 251771 4828 251805
rect 4964 251769 5024 253117
rect 4976 251699 5024 251769
rect 4646 251663 4828 251697
rect 4572 251613 4584 251625
rect 4630 251613 4632 251624
rect 4831 251613 4844 251624
rect 4890 251613 4902 251625
rect 4572 250437 4632 251613
rect 4842 250437 4902 251613
rect 4572 250425 4584 250437
rect 4890 250425 4902 250437
rect 4646 250353 4828 250387
rect 4964 250351 5024 251699
rect 4976 250281 5024 250351
rect 4646 250245 4828 250279
rect 4572 250195 4584 250207
rect 4630 250195 4632 250206
rect 4831 250195 4844 250206
rect 4890 250195 4902 250207
rect 4572 249019 4632 250195
rect 4842 249019 4902 250195
rect 4572 249007 4584 249019
rect 4890 249007 4902 249019
rect 4646 248935 4828 248969
rect 4964 248933 5024 250281
rect 4976 248863 5024 248933
rect 4646 248827 4828 248861
rect 4572 248777 4584 248789
rect 4630 248777 4632 248788
rect 4831 248777 4844 248788
rect 4890 248777 4902 248789
rect 4572 247601 4632 248777
rect 4842 247601 4902 248777
rect 4572 247589 4584 247601
rect 4890 247589 4902 247601
rect 4646 247517 4828 247551
rect 4964 247515 5024 248863
rect 4976 247445 5024 247515
rect 4646 247409 4828 247443
rect 4572 247359 4584 247371
rect 4630 247359 4632 247370
rect 4831 247359 4844 247370
rect 4890 247359 4902 247371
rect 4572 246231 4632 247359
rect 4842 246231 4902 247359
rect 4964 246231 5024 247445
rect 5041 343844 5058 343940
rect 5137 343906 5519 343940
rect 5041 343804 5089 343844
rect 5567 343804 5615 343844
rect 5041 342456 5101 343804
rect 5237 343768 5419 343802
rect 5163 343718 5175 343730
rect 5221 343718 5223 343729
rect 5422 343718 5435 343729
rect 5481 343718 5493 343730
rect 5163 342542 5223 343718
rect 5433 342542 5493 343718
rect 5163 342530 5175 342542
rect 5481 342530 5493 342542
rect 5237 342458 5419 342492
rect 5555 342456 5615 343804
rect 5041 342386 5089 342456
rect 5567 342386 5615 342456
rect 5041 341038 5101 342386
rect 5237 342350 5419 342384
rect 5163 342300 5175 342312
rect 5221 342300 5223 342311
rect 5422 342300 5435 342311
rect 5481 342300 5493 342312
rect 5163 341124 5223 342300
rect 5433 341124 5493 342300
rect 5163 341112 5175 341124
rect 5481 341112 5493 341124
rect 5237 341040 5419 341074
rect 5555 341038 5615 342386
rect 5041 340968 5089 341038
rect 5567 340968 5615 341038
rect 5041 339620 5101 340968
rect 5237 340932 5419 340966
rect 5163 340882 5175 340894
rect 5221 340882 5223 340893
rect 5422 340882 5435 340893
rect 5481 340882 5493 340894
rect 5163 339706 5223 340882
rect 5433 339706 5493 340882
rect 5163 339694 5175 339706
rect 5481 339694 5493 339706
rect 5237 339622 5419 339656
rect 5555 339620 5615 340968
rect 5041 339550 5089 339620
rect 5567 339550 5615 339620
rect 5041 338202 5101 339550
rect 5237 339514 5419 339548
rect 5163 339464 5175 339476
rect 5221 339464 5223 339475
rect 5422 339464 5435 339475
rect 5481 339464 5493 339476
rect 5163 338288 5223 339464
rect 5433 338288 5493 339464
rect 5163 338276 5175 338288
rect 5481 338276 5493 338288
rect 5237 338204 5419 338238
rect 5555 338202 5615 339550
rect 5041 338132 5089 338202
rect 5567 338132 5615 338202
rect 5041 336784 5101 338132
rect 5237 338096 5419 338130
rect 5163 338046 5175 338058
rect 5221 338046 5223 338057
rect 5422 338046 5435 338057
rect 5481 338046 5493 338058
rect 5163 336870 5223 338046
rect 5433 336870 5493 338046
rect 5163 336858 5175 336870
rect 5481 336858 5493 336870
rect 5237 336786 5419 336820
rect 5555 336784 5615 338132
rect 5041 336714 5089 336784
rect 5567 336714 5615 336784
rect 5041 335366 5101 336714
rect 5237 336678 5419 336712
rect 5163 336628 5175 336640
rect 5221 336628 5223 336639
rect 5422 336628 5435 336639
rect 5481 336628 5493 336640
rect 5163 335452 5223 336628
rect 5433 335452 5493 336628
rect 5163 335440 5175 335452
rect 5481 335440 5493 335452
rect 5237 335368 5419 335402
rect 5555 335366 5615 336714
rect 5041 335296 5089 335366
rect 5567 335296 5615 335366
rect 5041 333948 5101 335296
rect 5237 335260 5419 335294
rect 5163 335210 5175 335222
rect 5221 335210 5223 335221
rect 5422 335210 5435 335221
rect 5481 335210 5493 335222
rect 5163 334034 5223 335210
rect 5433 334034 5493 335210
rect 5163 334022 5175 334034
rect 5481 334022 5493 334034
rect 5237 333950 5419 333984
rect 5555 333948 5615 335296
rect 5041 333878 5089 333948
rect 5567 333878 5615 333948
rect 5041 332530 5101 333878
rect 5237 333842 5419 333876
rect 5163 333792 5175 333804
rect 5221 333792 5223 333803
rect 5422 333792 5435 333803
rect 5481 333792 5493 333804
rect 5163 332616 5223 333792
rect 5433 332616 5493 333792
rect 5163 332604 5175 332616
rect 5481 332604 5493 332616
rect 5237 332532 5419 332566
rect 5555 332530 5615 333878
rect 5041 332460 5089 332530
rect 5567 332460 5615 332530
rect 5041 331112 5101 332460
rect 5237 332424 5419 332458
rect 5163 332374 5175 332386
rect 5221 332374 5223 332385
rect 5422 332374 5435 332385
rect 5481 332374 5493 332386
rect 5163 331198 5223 332374
rect 5433 331198 5493 332374
rect 5163 331186 5175 331198
rect 5481 331186 5493 331198
rect 5237 331114 5419 331148
rect 5555 331112 5615 332460
rect 5041 331042 5089 331112
rect 5567 331042 5615 331112
rect 5041 329694 5101 331042
rect 5237 331006 5419 331040
rect 5163 330956 5175 330968
rect 5221 330956 5223 330967
rect 5422 330956 5435 330967
rect 5481 330956 5493 330968
rect 5163 329780 5223 330956
rect 5433 329780 5493 330956
rect 5163 329768 5175 329780
rect 5481 329768 5493 329780
rect 5237 329696 5419 329730
rect 5555 329694 5615 331042
rect 5041 329624 5089 329694
rect 5567 329624 5615 329694
rect 5041 328276 5101 329624
rect 5237 329588 5419 329622
rect 5163 329538 5175 329550
rect 5221 329538 5223 329549
rect 5422 329538 5435 329549
rect 5481 329538 5493 329550
rect 5163 328362 5223 329538
rect 5433 328362 5493 329538
rect 5163 328350 5175 328362
rect 5481 328350 5493 328362
rect 5237 328278 5419 328312
rect 5555 328276 5615 329624
rect 5041 328206 5089 328276
rect 5567 328206 5615 328276
rect 5041 326858 5101 328206
rect 5237 328170 5419 328204
rect 5163 328120 5175 328132
rect 5221 328120 5223 328131
rect 5422 328120 5435 328131
rect 5481 328120 5493 328132
rect 5163 326944 5223 328120
rect 5433 326944 5493 328120
rect 5163 326932 5175 326944
rect 5481 326932 5493 326944
rect 5237 326860 5419 326894
rect 5555 326858 5615 328206
rect 5041 326788 5089 326858
rect 5567 326788 5615 326858
rect 5041 325440 5101 326788
rect 5237 326752 5419 326786
rect 5163 326702 5175 326714
rect 5221 326702 5223 326713
rect 5422 326702 5435 326713
rect 5481 326702 5493 326714
rect 5163 325526 5223 326702
rect 5433 325526 5493 326702
rect 5163 325514 5175 325526
rect 5481 325514 5493 325526
rect 5237 325442 5419 325476
rect 5555 325440 5615 326788
rect 5041 325370 5089 325440
rect 5567 325370 5615 325440
rect 5041 324022 5101 325370
rect 5237 325334 5419 325368
rect 5163 325284 5175 325296
rect 5221 325284 5223 325295
rect 5422 325284 5435 325295
rect 5481 325284 5493 325296
rect 5163 324108 5223 325284
rect 5433 324108 5493 325284
rect 5163 324096 5175 324108
rect 5481 324096 5493 324108
rect 5237 324024 5419 324058
rect 5555 324022 5615 325370
rect 5041 323952 5089 324022
rect 5567 323952 5615 324022
rect 5041 322604 5101 323952
rect 5237 323916 5419 323950
rect 5163 323866 5175 323878
rect 5221 323866 5223 323877
rect 5422 323866 5435 323877
rect 5481 323866 5493 323878
rect 5163 322690 5223 323866
rect 5433 322690 5493 323866
rect 5163 322678 5175 322690
rect 5481 322678 5493 322690
rect 5237 322606 5419 322640
rect 5555 322604 5615 323952
rect 5041 322534 5089 322604
rect 5567 322534 5615 322604
rect 5041 321186 5101 322534
rect 5237 322498 5419 322532
rect 5163 322448 5175 322460
rect 5221 322448 5223 322459
rect 5422 322448 5435 322459
rect 5481 322448 5493 322460
rect 5163 321272 5223 322448
rect 5433 321272 5493 322448
rect 5163 321260 5175 321272
rect 5481 321260 5493 321272
rect 5237 321188 5419 321222
rect 5555 321186 5615 322534
rect 5041 321116 5089 321186
rect 5567 321116 5615 321186
rect 5041 319768 5101 321116
rect 5237 321080 5419 321114
rect 5163 321030 5175 321042
rect 5221 321030 5223 321041
rect 5422 321030 5435 321041
rect 5481 321030 5493 321042
rect 5163 319854 5223 321030
rect 5433 319854 5493 321030
rect 5163 319842 5175 319854
rect 5481 319842 5493 319854
rect 5237 319770 5419 319804
rect 5555 319768 5615 321116
rect 5041 319698 5089 319768
rect 5567 319698 5615 319768
rect 5041 318350 5101 319698
rect 5237 319662 5419 319696
rect 5163 319612 5175 319624
rect 5221 319612 5223 319623
rect 5422 319612 5435 319623
rect 5481 319612 5493 319624
rect 5163 318436 5223 319612
rect 5433 318436 5493 319612
rect 5163 318424 5175 318436
rect 5481 318424 5493 318436
rect 5237 318352 5419 318386
rect 5555 318350 5615 319698
rect 5041 318280 5089 318350
rect 5567 318280 5615 318350
rect 5041 316932 5101 318280
rect 5237 318244 5419 318278
rect 5163 318194 5175 318206
rect 5221 318194 5223 318205
rect 5422 318194 5435 318205
rect 5481 318194 5493 318206
rect 5163 317018 5223 318194
rect 5433 317018 5493 318194
rect 5163 317006 5175 317018
rect 5481 317006 5493 317018
rect 5237 316934 5419 316968
rect 5555 316932 5615 318280
rect 5041 316862 5089 316932
rect 5567 316862 5615 316932
rect 5041 315514 5101 316862
rect 5237 316826 5419 316860
rect 5163 316776 5175 316788
rect 5221 316776 5223 316787
rect 5422 316776 5435 316787
rect 5481 316776 5493 316788
rect 5163 315600 5223 316776
rect 5433 315600 5493 316776
rect 5163 315588 5175 315600
rect 5481 315588 5493 315600
rect 5237 315516 5419 315550
rect 5555 315514 5615 316862
rect 5041 315444 5089 315514
rect 5567 315444 5615 315514
rect 5041 314096 5101 315444
rect 5237 315408 5419 315442
rect 5163 315358 5175 315370
rect 5221 315358 5223 315369
rect 5422 315358 5435 315369
rect 5481 315358 5493 315370
rect 5163 314182 5223 315358
rect 5433 314182 5493 315358
rect 5163 314170 5175 314182
rect 5481 314170 5493 314182
rect 5237 314098 5419 314132
rect 5555 314096 5615 315444
rect 5041 314026 5089 314096
rect 5567 314026 5615 314096
rect 5041 312678 5101 314026
rect 5237 313990 5419 314024
rect 5163 313940 5175 313952
rect 5221 313940 5223 313951
rect 5422 313940 5435 313951
rect 5481 313940 5493 313952
rect 5163 312764 5223 313940
rect 5433 312764 5493 313940
rect 5163 312752 5175 312764
rect 5481 312752 5493 312764
rect 5237 312680 5419 312714
rect 5555 312678 5615 314026
rect 5041 312608 5089 312678
rect 5567 312608 5615 312678
rect 5041 311260 5101 312608
rect 5237 312572 5419 312606
rect 5163 312522 5175 312534
rect 5221 312522 5223 312533
rect 5422 312522 5435 312533
rect 5481 312522 5493 312534
rect 5163 311346 5223 312522
rect 5433 311346 5493 312522
rect 5163 311334 5175 311346
rect 5481 311334 5493 311346
rect 5237 311262 5419 311296
rect 5555 311260 5615 312608
rect 5041 311190 5089 311260
rect 5567 311190 5615 311260
rect 5041 309842 5101 311190
rect 5237 311154 5419 311188
rect 5163 311104 5175 311116
rect 5221 311104 5223 311115
rect 5422 311104 5435 311115
rect 5481 311104 5493 311116
rect 5163 309928 5223 311104
rect 5433 309928 5493 311104
rect 5163 309916 5175 309928
rect 5481 309916 5493 309928
rect 5237 309844 5419 309878
rect 5555 309842 5615 311190
rect 5041 309772 5089 309842
rect 5567 309772 5615 309842
rect 5041 308424 5101 309772
rect 5237 309736 5419 309770
rect 5163 309686 5175 309698
rect 5221 309686 5223 309697
rect 5422 309686 5435 309697
rect 5481 309686 5493 309698
rect 5163 308510 5223 309686
rect 5433 308510 5493 309686
rect 5163 308498 5175 308510
rect 5481 308498 5493 308510
rect 5237 308426 5419 308460
rect 5555 308424 5615 309772
rect 5041 308354 5089 308424
rect 5567 308354 5615 308424
rect 5041 307006 5101 308354
rect 5237 308318 5419 308352
rect 5163 308268 5175 308280
rect 5221 308268 5223 308279
rect 5422 308268 5435 308279
rect 5481 308268 5493 308280
rect 5163 307092 5223 308268
rect 5433 307092 5493 308268
rect 5163 307080 5175 307092
rect 5481 307080 5493 307092
rect 5237 307008 5419 307042
rect 5555 307006 5615 308354
rect 5041 306936 5089 307006
rect 5567 306936 5615 307006
rect 5041 305588 5101 306936
rect 5237 306900 5419 306934
rect 5163 306850 5175 306862
rect 5221 306850 5223 306861
rect 5422 306850 5435 306861
rect 5481 306850 5493 306862
rect 5163 305674 5223 306850
rect 5433 305674 5493 306850
rect 5163 305662 5175 305674
rect 5481 305662 5493 305674
rect 5237 305590 5419 305624
rect 5555 305588 5615 306936
rect 5041 305518 5089 305588
rect 5567 305518 5615 305588
rect 5041 304170 5101 305518
rect 5237 305482 5419 305516
rect 5163 305432 5175 305444
rect 5221 305432 5223 305443
rect 5422 305432 5435 305443
rect 5481 305432 5493 305444
rect 5163 304256 5223 305432
rect 5433 304256 5493 305432
rect 5163 304244 5175 304256
rect 5481 304244 5493 304256
rect 5237 304172 5419 304206
rect 5555 304170 5615 305518
rect 5041 304100 5089 304170
rect 5567 304100 5615 304170
rect 5041 302752 5101 304100
rect 5237 304064 5419 304098
rect 5163 304014 5175 304026
rect 5221 304014 5223 304025
rect 5422 304014 5435 304025
rect 5481 304014 5493 304026
rect 5163 302838 5223 304014
rect 5433 302838 5493 304014
rect 5163 302826 5175 302838
rect 5481 302826 5493 302838
rect 5237 302754 5419 302788
rect 5555 302752 5615 304100
rect 5041 302682 5089 302752
rect 5567 302682 5615 302752
rect 5041 301334 5101 302682
rect 5237 302646 5419 302680
rect 5163 302596 5175 302608
rect 5221 302596 5223 302607
rect 5422 302596 5435 302607
rect 5481 302596 5493 302608
rect 5163 301420 5223 302596
rect 5433 301420 5493 302596
rect 5163 301408 5175 301420
rect 5481 301408 5493 301420
rect 5237 301336 5419 301370
rect 5555 301334 5615 302682
rect 5041 301264 5089 301334
rect 5567 301264 5615 301334
rect 5041 299916 5101 301264
rect 5237 301228 5419 301262
rect 5163 301178 5175 301190
rect 5221 301178 5223 301189
rect 5422 301178 5435 301189
rect 5481 301178 5493 301190
rect 5163 300002 5223 301178
rect 5433 300002 5493 301178
rect 5163 299990 5175 300002
rect 5481 299990 5493 300002
rect 5237 299918 5419 299952
rect 5555 299916 5615 301264
rect 5041 299846 5089 299916
rect 5567 299846 5615 299916
rect 5041 298498 5101 299846
rect 5237 299810 5419 299844
rect 5163 299760 5175 299772
rect 5221 299760 5223 299771
rect 5422 299760 5435 299771
rect 5481 299760 5493 299772
rect 5163 298584 5223 299760
rect 5433 298584 5493 299760
rect 5163 298572 5175 298584
rect 5481 298572 5493 298584
rect 5237 298500 5419 298534
rect 5555 298498 5615 299846
rect 5041 298428 5089 298498
rect 5567 298428 5615 298498
rect 5041 297080 5101 298428
rect 5237 298392 5419 298426
rect 5163 298342 5175 298354
rect 5221 298342 5223 298353
rect 5422 298342 5435 298353
rect 5481 298342 5493 298354
rect 5163 297166 5223 298342
rect 5433 297166 5493 298342
rect 5163 297154 5175 297166
rect 5481 297154 5493 297166
rect 5237 297082 5419 297116
rect 5555 297080 5615 298428
rect 5041 297010 5089 297080
rect 5567 297010 5615 297080
rect 5041 295662 5101 297010
rect 5237 296974 5419 297008
rect 5163 296924 5175 296936
rect 5221 296924 5223 296935
rect 5422 296924 5435 296935
rect 5481 296924 5493 296936
rect 5163 295748 5223 296924
rect 5433 295748 5493 296924
rect 5163 295736 5175 295748
rect 5481 295736 5493 295748
rect 5237 295664 5419 295698
rect 5555 295662 5615 297010
rect 5041 295592 5089 295662
rect 5567 295592 5615 295662
rect 5041 294244 5101 295592
rect 5237 295556 5419 295590
rect 5163 295506 5175 295518
rect 5221 295506 5223 295517
rect 5422 295506 5435 295517
rect 5481 295506 5493 295518
rect 5163 294330 5223 295506
rect 5433 294330 5493 295506
rect 5163 294318 5175 294330
rect 5481 294318 5493 294330
rect 5237 294246 5419 294280
rect 5555 294244 5615 295592
rect 5041 294174 5089 294244
rect 5567 294174 5615 294244
rect 5041 292826 5101 294174
rect 5237 294138 5419 294172
rect 5163 294088 5175 294100
rect 5221 294088 5223 294099
rect 5422 294088 5435 294099
rect 5481 294088 5493 294100
rect 5163 292912 5223 294088
rect 5433 292912 5493 294088
rect 5163 292900 5175 292912
rect 5481 292900 5493 292912
rect 5237 292828 5419 292862
rect 5555 292826 5615 294174
rect 5041 292756 5089 292826
rect 5567 292756 5615 292826
rect 5041 291408 5101 292756
rect 5237 292720 5419 292754
rect 5163 292670 5175 292682
rect 5221 292670 5223 292681
rect 5422 292670 5435 292681
rect 5481 292670 5493 292682
rect 5163 291494 5223 292670
rect 5433 291494 5493 292670
rect 5163 291482 5175 291494
rect 5481 291482 5493 291494
rect 5237 291410 5419 291444
rect 5555 291408 5615 292756
rect 5041 291338 5089 291408
rect 5567 291338 5615 291408
rect 5041 289990 5101 291338
rect 5237 291302 5419 291336
rect 5163 291252 5175 291264
rect 5221 291252 5223 291263
rect 5422 291252 5435 291263
rect 5481 291252 5493 291264
rect 5163 290076 5223 291252
rect 5433 290076 5493 291252
rect 5163 290064 5175 290076
rect 5481 290064 5493 290076
rect 5237 289992 5419 290026
rect 5555 289990 5615 291338
rect 5041 289920 5089 289990
rect 5567 289920 5615 289990
rect 5041 288572 5101 289920
rect 5237 289884 5419 289918
rect 5163 289834 5175 289846
rect 5221 289834 5223 289845
rect 5422 289834 5435 289845
rect 5481 289834 5493 289846
rect 5163 288658 5223 289834
rect 5433 288658 5493 289834
rect 5163 288646 5175 288658
rect 5481 288646 5493 288658
rect 5237 288574 5419 288608
rect 5555 288572 5615 289920
rect 5041 288502 5089 288572
rect 5567 288502 5615 288572
rect 5041 287154 5101 288502
rect 5237 288466 5419 288500
rect 5163 288416 5175 288428
rect 5221 288416 5223 288427
rect 5422 288416 5435 288427
rect 5481 288416 5493 288428
rect 5163 287240 5223 288416
rect 5433 287240 5493 288416
rect 5163 287228 5175 287240
rect 5481 287228 5493 287240
rect 5237 287156 5419 287190
rect 5555 287154 5615 288502
rect 5041 287084 5089 287154
rect 5567 287084 5615 287154
rect 5041 285736 5101 287084
rect 5237 287048 5419 287082
rect 5163 286998 5175 287010
rect 5221 286998 5223 287009
rect 5422 286998 5435 287009
rect 5481 286998 5493 287010
rect 5163 285822 5223 286998
rect 5433 285822 5493 286998
rect 5163 285810 5175 285822
rect 5481 285810 5493 285822
rect 5237 285738 5419 285772
rect 5555 285736 5615 287084
rect 5041 285666 5089 285736
rect 5567 285666 5615 285736
rect 5041 284318 5101 285666
rect 5237 285630 5419 285664
rect 5163 285580 5175 285592
rect 5221 285580 5223 285591
rect 5422 285580 5435 285591
rect 5481 285580 5493 285592
rect 5163 284404 5223 285580
rect 5433 284404 5493 285580
rect 5163 284392 5175 284404
rect 5481 284392 5493 284404
rect 5237 284320 5419 284354
rect 5555 284318 5615 285666
rect 5041 284248 5089 284318
rect 5567 284248 5615 284318
rect 5041 282900 5101 284248
rect 5237 284212 5419 284246
rect 5163 284162 5175 284174
rect 5221 284162 5223 284173
rect 5422 284162 5435 284173
rect 5481 284162 5493 284174
rect 5163 282986 5223 284162
rect 5433 282986 5493 284162
rect 5163 282974 5175 282986
rect 5481 282974 5493 282986
rect 5237 282902 5419 282936
rect 5555 282900 5615 284248
rect 5041 282830 5089 282900
rect 5567 282830 5615 282900
rect 5041 281482 5101 282830
rect 5237 282794 5419 282828
rect 5163 282744 5175 282756
rect 5221 282744 5223 282755
rect 5422 282744 5435 282755
rect 5481 282744 5493 282756
rect 5163 281568 5223 282744
rect 5433 281568 5493 282744
rect 5163 281556 5175 281568
rect 5481 281556 5493 281568
rect 5237 281484 5419 281518
rect 5555 281482 5615 282830
rect 5041 281412 5089 281482
rect 5567 281412 5615 281482
rect 5041 280064 5101 281412
rect 5237 281376 5419 281410
rect 5163 281326 5175 281338
rect 5221 281326 5223 281337
rect 5422 281326 5435 281337
rect 5481 281326 5493 281338
rect 5163 280150 5223 281326
rect 5433 280150 5493 281326
rect 5163 280138 5175 280150
rect 5481 280138 5493 280150
rect 5237 280066 5419 280100
rect 5555 280064 5615 281412
rect 5041 279994 5089 280064
rect 5567 279994 5615 280064
rect 5041 278646 5101 279994
rect 5237 279958 5419 279992
rect 5163 279908 5175 279920
rect 5221 279908 5223 279919
rect 5422 279908 5435 279919
rect 5481 279908 5493 279920
rect 5163 278732 5223 279908
rect 5433 278732 5493 279908
rect 5163 278720 5175 278732
rect 5481 278720 5493 278732
rect 5237 278648 5419 278682
rect 5555 278646 5615 279994
rect 5041 278576 5089 278646
rect 5567 278576 5615 278646
rect 5041 277228 5101 278576
rect 5237 278540 5419 278574
rect 5163 278490 5175 278502
rect 5221 278490 5223 278501
rect 5422 278490 5435 278501
rect 5481 278490 5493 278502
rect 5163 277314 5223 278490
rect 5433 277314 5493 278490
rect 5163 277302 5175 277314
rect 5481 277302 5493 277314
rect 5237 277230 5419 277264
rect 5555 277228 5615 278576
rect 5041 277158 5089 277228
rect 5567 277158 5615 277228
rect 5041 275810 5101 277158
rect 5237 277122 5419 277156
rect 5163 277072 5175 277084
rect 5221 277072 5223 277083
rect 5422 277072 5435 277083
rect 5481 277072 5493 277084
rect 5163 275896 5223 277072
rect 5433 275896 5493 277072
rect 5163 275884 5175 275896
rect 5481 275884 5493 275896
rect 5237 275812 5419 275846
rect 5555 275810 5615 277158
rect 5041 275740 5089 275810
rect 5567 275740 5615 275810
rect 5041 274392 5101 275740
rect 5237 275704 5419 275738
rect 5163 275654 5175 275666
rect 5221 275654 5223 275665
rect 5422 275654 5435 275665
rect 5481 275654 5493 275666
rect 5163 274478 5223 275654
rect 5433 274478 5493 275654
rect 5163 274466 5175 274478
rect 5481 274466 5493 274478
rect 5237 274394 5419 274428
rect 5555 274392 5615 275740
rect 5041 274322 5089 274392
rect 5567 274322 5615 274392
rect 5041 272974 5101 274322
rect 5237 274286 5419 274320
rect 5163 274236 5175 274248
rect 5221 274236 5223 274247
rect 5422 274236 5435 274247
rect 5481 274236 5493 274248
rect 5163 273060 5223 274236
rect 5433 273060 5493 274236
rect 5163 273048 5175 273060
rect 5481 273048 5493 273060
rect 5237 272976 5419 273010
rect 5555 272974 5615 274322
rect 5041 272904 5089 272974
rect 5567 272904 5615 272974
rect 5041 271556 5101 272904
rect 5237 272868 5419 272902
rect 5163 272818 5175 272830
rect 5221 272818 5223 272829
rect 5422 272818 5435 272829
rect 5481 272818 5493 272830
rect 5163 271642 5223 272818
rect 5433 271642 5493 272818
rect 5163 271630 5175 271642
rect 5481 271630 5493 271642
rect 5237 271558 5419 271592
rect 5555 271556 5615 272904
rect 5041 271486 5089 271556
rect 5567 271486 5615 271556
rect 5041 270138 5101 271486
rect 5237 271450 5419 271484
rect 5163 271400 5175 271412
rect 5221 271400 5223 271411
rect 5422 271400 5435 271411
rect 5481 271400 5493 271412
rect 5163 270224 5223 271400
rect 5433 270224 5493 271400
rect 5163 270212 5175 270224
rect 5481 270212 5493 270224
rect 5237 270140 5419 270174
rect 5555 270138 5615 271486
rect 5041 270068 5089 270138
rect 5567 270068 5615 270138
rect 5041 268720 5101 270068
rect 5237 270032 5419 270066
rect 5163 269982 5175 269994
rect 5221 269982 5223 269993
rect 5422 269982 5435 269993
rect 5481 269982 5493 269994
rect 5163 268806 5223 269982
rect 5433 268806 5493 269982
rect 5163 268794 5175 268806
rect 5481 268794 5493 268806
rect 5237 268722 5419 268756
rect 5555 268720 5615 270068
rect 5041 268650 5089 268720
rect 5567 268650 5615 268720
rect 5041 267302 5101 268650
rect 5237 268614 5419 268648
rect 5163 268564 5175 268576
rect 5221 268564 5223 268575
rect 5422 268564 5435 268575
rect 5481 268564 5493 268576
rect 5163 267388 5223 268564
rect 5433 267388 5493 268564
rect 5163 267376 5175 267388
rect 5481 267376 5493 267388
rect 5237 267304 5419 267338
rect 5555 267302 5615 268650
rect 5041 267232 5089 267302
rect 5567 267232 5615 267302
rect 5041 265884 5101 267232
rect 5237 267196 5419 267230
rect 5163 267146 5175 267158
rect 5221 267146 5223 267157
rect 5422 267146 5435 267157
rect 5481 267146 5493 267158
rect 5163 265970 5223 267146
rect 5433 265970 5493 267146
rect 5163 265958 5175 265970
rect 5481 265958 5493 265970
rect 5237 265886 5419 265920
rect 5555 265884 5615 267232
rect 5041 265814 5089 265884
rect 5567 265814 5615 265884
rect 5041 264466 5101 265814
rect 5237 265778 5419 265812
rect 5163 265728 5175 265740
rect 5221 265728 5223 265739
rect 5422 265728 5435 265739
rect 5481 265728 5493 265740
rect 5163 264552 5223 265728
rect 5433 264552 5493 265728
rect 5163 264540 5175 264552
rect 5481 264540 5493 264552
rect 5237 264468 5419 264502
rect 5555 264466 5615 265814
rect 5041 264396 5089 264466
rect 5567 264396 5615 264466
rect 5041 263048 5101 264396
rect 5237 264360 5419 264394
rect 5163 264310 5175 264322
rect 5221 264310 5223 264321
rect 5422 264310 5435 264321
rect 5481 264310 5493 264322
rect 5163 263134 5223 264310
rect 5433 263134 5493 264310
rect 5163 263122 5175 263134
rect 5481 263122 5493 263134
rect 5237 263050 5419 263084
rect 5555 263048 5615 264396
rect 5041 262978 5089 263048
rect 5567 262978 5615 263048
rect 5041 261630 5101 262978
rect 5237 262942 5419 262976
rect 5163 262892 5175 262904
rect 5221 262892 5223 262903
rect 5422 262892 5435 262903
rect 5481 262892 5493 262904
rect 5163 261716 5223 262892
rect 5433 261716 5493 262892
rect 5163 261704 5175 261716
rect 5481 261704 5493 261716
rect 5237 261632 5419 261666
rect 5555 261630 5615 262978
rect 5041 261560 5089 261630
rect 5567 261560 5615 261630
rect 5041 260212 5101 261560
rect 5237 261524 5419 261558
rect 5163 261474 5175 261486
rect 5221 261474 5223 261485
rect 5422 261474 5435 261485
rect 5481 261474 5493 261486
rect 5163 260298 5223 261474
rect 5433 260298 5493 261474
rect 5163 260286 5175 260298
rect 5481 260286 5493 260298
rect 5237 260214 5419 260248
rect 5555 260212 5615 261560
rect 5041 260142 5089 260212
rect 5567 260142 5615 260212
rect 5041 258794 5101 260142
rect 5237 260106 5419 260140
rect 5163 260056 5175 260068
rect 5221 260056 5223 260067
rect 5422 260056 5435 260067
rect 5481 260056 5493 260068
rect 5163 258880 5223 260056
rect 5433 258880 5493 260056
rect 5163 258868 5175 258880
rect 5481 258868 5493 258880
rect 5237 258796 5419 258830
rect 5555 258794 5615 260142
rect 5041 258724 5089 258794
rect 5567 258724 5615 258794
rect 5041 257376 5101 258724
rect 5237 258688 5419 258722
rect 5163 258638 5175 258650
rect 5221 258638 5223 258649
rect 5422 258638 5435 258649
rect 5481 258638 5493 258650
rect 5163 257462 5223 258638
rect 5433 257462 5493 258638
rect 5163 257450 5175 257462
rect 5481 257450 5493 257462
rect 5237 257378 5419 257412
rect 5555 257376 5615 258724
rect 5041 257306 5089 257376
rect 5567 257306 5615 257376
rect 5041 255958 5101 257306
rect 5237 257270 5419 257304
rect 5163 257220 5175 257232
rect 5221 257220 5223 257231
rect 5422 257220 5435 257231
rect 5481 257220 5493 257232
rect 5163 256044 5223 257220
rect 5433 256044 5493 257220
rect 5163 256032 5175 256044
rect 5481 256032 5493 256044
rect 5237 255960 5419 255994
rect 5555 255958 5615 257306
rect 5041 255888 5089 255958
rect 5567 255888 5615 255958
rect 5041 254540 5101 255888
rect 5237 255852 5419 255886
rect 5163 255802 5175 255814
rect 5221 255802 5223 255813
rect 5422 255802 5435 255813
rect 5481 255802 5493 255814
rect 5163 254626 5223 255802
rect 5433 254626 5493 255802
rect 5163 254614 5175 254626
rect 5481 254614 5493 254626
rect 5237 254542 5419 254576
rect 5555 254540 5615 255888
rect 5041 254470 5089 254540
rect 5567 254470 5615 254540
rect 5041 253122 5101 254470
rect 5237 254434 5419 254468
rect 5163 254384 5175 254396
rect 5221 254384 5223 254395
rect 5422 254384 5435 254395
rect 5481 254384 5493 254396
rect 5163 253208 5223 254384
rect 5433 253208 5493 254384
rect 5163 253196 5175 253208
rect 5481 253196 5493 253208
rect 5237 253124 5419 253158
rect 5555 253122 5615 254470
rect 5041 253052 5089 253122
rect 5567 253052 5615 253122
rect 5041 251704 5101 253052
rect 5237 253016 5419 253050
rect 5163 252966 5175 252978
rect 5221 252966 5223 252977
rect 5422 252966 5435 252977
rect 5481 252966 5493 252978
rect 5163 251790 5223 252966
rect 5433 251790 5493 252966
rect 5163 251778 5175 251790
rect 5481 251778 5493 251790
rect 5237 251706 5419 251740
rect 5555 251704 5615 253052
rect 5041 251634 5089 251704
rect 5567 251634 5615 251704
rect 5041 250286 5101 251634
rect 5237 251598 5419 251632
rect 5163 251548 5175 251560
rect 5221 251548 5223 251559
rect 5422 251548 5435 251559
rect 5481 251548 5493 251560
rect 5163 250372 5223 251548
rect 5433 250372 5493 251548
rect 5163 250360 5175 250372
rect 5481 250360 5493 250372
rect 5237 250288 5419 250322
rect 5555 250286 5615 251634
rect 5041 250216 5089 250286
rect 5567 250216 5615 250286
rect 5041 248868 5101 250216
rect 5237 250180 5419 250214
rect 5163 250130 5175 250142
rect 5221 250130 5223 250141
rect 5422 250130 5435 250141
rect 5481 250130 5493 250142
rect 5163 248954 5223 250130
rect 5433 248954 5493 250130
rect 5163 248942 5175 248954
rect 5481 248942 5493 248954
rect 5237 248870 5419 248904
rect 5555 248868 5615 250216
rect 5041 248798 5089 248868
rect 5567 248798 5615 248868
rect 5041 247450 5101 248798
rect 5237 248762 5419 248796
rect 5163 248712 5175 248724
rect 5221 248712 5223 248723
rect 5422 248712 5435 248723
rect 5481 248712 5493 248724
rect 5163 247536 5223 248712
rect 5433 247536 5493 248712
rect 5163 247524 5175 247536
rect 5481 247524 5493 247536
rect 5237 247452 5419 247486
rect 5555 247450 5615 248798
rect 5041 247380 5089 247450
rect 5567 247380 5615 247450
rect 5041 246231 5101 247380
rect 5237 247344 5419 247378
rect 5163 247294 5175 247306
rect 5221 247294 5223 247305
rect 5422 247294 5435 247305
rect 5481 247294 5493 247306
rect 5163 246231 5223 247294
rect 3795 246136 5223 246231
rect 5433 246136 5493 247294
rect 5555 246136 5615 247380
rect 3795 246012 5663 246136
rect 3465 245287 3647 245321
rect 3465 245179 3647 245213
rect 3449 245120 3451 245131
rect 3650 245120 3663 245131
rect 3403 243944 3451 245120
rect 3661 243944 3709 245120
rect 3465 243851 3647 243885
rect 3465 243743 3647 243777
rect 3449 243684 3451 243695
rect 3650 243684 3663 243695
rect 3403 242508 3451 243684
rect 3661 242508 3709 243684
rect 3465 242415 3647 242449
rect 3465 242307 3647 242341
rect 3449 242248 3451 242259
rect 3650 242248 3663 242259
rect 3403 241072 3451 242248
rect 3661 241072 3709 242248
rect 3465 240979 3647 241013
rect 3465 240871 3647 240905
rect 3449 240812 3451 240823
rect 3650 240812 3663 240823
rect 3403 239636 3451 240812
rect 3661 239636 3709 240812
rect 3465 239543 3647 239577
rect 3465 239435 3647 239469
rect 3449 239376 3451 239387
rect 3650 239376 3663 239387
rect 3403 238200 3451 239376
rect 3661 238200 3709 239376
rect 3465 238107 3647 238141
rect 3465 237999 3647 238033
rect 3449 237940 3451 237951
rect 3650 237940 3663 237951
rect 3403 236764 3451 237940
rect 3661 236764 3709 237940
rect 3465 236671 3647 236705
rect 3465 236563 3647 236597
rect 3449 236504 3451 236515
rect 3650 236504 3663 236515
rect 3403 235328 3451 236504
rect 3661 235328 3709 236504
rect 3465 235235 3647 235269
rect 3465 235127 3647 235161
rect 3449 235068 3451 235079
rect 3650 235068 3663 235079
rect 3403 233892 3451 235068
rect 3661 233892 3709 235068
rect 3465 233799 3647 233833
rect 3465 233691 3647 233725
rect 3449 233632 3451 233643
rect 3650 233632 3663 233643
rect 3403 232456 3451 233632
rect 3661 232456 3709 233632
rect 3465 232363 3647 232397
rect 3465 232255 3647 232289
rect 3449 232196 3451 232207
rect 3650 232196 3663 232207
rect 3403 231020 3451 232196
rect 3661 231020 3709 232196
rect 3465 230927 3647 230961
rect 3465 230819 3647 230853
rect 3449 230760 3451 230771
rect 3650 230760 3663 230771
rect 3403 229584 3451 230760
rect 3661 229584 3709 230760
rect 3465 229491 3647 229525
rect 3465 229383 3647 229417
rect 3449 229324 3451 229335
rect 3650 229324 3663 229335
rect 3403 228148 3451 229324
rect 3661 228148 3709 229324
rect 3465 228055 3647 228089
rect 3465 227947 3647 227981
rect 3449 227888 3451 227899
rect 3650 227888 3663 227899
rect 3403 226712 3451 227888
rect 3661 226712 3709 227888
rect 3465 226619 3647 226653
rect 3465 226511 3647 226545
rect 3449 226452 3451 226463
rect 3650 226452 3663 226463
rect 3403 225276 3451 226452
rect 3661 225276 3709 226452
rect 3465 225183 3647 225217
rect 3465 225075 3647 225109
rect 3449 225016 3451 225027
rect 3650 225016 3663 225027
rect 3403 223840 3451 225016
rect 3661 223840 3709 225016
rect 3465 223747 3647 223781
rect 3465 223639 3647 223673
rect 3449 223580 3451 223591
rect 3650 223580 3663 223591
rect 3403 222404 3451 223580
rect 3661 222404 3709 223580
rect 3465 222311 3647 222345
rect 3465 222203 3647 222237
rect 3449 222144 3451 222155
rect 3650 222144 3663 222155
rect 3403 220968 3451 222144
rect 3661 220968 3709 222144
rect 3465 220875 3647 220909
rect 3465 220767 3647 220801
rect 3449 220708 3451 220719
rect 3650 220708 3663 220719
rect 3403 219532 3451 220708
rect 3661 219532 3709 220708
rect 3465 219439 3647 219473
rect 3465 219331 3647 219365
rect 3449 219272 3451 219283
rect 3650 219272 3663 219283
rect 3403 218096 3451 219272
rect 3661 218096 3709 219272
rect 3465 218003 3647 218037
rect 3465 217895 3647 217929
rect 3449 217836 3451 217847
rect 3650 217836 3663 217847
rect 3403 216660 3451 217836
rect 3661 216660 3709 217836
rect 3465 216567 3647 216601
rect 3465 216459 3647 216493
rect 3449 216400 3451 216411
rect 3650 216400 3663 216411
rect 3403 215224 3451 216400
rect 3661 215224 3709 216400
rect 3465 215131 3647 215165
rect 3465 215023 3647 215057
rect 3449 214964 3451 214975
rect 3650 214964 3663 214975
rect 3403 213788 3451 214964
rect 3661 213788 3709 214964
rect 3465 213695 3647 213729
rect 3465 213587 3647 213621
rect 3449 213528 3451 213539
rect 3650 213528 3663 213539
rect 3403 212352 3451 213528
rect 3661 212352 3709 213528
rect 3465 212259 3647 212293
rect 3465 212151 3647 212185
rect 3449 212092 3451 212103
rect 3650 212092 3663 212103
rect 3403 210916 3451 212092
rect 3661 210916 3709 212092
rect 3465 210823 3647 210857
rect 3465 210715 3647 210749
rect 3449 210656 3451 210667
rect 3650 210656 3663 210667
rect 3403 209480 3451 210656
rect 3661 209480 3709 210656
rect 3465 209387 3647 209421
rect 3465 209279 3647 209313
rect 3449 209220 3451 209231
rect 3650 209220 3663 209231
rect 3403 208044 3451 209220
rect 3661 208044 3709 209220
rect 3465 207951 3647 207985
rect 3465 207843 3647 207877
rect 3449 207784 3451 207795
rect 3650 207784 3663 207795
rect 3403 206608 3451 207784
rect 3661 206608 3709 207784
rect 3465 206515 3647 206549
rect 3465 206407 3647 206441
rect 3449 206348 3451 206359
rect 3650 206348 3663 206359
rect 3403 205172 3451 206348
rect 3661 205172 3709 206348
rect 3465 205079 3647 205113
rect 3465 204971 3647 205005
rect 3449 204912 3451 204923
rect 3650 204912 3663 204923
rect 3403 203736 3451 204912
rect 3661 203736 3709 204912
rect 3465 203643 3647 203677
rect 3465 203535 3647 203569
rect 3449 203476 3451 203487
rect 3650 203476 3663 203487
rect 3403 202300 3451 203476
rect 3661 202300 3709 203476
rect 3465 202207 3647 202241
rect 3465 202099 3647 202133
rect 3449 202040 3451 202051
rect 3650 202040 3663 202051
rect 3403 200864 3451 202040
rect 3661 200864 3709 202040
rect 3465 200771 3647 200805
rect 3465 200663 3647 200697
rect 3449 200604 3451 200615
rect 3650 200604 3663 200615
rect 3403 199428 3451 200604
rect 3661 199428 3709 200604
rect 3465 199335 3647 199369
rect 3465 199227 3647 199261
rect 3449 199168 3451 199179
rect 3650 199168 3663 199179
rect 3403 197992 3451 199168
rect 3661 197992 3709 199168
rect 3465 197899 3647 197933
rect 3465 197791 3647 197825
rect 3449 197732 3451 197743
rect 3650 197732 3663 197743
rect 3403 196556 3451 197732
rect 3661 196556 3709 197732
rect 3465 196463 3647 196497
rect 3465 196355 3647 196389
rect 3449 196296 3451 196307
rect 3650 196296 3663 196307
rect 3403 195120 3451 196296
rect 3661 195120 3709 196296
rect 3465 195027 3647 195061
rect 3465 194919 3647 194953
rect 3449 194860 3451 194871
rect 3650 194860 3663 194871
rect 3403 193684 3451 194860
rect 3661 193684 3709 194860
rect 3465 193591 3647 193625
rect 3465 193483 3647 193517
rect 3449 193424 3451 193435
rect 3650 193424 3663 193435
rect 3403 192248 3451 193424
rect 3661 192248 3709 193424
rect 3465 192155 3647 192189
rect 3465 192047 3647 192081
rect 3449 191988 3451 191999
rect 3650 191988 3663 191999
rect 3403 190812 3451 191988
rect 3661 190812 3709 191988
rect 3465 190719 3647 190753
rect 3465 190611 3647 190645
rect 3795 190583 5718 246012
rect 3220 0 5718 190583
rect 40232 -16145 40274 -16111
rect 40328 -16145 40370 -16111
rect 40424 -16145 40466 -16111
rect 40520 -16145 40562 -16111
rect 40616 -16145 40658 -16111
rect 43576 -16145 43618 -16111
rect 43672 -16145 43714 -16111
rect 43768 -16145 43810 -16111
rect 43864 -16145 43906 -16111
rect 43960 -16145 44002 -16111
rect 46920 -16145 46962 -16111
rect 47016 -16145 47058 -16111
rect 47112 -16145 47154 -16111
rect 47208 -16145 47250 -16111
rect 47304 -16145 47346 -16111
rect 50264 -16145 50306 -16111
rect 50360 -16145 50402 -16111
rect 50456 -16145 50498 -16111
rect 50552 -16145 50594 -16111
rect 50648 -16145 50690 -16111
rect 53609 -16145 53650 -16111
rect 53705 -16145 53746 -16111
rect 53801 -16145 53842 -16111
rect 53897 -16145 53938 -16111
rect 53993 -16145 54034 -16111
rect 56953 -16145 56994 -16111
rect 57049 -16145 57090 -16111
rect 57145 -16145 57186 -16111
rect 57241 -16145 57282 -16111
rect 57337 -16145 57378 -16111
rect 60297 -16145 60338 -16111
rect 60393 -16145 60434 -16111
rect 60489 -16145 60530 -16111
rect 60585 -16145 60626 -16111
rect 60681 -16145 60722 -16111
rect 63641 -16145 63682 -16111
rect 63737 -16145 63778 -16111
rect 63833 -16145 63874 -16111
rect 63929 -16145 63970 -16111
rect 64025 -16145 64066 -16111
rect 66985 -16145 67026 -16111
rect 67081 -16145 67122 -16111
rect 67177 -16145 67218 -16111
rect 67273 -16145 67314 -16111
rect 67369 -16145 67410 -16111
rect 70329 -16145 70370 -16111
rect 70425 -16145 70466 -16111
rect 70521 -16145 70562 -16111
rect 70617 -16145 70658 -16111
rect 70713 -16145 70754 -16111
rect 73673 -16145 73714 -16111
rect 73769 -16145 73810 -16111
rect 73865 -16145 73906 -16111
rect 73961 -16145 74002 -16111
rect 74057 -16145 74098 -16111
rect 77017 -16145 77058 -16111
rect 77113 -16145 77154 -16111
rect 77209 -16145 77250 -16111
rect 77305 -16145 77346 -16111
rect 77401 -16145 77442 -16111
rect 80361 -16145 80402 -16111
rect 80457 -16145 80498 -16111
rect 80553 -16145 80594 -16111
rect 80649 -16145 80690 -16111
rect 80745 -16145 80786 -16111
rect 83705 -16145 83746 -16111
rect 83801 -16145 83842 -16111
rect 83897 -16145 83938 -16111
rect 83993 -16145 84034 -16111
rect 84089 -16145 84130 -16111
rect 87049 -16145 87090 -16111
rect 87145 -16145 87186 -16111
rect 87241 -16145 87282 -16111
rect 87337 -16145 87378 -16111
rect 87433 -16145 87474 -16111
rect 90393 -16145 90434 -16111
rect 90489 -16145 90530 -16111
rect 90585 -16145 90626 -16111
rect 90681 -16145 90722 -16111
rect 90777 -16145 90818 -16111
rect 93737 -16145 93778 -16111
rect 93833 -16145 93874 -16111
rect 93929 -16145 93970 -16111
rect 94025 -16145 94066 -16111
rect 94121 -16145 94162 -16111
rect 97081 -16145 97122 -16111
rect 97177 -16145 97218 -16111
rect 97273 -16145 97314 -16111
rect 97369 -16145 97410 -16111
rect 97465 -16145 97506 -16111
rect 100425 -16145 100466 -16111
rect 100521 -16145 100562 -16111
rect 100617 -16145 100658 -16111
rect 100713 -16145 100754 -16111
rect 100809 -16145 100850 -16111
rect 103769 -16145 103810 -16111
rect 103865 -16145 103906 -16111
rect 103961 -16145 104002 -16111
rect 104057 -16145 104098 -16111
rect 104153 -16145 104194 -16111
rect 107119 -16145 107154 -16111
rect 107215 -16145 107250 -16111
rect 107311 -16145 107346 -16111
rect 107407 -16145 107442 -16111
rect 107503 -16145 107538 -16111
rect 110463 -16145 110498 -16111
rect 110559 -16145 110594 -16111
rect 110655 -16145 110690 -16111
rect 110751 -16145 110786 -16111
rect 110847 -16145 110882 -16111
rect 113807 -16145 113842 -16111
rect 113903 -16145 113938 -16111
rect 113999 -16145 114034 -16111
rect 114095 -16145 114130 -16111
rect 114191 -16145 114226 -16111
rect 117151 -16145 117186 -16111
rect 117247 -16145 117282 -16111
rect 117343 -16145 117378 -16111
rect 117439 -16145 117474 -16111
rect 117535 -16145 117570 -16111
rect 120495 -16145 120530 -16111
rect 120591 -16145 120626 -16111
rect 120687 -16145 120722 -16111
rect 120783 -16145 120818 -16111
rect 120879 -16145 120914 -16111
rect 123839 -16145 123874 -16111
rect 123935 -16145 123970 -16111
rect 124031 -16145 124066 -16111
rect 124127 -16145 124162 -16111
rect 124223 -16145 124258 -16111
rect 127183 -16145 127218 -16111
rect 127279 -16145 127314 -16111
rect 127375 -16145 127410 -16111
rect 127471 -16145 127506 -16111
rect 127567 -16145 127602 -16111
rect 130527 -16145 130562 -16111
rect 130623 -16145 130658 -16111
rect 130719 -16145 130754 -16111
rect 130815 -16145 130850 -16111
rect 130911 -16145 130946 -16111
rect 133871 -16145 133906 -16111
rect 133967 -16145 134002 -16111
rect 134063 -16145 134098 -16111
rect 134159 -16145 134194 -16111
rect 134255 -16145 134290 -16111
rect 137215 -16145 137250 -16111
rect 137311 -16145 137346 -16111
rect 137407 -16145 137442 -16111
rect 137503 -16145 137538 -16111
rect 137599 -16145 137634 -16111
rect 140559 -16145 140594 -16111
rect 140655 -16145 140690 -16111
rect 140751 -16145 140786 -16111
rect 140847 -16145 140882 -16111
rect 140943 -16145 140978 -16111
rect 143903 -16145 143938 -16111
rect 143999 -16145 144034 -16111
rect 144095 -16145 144130 -16111
rect 144191 -16145 144226 -16111
rect 144287 -16145 144322 -16111
rect 147247 -16145 147282 -16111
rect 147343 -16145 147378 -16111
rect 147439 -16145 147474 -16111
rect 147535 -16145 147570 -16111
rect 147631 -16145 147666 -16111
rect 150591 -16145 150626 -16111
rect 150687 -16145 150722 -16111
rect 150783 -16145 150818 -16111
rect 150879 -16145 150914 -16111
rect 150975 -16145 151010 -16111
rect 153935 -16145 153970 -16111
rect 154031 -16145 154066 -16111
rect 154127 -16145 154162 -16111
rect 154223 -16145 154258 -16111
rect 154319 -16145 154354 -16111
rect 157279 -16145 157314 -16111
rect 157375 -16145 157410 -16111
rect 157471 -16145 157506 -16111
rect 157567 -16145 157602 -16111
rect 157663 -16145 157698 -16111
rect 160623 -16145 160658 -16111
rect 160719 -16145 160754 -16111
rect 160815 -16145 160850 -16111
rect 160911 -16145 160946 -16111
rect 161007 -16145 161042 -16111
rect 163967 -16145 164002 -16111
rect 164063 -16145 164098 -16111
rect 164159 -16145 164194 -16111
rect 164255 -16145 164290 -16111
rect 164351 -16145 164386 -16111
rect 167311 -16145 167346 -16111
rect 167407 -16145 167442 -16111
rect 167503 -16145 167538 -16111
rect 167599 -16145 167634 -16111
rect 167695 -16145 167730 -16111
rect 170655 -16145 170690 -16111
rect 170751 -16145 170786 -16111
rect 170847 -16145 170882 -16111
rect 170943 -16145 170978 -16111
rect 171039 -16145 171074 -16111
rect 173999 -16145 174034 -16111
rect 174095 -16145 174130 -16111
rect 174191 -16145 174226 -16111
rect 174287 -16145 174322 -16111
rect 174383 -16145 174418 -16111
rect 177343 -16145 177378 -16111
rect 177439 -16145 177474 -16111
rect 177535 -16145 177570 -16111
rect 177631 -16145 177666 -16111
rect 177727 -16145 177762 -16111
rect 180687 -16145 180722 -16111
rect 180783 -16145 180818 -16111
rect 180879 -16145 180914 -16111
rect 180975 -16145 181010 -16111
rect 181071 -16145 181106 -16111
rect 184031 -16145 184066 -16111
rect 184127 -16145 184162 -16111
rect 184223 -16145 184258 -16111
rect 184319 -16145 184354 -16111
rect 184415 -16145 184450 -16111
rect 187375 -16145 187410 -16111
rect 187471 -16145 187506 -16111
rect 187567 -16145 187602 -16111
rect 187663 -16145 187698 -16111
rect 187759 -16145 187794 -16111
rect 190719 -16145 190754 -16111
rect 190815 -16145 190850 -16111
rect 190911 -16145 190946 -16111
rect 191007 -16145 191042 -16111
rect 191103 -16145 191138 -16111
rect 194063 -16145 194098 -16111
rect 194159 -16145 194194 -16111
rect 194255 -16145 194290 -16111
rect 194351 -16145 194386 -16111
rect 194447 -16145 194482 -16111
rect 197407 -16145 197442 -16111
rect 197503 -16145 197538 -16111
rect 197599 -16145 197634 -16111
rect 197695 -16145 197730 -16111
rect 197791 -16145 197826 -16111
rect 200751 -16145 200786 -16111
rect 200847 -16145 200882 -16111
rect 200943 -16145 200978 -16111
rect 201039 -16145 201074 -16111
rect 201135 -16145 201170 -16111
rect 204095 -16145 204130 -16111
rect 204191 -16145 204226 -16111
rect 204287 -16145 204322 -16111
rect 204383 -16145 204418 -16111
rect 204479 -16145 204514 -16111
rect 207439 -16145 207474 -16111
rect 207535 -16145 207570 -16111
rect 207631 -16145 207666 -16111
rect 207727 -16145 207762 -16111
rect 207823 -16145 207858 -16111
rect 210783 -16145 210818 -16111
rect 210879 -16145 210914 -16111
rect 210975 -16145 211010 -16111
rect 211071 -16145 211106 -16111
rect 211167 -16145 211202 -16111
rect 40778 -16188 40820 -16154
rect 40874 -16188 40916 -16154
rect 40970 -16188 41012 -16154
rect 41066 -16188 41108 -16154
rect 41162 -16188 41204 -16154
rect 41258 -16188 41300 -16154
rect 41354 -16188 41396 -16154
rect 44122 -16188 44164 -16154
rect 44218 -16188 44260 -16154
rect 44314 -16188 44356 -16154
rect 44410 -16188 44452 -16154
rect 44506 -16188 44548 -16154
rect 44602 -16188 44644 -16154
rect 44698 -16188 44740 -16154
rect 47466 -16188 47508 -16154
rect 47562 -16188 47604 -16154
rect 47658 -16188 47700 -16154
rect 47754 -16188 47796 -16154
rect 47850 -16188 47892 -16154
rect 47946 -16188 47988 -16154
rect 48042 -16188 48084 -16154
rect 50810 -16188 50852 -16154
rect 50906 -16188 50948 -16154
rect 51002 -16188 51044 -16154
rect 51098 -16188 51140 -16154
rect 51194 -16188 51236 -16154
rect 51290 -16188 51332 -16154
rect 51386 -16188 51428 -16154
rect 54155 -16188 54196 -16154
rect 54251 -16188 54292 -16154
rect 54347 -16188 54388 -16154
rect 54443 -16188 54484 -16154
rect 54539 -16188 54580 -16154
rect 54635 -16188 54676 -16154
rect 54731 -16188 54772 -16154
rect 57499 -16188 57540 -16154
rect 57595 -16188 57636 -16154
rect 57691 -16188 57732 -16154
rect 57787 -16188 57828 -16154
rect 57883 -16188 57924 -16154
rect 57979 -16188 58020 -16154
rect 58075 -16188 58116 -16154
rect 60843 -16188 60884 -16154
rect 60939 -16188 60980 -16154
rect 61035 -16188 61076 -16154
rect 61131 -16188 61172 -16154
rect 61227 -16188 61268 -16154
rect 61323 -16188 61364 -16154
rect 61419 -16188 61460 -16154
rect 64187 -16188 64228 -16154
rect 64283 -16188 64324 -16154
rect 64379 -16188 64420 -16154
rect 64475 -16188 64516 -16154
rect 64571 -16188 64612 -16154
rect 64667 -16188 64708 -16154
rect 64763 -16188 64804 -16154
rect 67531 -16188 67572 -16154
rect 67627 -16188 67668 -16154
rect 67723 -16188 67764 -16154
rect 67819 -16188 67860 -16154
rect 67915 -16188 67956 -16154
rect 68011 -16188 68052 -16154
rect 68107 -16188 68148 -16154
rect 70875 -16188 70916 -16154
rect 70971 -16188 71012 -16154
rect 71067 -16188 71108 -16154
rect 71163 -16188 71204 -16154
rect 71259 -16188 71300 -16154
rect 71355 -16188 71396 -16154
rect 71451 -16188 71492 -16154
rect 74219 -16188 74260 -16154
rect 74315 -16188 74356 -16154
rect 74411 -16188 74452 -16154
rect 74507 -16188 74548 -16154
rect 74603 -16188 74644 -16154
rect 74699 -16188 74740 -16154
rect 74795 -16188 74836 -16154
rect 77563 -16188 77604 -16154
rect 77659 -16188 77700 -16154
rect 77755 -16188 77796 -16154
rect 77851 -16188 77892 -16154
rect 77947 -16188 77988 -16154
rect 78043 -16188 78084 -16154
rect 78139 -16188 78180 -16154
rect 80907 -16188 80948 -16154
rect 81003 -16188 81044 -16154
rect 81099 -16188 81140 -16154
rect 81195 -16188 81236 -16154
rect 81291 -16188 81332 -16154
rect 81387 -16188 81428 -16154
rect 81483 -16188 81524 -16154
rect 84251 -16188 84292 -16154
rect 84347 -16188 84388 -16154
rect 84443 -16188 84484 -16154
rect 84539 -16188 84580 -16154
rect 84635 -16188 84676 -16154
rect 84731 -16188 84772 -16154
rect 84827 -16188 84868 -16154
rect 87595 -16188 87636 -16154
rect 87691 -16188 87732 -16154
rect 87787 -16188 87828 -16154
rect 87883 -16188 87924 -16154
rect 87979 -16188 88020 -16154
rect 88075 -16188 88116 -16154
rect 88171 -16188 88212 -16154
rect 90939 -16188 90980 -16154
rect 91035 -16188 91076 -16154
rect 91131 -16188 91172 -16154
rect 91227 -16188 91268 -16154
rect 91323 -16188 91364 -16154
rect 91419 -16188 91460 -16154
rect 91515 -16188 91556 -16154
rect 94283 -16188 94324 -16154
rect 94379 -16188 94420 -16154
rect 94475 -16188 94516 -16154
rect 94571 -16188 94612 -16154
rect 94667 -16188 94708 -16154
rect 94763 -16188 94804 -16154
rect 94859 -16188 94900 -16154
rect 97627 -16188 97668 -16154
rect 97723 -16188 97764 -16154
rect 97819 -16188 97860 -16154
rect 97915 -16188 97956 -16154
rect 98011 -16188 98052 -16154
rect 98107 -16188 98148 -16154
rect 98203 -16188 98244 -16154
rect 100971 -16188 101012 -16154
rect 101067 -16188 101108 -16154
rect 101163 -16188 101204 -16154
rect 101259 -16188 101300 -16154
rect 101355 -16188 101396 -16154
rect 101451 -16188 101492 -16154
rect 101547 -16188 101588 -16154
rect 104315 -16188 104356 -16154
rect 104411 -16188 104452 -16154
rect 104507 -16188 104548 -16154
rect 104603 -16188 104644 -16154
rect 104699 -16188 104740 -16154
rect 104795 -16188 104836 -16154
rect 104891 -16188 104932 -16154
rect 107665 -16188 107700 -16154
rect 107761 -16188 107796 -16154
rect 107857 -16188 107892 -16154
rect 107953 -16188 107988 -16154
rect 108049 -16188 108084 -16154
rect 108145 -16188 108180 -16154
rect 108241 -16188 108276 -16154
rect 111009 -16188 111044 -16154
rect 111105 -16188 111140 -16154
rect 111201 -16188 111236 -16154
rect 111297 -16188 111332 -16154
rect 111393 -16188 111428 -16154
rect 111489 -16188 111524 -16154
rect 111585 -16188 111620 -16154
rect 114353 -16188 114388 -16154
rect 114449 -16188 114484 -16154
rect 114545 -16188 114580 -16154
rect 114641 -16188 114676 -16154
rect 114737 -16188 114772 -16154
rect 114833 -16188 114868 -16154
rect 114929 -16188 114964 -16154
rect 117697 -16188 117732 -16154
rect 117793 -16188 117828 -16154
rect 117889 -16188 117924 -16154
rect 117985 -16188 118020 -16154
rect 118081 -16188 118116 -16154
rect 118177 -16188 118212 -16154
rect 118273 -16188 118308 -16154
rect 121041 -16188 121076 -16154
rect 121137 -16188 121172 -16154
rect 121233 -16188 121268 -16154
rect 121329 -16188 121364 -16154
rect 121425 -16188 121460 -16154
rect 121521 -16188 121556 -16154
rect 121617 -16188 121652 -16154
rect 124385 -16188 124420 -16154
rect 124481 -16188 124516 -16154
rect 124577 -16188 124612 -16154
rect 124673 -16188 124708 -16154
rect 124769 -16188 124804 -16154
rect 124865 -16188 124900 -16154
rect 124961 -16188 124996 -16154
rect 127729 -16188 127764 -16154
rect 127825 -16188 127860 -16154
rect 127921 -16188 127956 -16154
rect 128017 -16188 128052 -16154
rect 128113 -16188 128148 -16154
rect 128209 -16188 128244 -16154
rect 128305 -16188 128340 -16154
rect 131073 -16188 131108 -16154
rect 131169 -16188 131204 -16154
rect 131265 -16188 131300 -16154
rect 131361 -16188 131396 -16154
rect 131457 -16188 131492 -16154
rect 131553 -16188 131588 -16154
rect 131649 -16188 131684 -16154
rect 134417 -16188 134452 -16154
rect 134513 -16188 134548 -16154
rect 134609 -16188 134644 -16154
rect 134705 -16188 134740 -16154
rect 134801 -16188 134836 -16154
rect 134897 -16188 134932 -16154
rect 134993 -16188 135028 -16154
rect 137761 -16188 137796 -16154
rect 137857 -16188 137892 -16154
rect 137953 -16188 137988 -16154
rect 138049 -16188 138084 -16154
rect 138145 -16188 138180 -16154
rect 138241 -16188 138276 -16154
rect 138337 -16188 138372 -16154
rect 141105 -16188 141140 -16154
rect 141201 -16188 141236 -16154
rect 141297 -16188 141332 -16154
rect 141393 -16188 141428 -16154
rect 141489 -16188 141524 -16154
rect 141585 -16188 141620 -16154
rect 141681 -16188 141716 -16154
rect 144449 -16188 144484 -16154
rect 144545 -16188 144580 -16154
rect 144641 -16188 144676 -16154
rect 144737 -16188 144772 -16154
rect 144833 -16188 144868 -16154
rect 144929 -16188 144964 -16154
rect 145025 -16188 145060 -16154
rect 147793 -16188 147828 -16154
rect 147889 -16188 147924 -16154
rect 147985 -16188 148020 -16154
rect 148081 -16188 148116 -16154
rect 148177 -16188 148212 -16154
rect 148273 -16188 148308 -16154
rect 148369 -16188 148404 -16154
rect 151137 -16188 151172 -16154
rect 151233 -16188 151268 -16154
rect 151329 -16188 151364 -16154
rect 151425 -16188 151460 -16154
rect 151521 -16188 151556 -16154
rect 151617 -16188 151652 -16154
rect 151713 -16188 151748 -16154
rect 154481 -16188 154516 -16154
rect 154577 -16188 154612 -16154
rect 154673 -16188 154708 -16154
rect 154769 -16188 154804 -16154
rect 154865 -16188 154900 -16154
rect 154961 -16188 154996 -16154
rect 155057 -16188 155092 -16154
rect 157825 -16188 157860 -16154
rect 157921 -16188 157956 -16154
rect 158017 -16188 158052 -16154
rect 158113 -16188 158148 -16154
rect 158209 -16188 158244 -16154
rect 158305 -16188 158340 -16154
rect 158401 -16188 158436 -16154
rect 161169 -16188 161204 -16154
rect 161265 -16188 161300 -16154
rect 161361 -16188 161396 -16154
rect 161457 -16188 161492 -16154
rect 161553 -16188 161588 -16154
rect 161649 -16188 161684 -16154
rect 161745 -16188 161780 -16154
rect 164513 -16188 164548 -16154
rect 164609 -16188 164644 -16154
rect 164705 -16188 164740 -16154
rect 164801 -16188 164836 -16154
rect 164897 -16188 164932 -16154
rect 164993 -16188 165028 -16154
rect 165089 -16188 165124 -16154
rect 167857 -16188 167892 -16154
rect 167953 -16188 167988 -16154
rect 168049 -16188 168084 -16154
rect 168145 -16188 168180 -16154
rect 168241 -16188 168276 -16154
rect 168337 -16188 168372 -16154
rect 168433 -16188 168468 -16154
rect 171201 -16188 171236 -16154
rect 171297 -16188 171332 -16154
rect 171393 -16188 171428 -16154
rect 171489 -16188 171524 -16154
rect 171585 -16188 171620 -16154
rect 171681 -16188 171716 -16154
rect 171777 -16188 171812 -16154
rect 174545 -16188 174580 -16154
rect 174641 -16188 174676 -16154
rect 174737 -16188 174772 -16154
rect 174833 -16188 174868 -16154
rect 174929 -16188 174964 -16154
rect 175025 -16188 175060 -16154
rect 175121 -16188 175156 -16154
rect 177889 -16188 177924 -16154
rect 177985 -16188 178020 -16154
rect 178081 -16188 178116 -16154
rect 178177 -16188 178212 -16154
rect 178273 -16188 178308 -16154
rect 178369 -16188 178404 -16154
rect 178465 -16188 178500 -16154
rect 181233 -16188 181268 -16154
rect 181329 -16188 181364 -16154
rect 181425 -16188 181460 -16154
rect 181521 -16188 181556 -16154
rect 181617 -16188 181652 -16154
rect 181713 -16188 181748 -16154
rect 181809 -16188 181844 -16154
rect 184577 -16188 184612 -16154
rect 184673 -16188 184708 -16154
rect 184769 -16188 184804 -16154
rect 184865 -16188 184900 -16154
rect 184961 -16188 184996 -16154
rect 185057 -16188 185092 -16154
rect 185153 -16188 185188 -16154
rect 187921 -16188 187956 -16154
rect 188017 -16188 188052 -16154
rect 188113 -16188 188148 -16154
rect 188209 -16188 188244 -16154
rect 188305 -16188 188340 -16154
rect 188401 -16188 188436 -16154
rect 188497 -16188 188532 -16154
rect 191265 -16188 191300 -16154
rect 191361 -16188 191396 -16154
rect 191457 -16188 191492 -16154
rect 191553 -16188 191588 -16154
rect 191649 -16188 191684 -16154
rect 191745 -16188 191780 -16154
rect 191841 -16188 191876 -16154
rect 194609 -16188 194644 -16154
rect 194705 -16188 194740 -16154
rect 194801 -16188 194836 -16154
rect 194897 -16188 194932 -16154
rect 194993 -16188 195028 -16154
rect 195089 -16188 195124 -16154
rect 195185 -16188 195220 -16154
rect 197953 -16188 197988 -16154
rect 198049 -16188 198084 -16154
rect 198145 -16188 198180 -16154
rect 198241 -16188 198276 -16154
rect 198337 -16188 198372 -16154
rect 198433 -16188 198468 -16154
rect 198529 -16188 198564 -16154
rect 201297 -16188 201332 -16154
rect 201393 -16188 201428 -16154
rect 201489 -16188 201524 -16154
rect 201585 -16188 201620 -16154
rect 201681 -16188 201716 -16154
rect 201777 -16188 201812 -16154
rect 201873 -16188 201908 -16154
rect 204641 -16188 204676 -16154
rect 204737 -16188 204772 -16154
rect 204833 -16188 204868 -16154
rect 204929 -16188 204964 -16154
rect 205025 -16188 205060 -16154
rect 205121 -16188 205156 -16154
rect 205217 -16188 205252 -16154
rect 207985 -16188 208020 -16154
rect 208081 -16188 208116 -16154
rect 208177 -16188 208212 -16154
rect 208273 -16188 208308 -16154
rect 208369 -16188 208404 -16154
rect 208465 -16188 208500 -16154
rect 208561 -16188 208596 -16154
rect 211329 -16188 211364 -16154
rect 211425 -16188 211460 -16154
rect 211521 -16188 211556 -16154
rect 211617 -16188 211652 -16154
rect 211713 -16188 211748 -16154
rect 211809 -16188 211844 -16154
rect 211905 -16188 211940 -16154
rect 38274 -16231 38310 -16197
rect 38364 -16231 38406 -16197
rect 40334 -16207 40342 -16199
rect 40411 -16207 40417 -16191
rect 40434 -16207 40442 -16199
rect 40445 -16207 40451 -16191
rect 38526 -16274 38568 -16240
rect 38622 -16274 38664 -16240
rect 38718 -16274 38760 -16240
rect 40225 -16241 40267 -16207
rect 40289 -16241 40342 -16207
rect 40369 -16241 40417 -16207
rect 38338 -16293 38346 -16285
rect 38274 -16327 38279 -16293
rect 38349 -16327 38391 -16293
rect 38880 -16317 38922 -16283
rect 38976 -16317 39018 -16283
rect 39072 -16317 39114 -16283
rect 39168 -16317 39210 -16283
rect 39264 -16317 39306 -16283
rect 40289 -16324 40331 -16290
rect 40334 -16324 40342 -16279
rect 38592 -16336 38600 -16328
rect 38692 -16336 38700 -16328
rect 38338 -16376 38346 -16365
rect 38519 -16370 38589 -16336
rect 38591 -16370 38633 -16336
rect 38703 -16370 38745 -16336
rect 39428 -16360 39470 -16326
rect 39524 -16360 39566 -16326
rect 39620 -16360 39662 -16326
rect 39716 -16360 39758 -16326
rect 39812 -16360 39854 -16326
rect 39908 -16360 39950 -16326
rect 40004 -16360 40046 -16326
rect 38349 -16410 38391 -16376
rect 38982 -16379 38990 -16371
rect 39059 -16379 39065 -16363
rect 39082 -16379 39090 -16371
rect 39093 -16379 39099 -16363
rect 38338 -16460 38346 -16449
rect 38547 -16453 38589 -16419
rect 38592 -16453 38600 -16408
rect 38692 -16419 38700 -16408
rect 38873 -16413 38915 -16379
rect 38937 -16413 38990 -16379
rect 39017 -16413 39065 -16379
rect 38703 -16453 38745 -16419
rect 38349 -16494 38391 -16460
rect 38338 -16543 38346 -16532
rect 38547 -16537 38589 -16503
rect 38592 -16537 38600 -16492
rect 38692 -16503 38700 -16492
rect 38937 -16496 38979 -16462
rect 38982 -16496 38990 -16451
rect 38703 -16537 38745 -16503
rect 38349 -16577 38391 -16543
rect 38274 -16691 38300 -16657
rect 38310 -16718 38316 -16641
rect 38344 -16752 38350 -16607
rect 38547 -16620 38589 -16586
rect 38592 -16620 38600 -16575
rect 38692 -16586 38700 -16575
rect 38937 -16580 38979 -16546
rect 38982 -16580 38990 -16535
rect 38703 -16620 38745 -16586
rect 38612 -16734 38654 -16700
rect 38664 -16761 38670 -16684
rect 38342 -16779 38350 -16771
rect 38353 -16813 38395 -16779
rect 38698 -16795 38704 -16650
rect 38937 -16663 38979 -16629
rect 38982 -16663 38990 -16618
rect 39059 -16679 39065 -16413
rect 39093 -16413 39135 -16379
rect 39138 -16413 39146 -16371
rect 39082 -16462 39090 -16451
rect 39093 -16462 39099 -16413
rect 39093 -16496 39135 -16462
rect 39138 -16496 39146 -16451
rect 39082 -16546 39090 -16535
rect 39093 -16546 39099 -16496
rect 39093 -16580 39135 -16546
rect 39138 -16580 39146 -16535
rect 39082 -16629 39090 -16618
rect 39093 -16629 39099 -16580
rect 39093 -16663 39135 -16629
rect 39138 -16663 39146 -16618
rect 39082 -16697 39090 -16671
rect 39093 -16713 39099 -16663
rect 39002 -16777 39044 -16743
rect 39059 -16804 39060 -16727
rect 39093 -16809 39094 -16713
rect 38551 -16856 38593 -16822
rect 38596 -16856 38604 -16814
rect 38696 -16822 38704 -16814
rect 38707 -16856 38749 -16822
rect 39124 -16845 39132 -16697
rect 39147 -16713 39151 -16363
rect 39181 -16679 39185 -16363
rect 39238 -16379 39246 -16371
rect 39187 -16413 39229 -16379
rect 39249 -16413 39301 -16379
rect 39959 -16422 39965 -16406
rect 39982 -16422 39990 -16414
rect 39993 -16422 39999 -16406
rect 40289 -16408 40331 -16374
rect 40334 -16408 40342 -16363
rect 39238 -16462 39246 -16451
rect 39419 -16456 39461 -16422
rect 39491 -16456 39533 -16422
rect 39563 -16456 39605 -16422
rect 39707 -16456 39749 -16422
rect 39779 -16456 39893 -16422
rect 39923 -16456 39965 -16422
rect 39249 -16496 39291 -16462
rect 39238 -16546 39246 -16535
rect 39816 -16539 39858 -16505
rect 39249 -16580 39291 -16546
rect 39238 -16629 39246 -16618
rect 39249 -16663 39291 -16629
rect 39481 -16689 39523 -16655
rect 39526 -16689 39534 -16644
rect 39603 -16706 39609 -16588
rect 39626 -16655 39634 -16644
rect 39637 -16655 39643 -16622
rect 39673 -16655 39679 -16622
rect 39637 -16689 39679 -16655
rect 39682 -16689 39690 -16644
rect 39637 -16740 39643 -16689
rect 39673 -16740 39679 -16689
rect 39707 -16706 39713 -16589
rect 39804 -16630 39805 -16589
rect 39816 -16623 39858 -16589
rect 39816 -16706 39858 -16672
rect 39959 -16706 39965 -16456
rect 39993 -16456 40035 -16422
rect 39982 -16505 39990 -16494
rect 39993 -16505 39999 -16456
rect 40289 -16491 40331 -16457
rect 40334 -16491 40342 -16446
rect 39993 -16539 40035 -16505
rect 39982 -16589 39990 -16578
rect 39993 -16589 39999 -16539
rect 40143 -16565 40251 -16499
rect 40411 -16507 40417 -16241
rect 40445 -16241 40487 -16207
rect 40490 -16241 40498 -16199
rect 40434 -16290 40442 -16279
rect 40445 -16290 40451 -16241
rect 40445 -16324 40487 -16290
rect 40490 -16324 40498 -16279
rect 40434 -16374 40442 -16363
rect 40445 -16374 40451 -16324
rect 40445 -16408 40487 -16374
rect 40490 -16408 40498 -16363
rect 40434 -16457 40442 -16446
rect 40445 -16457 40451 -16408
rect 40445 -16491 40487 -16457
rect 40490 -16491 40498 -16446
rect 40434 -16525 40442 -16499
rect 40445 -16541 40451 -16491
rect 39993 -16623 40035 -16589
rect 40354 -16605 40396 -16571
rect 39982 -16672 39990 -16661
rect 39993 -16672 39999 -16623
rect 40411 -16632 40412 -16555
rect 40445 -16637 40446 -16541
rect 39993 -16706 40035 -16672
rect 40476 -16673 40484 -16525
rect 40499 -16541 40503 -16191
rect 40533 -16507 40537 -16191
rect 40590 -16207 40598 -16199
rect 40539 -16241 40581 -16207
rect 40601 -16241 40653 -16207
rect 41516 -16231 41558 -16197
rect 41612 -16231 41654 -16197
rect 41708 -16231 41750 -16197
rect 43678 -16207 43686 -16199
rect 43755 -16207 43761 -16191
rect 43778 -16207 43786 -16199
rect 43789 -16207 43795 -16191
rect 41309 -16250 41315 -16234
rect 41332 -16250 41340 -16242
rect 41343 -16250 41349 -16234
rect 40590 -16290 40598 -16279
rect 40769 -16284 40811 -16250
rect 40841 -16284 40883 -16250
rect 40913 -16284 40955 -16250
rect 41057 -16284 41099 -16250
rect 41129 -16284 41243 -16250
rect 41273 -16284 41315 -16250
rect 40601 -16324 40643 -16290
rect 40590 -16374 40598 -16363
rect 41166 -16367 41208 -16333
rect 40601 -16408 40643 -16374
rect 40590 -16457 40598 -16446
rect 40601 -16491 40643 -16457
rect 40831 -16517 40873 -16483
rect 40876 -16517 40884 -16472
rect 40953 -16534 40959 -16416
rect 40976 -16483 40984 -16472
rect 40987 -16483 40993 -16450
rect 41023 -16483 41029 -16450
rect 40987 -16517 41029 -16483
rect 41032 -16517 41040 -16472
rect 40987 -16568 40993 -16517
rect 41023 -16568 41029 -16517
rect 41057 -16534 41063 -16417
rect 41154 -16458 41155 -16417
rect 41166 -16451 41208 -16417
rect 41166 -16534 41208 -16500
rect 41309 -16534 41315 -16284
rect 41343 -16284 41385 -16250
rect 41870 -16274 41912 -16240
rect 41966 -16274 42008 -16240
rect 42062 -16274 42104 -16240
rect 43569 -16241 43611 -16207
rect 43633 -16241 43686 -16207
rect 43713 -16241 43761 -16207
rect 41332 -16333 41340 -16322
rect 41343 -16333 41349 -16284
rect 41582 -16293 41590 -16285
rect 41682 -16293 41690 -16285
rect 41509 -16327 41579 -16293
rect 41581 -16327 41623 -16293
rect 41693 -16327 41735 -16293
rect 42224 -16317 42266 -16283
rect 42320 -16317 42362 -16283
rect 42416 -16317 42458 -16283
rect 42512 -16317 42554 -16283
rect 42608 -16317 42650 -16283
rect 43633 -16324 43675 -16290
rect 43678 -16324 43686 -16279
rect 41343 -16367 41385 -16333
rect 41936 -16336 41944 -16328
rect 42036 -16336 42044 -16328
rect 41332 -16417 41340 -16406
rect 41343 -16417 41349 -16367
rect 41537 -16410 41579 -16376
rect 41582 -16410 41590 -16365
rect 41682 -16376 41690 -16365
rect 41863 -16370 41933 -16336
rect 41935 -16370 41977 -16336
rect 42047 -16370 42089 -16336
rect 42772 -16360 42814 -16326
rect 42868 -16360 42910 -16326
rect 42964 -16360 43006 -16326
rect 43060 -16360 43102 -16326
rect 43156 -16360 43198 -16326
rect 43252 -16360 43294 -16326
rect 43348 -16360 43390 -16326
rect 41693 -16410 41735 -16376
rect 42326 -16379 42334 -16371
rect 42403 -16379 42409 -16363
rect 42426 -16379 42434 -16371
rect 42437 -16379 42443 -16363
rect 41343 -16451 41385 -16417
rect 41332 -16500 41340 -16489
rect 41343 -16500 41349 -16451
rect 41537 -16494 41579 -16460
rect 41582 -16494 41590 -16449
rect 41682 -16460 41690 -16449
rect 41891 -16453 41933 -16419
rect 41936 -16453 41944 -16408
rect 42036 -16419 42044 -16408
rect 42217 -16413 42259 -16379
rect 42281 -16413 42334 -16379
rect 42361 -16413 42409 -16379
rect 42047 -16453 42089 -16419
rect 41693 -16494 41735 -16460
rect 41343 -16534 41385 -16500
rect 41343 -16568 41349 -16534
rect 39993 -16740 39999 -16706
rect 40289 -16723 40331 -16689
rect 40334 -16723 40342 -16681
rect 38342 -16879 38350 -16868
rect 38353 -16913 38395 -16879
rect 38937 -16895 38979 -16861
rect 38982 -16895 38990 -16853
rect 38274 -16949 38279 -16915
rect 38551 -16956 38593 -16922
rect 38596 -16956 38604 -16911
rect 38696 -16922 38704 -16911
rect 39124 -16913 39137 -16845
rect 39165 -16879 39171 -16811
rect 39210 -16843 39216 -16775
rect 39244 -16809 39250 -16743
rect 39254 -16793 39296 -16759
rect 39457 -16838 39499 -16804
rect 39224 -16861 39232 -16853
rect 39235 -16895 39277 -16861
rect 39457 -16906 39499 -16872
rect 38707 -16956 38749 -16922
rect 38519 -16992 38561 -16958
rect 38591 -16992 38633 -16958
rect 38937 -16995 38979 -16961
rect 38982 -16995 38990 -16950
rect 39124 -17001 39132 -16913
rect 39506 -16922 39512 -16788
rect 39224 -16961 39232 -16950
rect 39540 -16956 39546 -16762
rect 39580 -16778 39588 -16767
rect 39576 -16809 39588 -16778
rect 39902 -16796 39944 -16762
rect 39235 -16995 39277 -16961
rect 38274 -17045 38310 -17011
rect 38364 -17045 38406 -17011
rect 38873 -17035 38915 -17001
rect 38945 -17035 38987 -17001
rect 39017 -17035 39059 -17001
rect 39089 -17029 39132 -17001
rect 39435 -17025 39477 -16991
rect 39480 -17025 39488 -16980
rect 39576 -16992 39582 -16809
rect 39610 -16995 39616 -16812
rect 39089 -17035 39131 -17029
rect 38526 -17088 38568 -17054
rect 38622 -17088 38664 -17054
rect 38718 -17088 38760 -17054
rect 39622 -17076 39630 -16809
rect 39959 -16812 39960 -16742
rect 39993 -16819 39994 -16740
rect 40476 -16741 40489 -16673
rect 40517 -16707 40523 -16639
rect 40562 -16671 40568 -16603
rect 40596 -16637 40602 -16571
rect 40606 -16621 40648 -16587
rect 40807 -16666 40849 -16632
rect 40576 -16689 40584 -16681
rect 40587 -16723 40629 -16689
rect 40807 -16734 40849 -16700
rect 40476 -16753 40484 -16741
rect 40856 -16750 40862 -16616
rect 40251 -16819 40645 -16753
rect 40890 -16784 40896 -16590
rect 40930 -16606 40938 -16595
rect 40926 -16637 40938 -16606
rect 41252 -16624 41294 -16590
rect 39638 -16860 39680 -16826
rect 39987 -16830 40005 -16819
rect 39987 -16832 39994 -16830
rect 39638 -16928 39680 -16894
rect 39690 -16995 39696 -16860
rect 39921 -16874 39994 -16832
rect 40049 -16874 40645 -16819
rect 40785 -16853 40827 -16819
rect 40830 -16853 40838 -16808
rect 40926 -16820 40932 -16637
rect 40960 -16823 40966 -16640
rect 39921 -16877 40645 -16874
rect 39724 -16980 39730 -16892
rect 39841 -16942 39883 -16908
rect 39886 -16942 39894 -16900
rect 39722 -16991 39730 -16980
rect 39724 -17025 39730 -16991
rect 39733 -17025 39775 -16991
rect 39841 -17042 39883 -17008
rect 39886 -17042 39894 -16997
rect 39734 -17078 39776 -17044
rect 39806 -17078 39848 -17044
rect 39878 -17078 39920 -17044
rect 38880 -17131 38922 -17097
rect 38976 -17131 39018 -17097
rect 39072 -17131 39114 -17097
rect 39168 -17131 39210 -17097
rect 39264 -17131 39306 -17097
rect 39921 -17114 40073 -16877
rect 40251 -16899 40645 -16877
rect 40175 -16925 40645 -16899
rect 40972 -16904 40980 -16637
rect 41309 -16640 41310 -16570
rect 40988 -16688 41030 -16654
rect 41343 -16674 41344 -16568
rect 41537 -16577 41579 -16543
rect 41582 -16577 41590 -16532
rect 41682 -16543 41690 -16532
rect 41891 -16537 41933 -16503
rect 41936 -16537 41944 -16492
rect 42036 -16503 42044 -16492
rect 42281 -16496 42323 -16462
rect 42326 -16496 42334 -16451
rect 42047 -16537 42089 -16503
rect 41693 -16577 41735 -16543
rect 40988 -16756 41030 -16722
rect 41040 -16823 41046 -16688
rect 41602 -16691 41644 -16657
rect 41654 -16718 41660 -16641
rect 41074 -16808 41080 -16720
rect 41191 -16770 41233 -16736
rect 41236 -16770 41244 -16728
rect 41336 -16740 41344 -16729
rect 41347 -16774 41389 -16740
rect 41688 -16752 41694 -16607
rect 41891 -16620 41933 -16586
rect 41936 -16620 41944 -16575
rect 42036 -16586 42044 -16575
rect 42281 -16580 42323 -16546
rect 42326 -16580 42334 -16535
rect 42047 -16620 42089 -16586
rect 41956 -16734 41998 -16700
rect 42008 -16761 42014 -16684
rect 41072 -16819 41080 -16808
rect 41541 -16813 41583 -16779
rect 41586 -16813 41594 -16771
rect 41686 -16779 41694 -16771
rect 41697 -16813 41739 -16779
rect 42042 -16795 42048 -16650
rect 42281 -16663 42323 -16629
rect 42326 -16663 42334 -16618
rect 42403 -16679 42409 -16413
rect 42437 -16413 42479 -16379
rect 42482 -16413 42490 -16371
rect 42426 -16462 42434 -16451
rect 42437 -16462 42443 -16413
rect 42437 -16496 42479 -16462
rect 42482 -16496 42490 -16451
rect 42426 -16546 42434 -16535
rect 42437 -16546 42443 -16496
rect 42437 -16580 42479 -16546
rect 42482 -16580 42490 -16535
rect 42426 -16629 42434 -16618
rect 42437 -16629 42443 -16580
rect 42437 -16663 42479 -16629
rect 42482 -16663 42490 -16618
rect 42426 -16697 42434 -16671
rect 42437 -16713 42443 -16663
rect 42346 -16777 42388 -16743
rect 42403 -16804 42404 -16727
rect 42437 -16809 42438 -16713
rect 41074 -16853 41080 -16819
rect 41083 -16853 41125 -16819
rect 41191 -16870 41233 -16836
rect 41236 -16870 41244 -16825
rect 41336 -16832 41344 -16821
rect 41347 -16866 41389 -16832
rect 41895 -16856 41937 -16822
rect 41940 -16856 41948 -16814
rect 42040 -16822 42048 -16814
rect 42051 -16856 42093 -16822
rect 42468 -16845 42476 -16697
rect 42491 -16713 42495 -16363
rect 42525 -16679 42529 -16363
rect 42582 -16379 42590 -16371
rect 42531 -16413 42573 -16379
rect 42593 -16413 42645 -16379
rect 43303 -16422 43309 -16406
rect 43326 -16422 43334 -16414
rect 43337 -16422 43343 -16406
rect 43633 -16408 43675 -16374
rect 43678 -16408 43686 -16363
rect 42582 -16462 42590 -16451
rect 42763 -16456 42805 -16422
rect 42835 -16456 42877 -16422
rect 42907 -16456 42949 -16422
rect 43051 -16456 43093 -16422
rect 43123 -16456 43237 -16422
rect 43267 -16456 43309 -16422
rect 42593 -16496 42635 -16462
rect 42582 -16546 42590 -16535
rect 43160 -16539 43202 -16505
rect 42593 -16580 42635 -16546
rect 42582 -16629 42590 -16618
rect 42593 -16663 42635 -16629
rect 42825 -16689 42867 -16655
rect 42870 -16689 42878 -16644
rect 42947 -16706 42953 -16588
rect 42970 -16655 42978 -16644
rect 42981 -16655 42987 -16622
rect 43017 -16655 43023 -16622
rect 42981 -16689 43023 -16655
rect 43026 -16689 43034 -16644
rect 42981 -16740 42987 -16689
rect 43017 -16740 43023 -16689
rect 43051 -16706 43057 -16589
rect 43148 -16630 43149 -16589
rect 43160 -16623 43202 -16589
rect 43160 -16706 43202 -16672
rect 43303 -16706 43309 -16456
rect 43337 -16456 43379 -16422
rect 43326 -16505 43334 -16494
rect 43337 -16505 43343 -16456
rect 43633 -16491 43675 -16457
rect 43678 -16491 43686 -16446
rect 43337 -16539 43379 -16505
rect 43326 -16589 43334 -16578
rect 43337 -16589 43343 -16539
rect 43487 -16565 43595 -16499
rect 43755 -16507 43761 -16241
rect 43789 -16241 43831 -16207
rect 43834 -16241 43842 -16199
rect 43778 -16290 43786 -16279
rect 43789 -16290 43795 -16241
rect 43789 -16324 43831 -16290
rect 43834 -16324 43842 -16279
rect 43778 -16374 43786 -16363
rect 43789 -16374 43795 -16324
rect 43789 -16408 43831 -16374
rect 43834 -16408 43842 -16363
rect 43778 -16457 43786 -16446
rect 43789 -16457 43795 -16408
rect 43789 -16491 43831 -16457
rect 43834 -16491 43842 -16446
rect 43778 -16525 43786 -16499
rect 43789 -16541 43795 -16491
rect 43337 -16623 43379 -16589
rect 43698 -16605 43740 -16571
rect 43326 -16672 43334 -16661
rect 43337 -16672 43343 -16623
rect 43755 -16632 43756 -16555
rect 43789 -16637 43790 -16541
rect 43337 -16706 43379 -16672
rect 43820 -16673 43828 -16525
rect 43843 -16541 43847 -16191
rect 43877 -16507 43881 -16191
rect 43934 -16207 43942 -16199
rect 43883 -16241 43925 -16207
rect 43945 -16241 43997 -16207
rect 44860 -16231 44902 -16197
rect 44956 -16231 44998 -16197
rect 45052 -16231 45094 -16197
rect 47022 -16207 47030 -16199
rect 47099 -16207 47105 -16191
rect 47122 -16207 47130 -16199
rect 47133 -16207 47139 -16191
rect 44653 -16250 44659 -16234
rect 44676 -16250 44684 -16242
rect 44687 -16250 44693 -16234
rect 43934 -16290 43942 -16279
rect 44113 -16284 44155 -16250
rect 44185 -16284 44227 -16250
rect 44257 -16284 44299 -16250
rect 44401 -16284 44443 -16250
rect 44473 -16284 44587 -16250
rect 44617 -16284 44659 -16250
rect 43945 -16324 43987 -16290
rect 43934 -16374 43942 -16363
rect 44510 -16367 44552 -16333
rect 43945 -16408 43987 -16374
rect 43934 -16457 43942 -16446
rect 43945 -16491 43987 -16457
rect 44175 -16517 44217 -16483
rect 44220 -16517 44228 -16472
rect 44297 -16534 44303 -16416
rect 44320 -16483 44328 -16472
rect 44331 -16483 44337 -16450
rect 44367 -16483 44373 -16450
rect 44331 -16517 44373 -16483
rect 44376 -16517 44384 -16472
rect 44331 -16568 44337 -16517
rect 44367 -16568 44373 -16517
rect 44401 -16534 44407 -16417
rect 44498 -16458 44499 -16417
rect 44510 -16451 44552 -16417
rect 44510 -16534 44552 -16500
rect 44653 -16534 44659 -16284
rect 44687 -16284 44729 -16250
rect 45214 -16274 45256 -16240
rect 45310 -16274 45352 -16240
rect 45406 -16274 45448 -16240
rect 46913 -16241 46955 -16207
rect 46977 -16241 47030 -16207
rect 47057 -16241 47105 -16207
rect 44676 -16333 44684 -16322
rect 44687 -16333 44693 -16284
rect 44926 -16293 44934 -16285
rect 45026 -16293 45034 -16285
rect 44853 -16327 44923 -16293
rect 44925 -16327 44967 -16293
rect 45037 -16327 45079 -16293
rect 45568 -16317 45610 -16283
rect 45664 -16317 45706 -16283
rect 45760 -16317 45802 -16283
rect 45856 -16317 45898 -16283
rect 45952 -16317 45994 -16283
rect 46977 -16324 47019 -16290
rect 47022 -16324 47030 -16279
rect 44687 -16367 44729 -16333
rect 45280 -16336 45288 -16328
rect 45380 -16336 45388 -16328
rect 44676 -16417 44684 -16406
rect 44687 -16417 44693 -16367
rect 44881 -16410 44923 -16376
rect 44926 -16410 44934 -16365
rect 45026 -16376 45034 -16365
rect 45207 -16370 45277 -16336
rect 45279 -16370 45321 -16336
rect 45391 -16370 45433 -16336
rect 46116 -16360 46158 -16326
rect 46212 -16360 46254 -16326
rect 46308 -16360 46350 -16326
rect 46404 -16360 46446 -16326
rect 46500 -16360 46542 -16326
rect 46596 -16360 46638 -16326
rect 46692 -16360 46734 -16326
rect 45037 -16410 45079 -16376
rect 45670 -16379 45678 -16371
rect 45747 -16379 45753 -16363
rect 45770 -16379 45778 -16371
rect 45781 -16379 45787 -16363
rect 44687 -16451 44729 -16417
rect 44676 -16500 44684 -16489
rect 44687 -16500 44693 -16451
rect 44881 -16494 44923 -16460
rect 44926 -16494 44934 -16449
rect 45026 -16460 45034 -16449
rect 45235 -16453 45277 -16419
rect 45280 -16453 45288 -16408
rect 45380 -16419 45388 -16408
rect 45561 -16413 45603 -16379
rect 45625 -16413 45678 -16379
rect 45705 -16413 45753 -16379
rect 45391 -16453 45433 -16419
rect 45037 -16494 45079 -16460
rect 44687 -16534 44729 -16500
rect 44687 -16568 44693 -16534
rect 43337 -16740 43343 -16706
rect 43633 -16723 43675 -16689
rect 43678 -16723 43686 -16681
rect 41084 -16906 41126 -16872
rect 41156 -16906 41198 -16872
rect 41228 -16906 41270 -16872
rect 41541 -16913 41583 -16879
rect 41586 -16913 41594 -16868
rect 41686 -16879 41694 -16868
rect 41697 -16913 41739 -16879
rect 42281 -16895 42323 -16861
rect 42326 -16895 42334 -16853
rect 40175 -16959 40658 -16925
rect 41509 -16949 41551 -16915
rect 41581 -16949 41623 -16915
rect 41895 -16956 41937 -16922
rect 41940 -16956 41948 -16911
rect 42040 -16922 42048 -16911
rect 42468 -16913 42481 -16845
rect 42509 -16879 42515 -16811
rect 42554 -16843 42560 -16775
rect 42588 -16809 42594 -16743
rect 42598 -16793 42640 -16759
rect 42801 -16838 42843 -16804
rect 42568 -16861 42576 -16853
rect 42579 -16895 42621 -16861
rect 42801 -16906 42843 -16872
rect 42051 -16956 42093 -16922
rect 40175 -16985 40645 -16959
rect 40179 -16993 40387 -16985
rect 40195 -17003 40371 -16993
rect 39921 -17140 40103 -17114
rect 39428 -17174 39470 -17140
rect 39524 -17174 39566 -17140
rect 39620 -17174 39662 -17140
rect 39716 -17174 39758 -17140
rect 39812 -17174 39854 -17140
rect 39908 -17174 40103 -17140
rect 39921 -17200 40103 -17174
rect 40121 -17174 40229 -17050
rect 40380 -17062 40387 -17051
rect 39999 -17870 40041 -17200
rect 40121 -17228 40131 -17174
rect 39806 -17936 39958 -17924
rect 39474 -17970 39958 -17936
rect 39806 -17971 39958 -17970
rect 39987 -17971 40041 -17870
rect 40133 -17971 40175 -17174
rect 40179 -17971 40186 -17174
rect 40391 -17971 40433 -17062
rect 40525 -17971 40567 -16985
rect 40778 -17002 40820 -16968
rect 40874 -17002 40916 -16968
rect 40970 -17002 41012 -16968
rect 41066 -17002 41108 -16968
rect 41162 -17002 41204 -16968
rect 41258 -17002 41300 -16968
rect 41354 -17002 41396 -16968
rect 41863 -16992 41905 -16958
rect 41935 -16992 41977 -16958
rect 42281 -16995 42323 -16961
rect 42326 -16995 42334 -16950
rect 42468 -17001 42476 -16913
rect 42850 -16922 42856 -16788
rect 42568 -16961 42576 -16950
rect 42884 -16956 42890 -16762
rect 42924 -16778 42932 -16767
rect 42920 -16809 42932 -16778
rect 43246 -16796 43288 -16762
rect 42579 -16995 42621 -16961
rect 41516 -17045 41558 -17011
rect 41612 -17045 41654 -17011
rect 41708 -17045 41750 -17011
rect 42217 -17035 42259 -17001
rect 42289 -17035 42331 -17001
rect 42361 -17035 42403 -17001
rect 42433 -17029 42476 -17001
rect 42779 -17025 42821 -16991
rect 42824 -17025 42832 -16980
rect 42920 -16992 42926 -16809
rect 42954 -16995 42960 -16812
rect 42433 -17035 42475 -17029
rect 41870 -17088 41912 -17054
rect 41966 -17088 42008 -17054
rect 42062 -17088 42104 -17054
rect 42966 -17076 42974 -16809
rect 43303 -16812 43304 -16742
rect 43337 -16819 43338 -16740
rect 43820 -16741 43833 -16673
rect 43861 -16707 43867 -16639
rect 43906 -16671 43912 -16603
rect 43940 -16637 43946 -16571
rect 43950 -16621 43992 -16587
rect 44151 -16666 44193 -16632
rect 43920 -16689 43928 -16681
rect 43931 -16723 43973 -16689
rect 44151 -16734 44193 -16700
rect 43820 -16753 43828 -16741
rect 44200 -16750 44206 -16616
rect 43595 -16819 43989 -16753
rect 44234 -16784 44240 -16590
rect 44274 -16606 44282 -16595
rect 44270 -16637 44282 -16606
rect 44596 -16624 44638 -16590
rect 42982 -16860 43024 -16826
rect 43331 -16830 43349 -16819
rect 43331 -16832 43338 -16830
rect 42982 -16928 43024 -16894
rect 43034 -16995 43040 -16860
rect 43265 -16874 43338 -16832
rect 43393 -16874 43989 -16819
rect 44129 -16853 44171 -16819
rect 44174 -16853 44182 -16808
rect 44270 -16820 44276 -16637
rect 44304 -16823 44310 -16640
rect 43265 -16877 43989 -16874
rect 43068 -16980 43074 -16892
rect 43185 -16942 43227 -16908
rect 43230 -16942 43238 -16900
rect 43066 -16991 43074 -16980
rect 43068 -17025 43074 -16991
rect 43077 -17025 43119 -16991
rect 43185 -17042 43227 -17008
rect 43230 -17042 43238 -16997
rect 43078 -17078 43120 -17044
rect 43150 -17078 43192 -17044
rect 43222 -17078 43264 -17044
rect 42224 -17131 42266 -17097
rect 42320 -17131 42362 -17097
rect 42416 -17131 42458 -17097
rect 42512 -17131 42554 -17097
rect 42608 -17131 42650 -17097
rect 43265 -17114 43417 -16877
rect 43595 -16899 43989 -16877
rect 43519 -16925 43989 -16899
rect 44316 -16904 44324 -16637
rect 44653 -16640 44654 -16570
rect 44332 -16688 44374 -16654
rect 44687 -16674 44688 -16568
rect 44881 -16577 44923 -16543
rect 44926 -16577 44934 -16532
rect 45026 -16543 45034 -16532
rect 45235 -16537 45277 -16503
rect 45280 -16537 45288 -16492
rect 45380 -16503 45388 -16492
rect 45625 -16496 45667 -16462
rect 45670 -16496 45678 -16451
rect 45391 -16537 45433 -16503
rect 45037 -16577 45079 -16543
rect 44332 -16756 44374 -16722
rect 44384 -16823 44390 -16688
rect 44946 -16691 44988 -16657
rect 44998 -16718 45004 -16641
rect 44418 -16808 44424 -16720
rect 44535 -16770 44577 -16736
rect 44580 -16770 44588 -16728
rect 44680 -16740 44688 -16729
rect 44691 -16774 44733 -16740
rect 45032 -16752 45038 -16607
rect 45235 -16620 45277 -16586
rect 45280 -16620 45288 -16575
rect 45380 -16586 45388 -16575
rect 45625 -16580 45667 -16546
rect 45670 -16580 45678 -16535
rect 45391 -16620 45433 -16586
rect 45300 -16734 45342 -16700
rect 45352 -16761 45358 -16684
rect 44416 -16819 44424 -16808
rect 44885 -16813 44927 -16779
rect 44930 -16813 44938 -16771
rect 45030 -16779 45038 -16771
rect 45041 -16813 45083 -16779
rect 45386 -16795 45392 -16650
rect 45625 -16663 45667 -16629
rect 45670 -16663 45678 -16618
rect 45747 -16679 45753 -16413
rect 45781 -16413 45823 -16379
rect 45826 -16413 45834 -16371
rect 45770 -16462 45778 -16451
rect 45781 -16462 45787 -16413
rect 45781 -16496 45823 -16462
rect 45826 -16496 45834 -16451
rect 45770 -16546 45778 -16535
rect 45781 -16546 45787 -16496
rect 45781 -16580 45823 -16546
rect 45826 -16580 45834 -16535
rect 45770 -16629 45778 -16618
rect 45781 -16629 45787 -16580
rect 45781 -16663 45823 -16629
rect 45826 -16663 45834 -16618
rect 45770 -16697 45778 -16671
rect 45781 -16713 45787 -16663
rect 45690 -16777 45732 -16743
rect 45747 -16804 45748 -16727
rect 45781 -16809 45782 -16713
rect 44418 -16853 44424 -16819
rect 44427 -16853 44469 -16819
rect 44535 -16870 44577 -16836
rect 44580 -16870 44588 -16825
rect 44680 -16832 44688 -16821
rect 44691 -16866 44733 -16832
rect 45239 -16856 45281 -16822
rect 45284 -16856 45292 -16814
rect 45384 -16822 45392 -16814
rect 45395 -16856 45437 -16822
rect 45812 -16845 45820 -16697
rect 45835 -16713 45839 -16363
rect 45869 -16679 45873 -16363
rect 45926 -16379 45934 -16371
rect 45875 -16413 45917 -16379
rect 45937 -16413 45989 -16379
rect 46647 -16422 46653 -16406
rect 46670 -16422 46678 -16414
rect 46681 -16422 46687 -16406
rect 46977 -16408 47019 -16374
rect 47022 -16408 47030 -16363
rect 45926 -16462 45934 -16451
rect 46107 -16456 46149 -16422
rect 46179 -16456 46221 -16422
rect 46251 -16456 46293 -16422
rect 46395 -16456 46437 -16422
rect 46467 -16456 46581 -16422
rect 46611 -16456 46653 -16422
rect 45937 -16496 45979 -16462
rect 45926 -16546 45934 -16535
rect 46504 -16539 46546 -16505
rect 45937 -16580 45979 -16546
rect 45926 -16629 45934 -16618
rect 45937 -16663 45979 -16629
rect 46169 -16689 46211 -16655
rect 46214 -16689 46222 -16644
rect 46291 -16706 46297 -16588
rect 46314 -16655 46322 -16644
rect 46325 -16655 46331 -16622
rect 46361 -16655 46367 -16622
rect 46325 -16689 46367 -16655
rect 46370 -16689 46378 -16644
rect 46325 -16740 46331 -16689
rect 46361 -16740 46367 -16689
rect 46395 -16706 46401 -16589
rect 46492 -16630 46493 -16589
rect 46504 -16623 46546 -16589
rect 46504 -16706 46546 -16672
rect 46647 -16706 46653 -16456
rect 46681 -16456 46723 -16422
rect 46670 -16505 46678 -16494
rect 46681 -16505 46687 -16456
rect 46977 -16491 47019 -16457
rect 47022 -16491 47030 -16446
rect 46681 -16539 46723 -16505
rect 46670 -16589 46678 -16578
rect 46681 -16589 46687 -16539
rect 46831 -16565 46939 -16499
rect 47099 -16507 47105 -16241
rect 47133 -16241 47175 -16207
rect 47178 -16241 47186 -16199
rect 47122 -16290 47130 -16279
rect 47133 -16290 47139 -16241
rect 47133 -16324 47175 -16290
rect 47178 -16324 47186 -16279
rect 47122 -16374 47130 -16363
rect 47133 -16374 47139 -16324
rect 47133 -16408 47175 -16374
rect 47178 -16408 47186 -16363
rect 47122 -16457 47130 -16446
rect 47133 -16457 47139 -16408
rect 47133 -16491 47175 -16457
rect 47178 -16491 47186 -16446
rect 47122 -16525 47130 -16499
rect 47133 -16541 47139 -16491
rect 46681 -16623 46723 -16589
rect 47042 -16605 47084 -16571
rect 46670 -16672 46678 -16661
rect 46681 -16672 46687 -16623
rect 47099 -16632 47100 -16555
rect 47133 -16637 47134 -16541
rect 46681 -16706 46723 -16672
rect 47164 -16673 47172 -16525
rect 47187 -16541 47191 -16191
rect 47221 -16507 47225 -16191
rect 47278 -16207 47286 -16199
rect 47227 -16241 47269 -16207
rect 47289 -16241 47341 -16207
rect 48204 -16231 48246 -16197
rect 48300 -16231 48342 -16197
rect 48396 -16231 48438 -16197
rect 50366 -16207 50374 -16199
rect 50443 -16207 50449 -16191
rect 50466 -16207 50474 -16199
rect 50477 -16207 50483 -16191
rect 47997 -16250 48003 -16234
rect 48020 -16250 48028 -16242
rect 48031 -16250 48037 -16234
rect 47278 -16290 47286 -16279
rect 47457 -16284 47499 -16250
rect 47529 -16284 47571 -16250
rect 47601 -16284 47643 -16250
rect 47745 -16284 47787 -16250
rect 47817 -16284 47931 -16250
rect 47961 -16284 48003 -16250
rect 47289 -16324 47331 -16290
rect 47278 -16374 47286 -16363
rect 47854 -16367 47896 -16333
rect 47289 -16408 47331 -16374
rect 47278 -16457 47286 -16446
rect 47289 -16491 47331 -16457
rect 47519 -16517 47561 -16483
rect 47564 -16517 47572 -16472
rect 47641 -16534 47647 -16416
rect 47664 -16483 47672 -16472
rect 47675 -16483 47681 -16450
rect 47711 -16483 47717 -16450
rect 47675 -16517 47717 -16483
rect 47720 -16517 47728 -16472
rect 47675 -16568 47681 -16517
rect 47711 -16568 47717 -16517
rect 47745 -16534 47751 -16417
rect 47842 -16458 47843 -16417
rect 47854 -16451 47896 -16417
rect 47854 -16534 47896 -16500
rect 47997 -16534 48003 -16284
rect 48031 -16284 48073 -16250
rect 48558 -16274 48600 -16240
rect 48654 -16274 48696 -16240
rect 48750 -16274 48792 -16240
rect 50257 -16241 50299 -16207
rect 50321 -16241 50374 -16207
rect 50401 -16241 50449 -16207
rect 48020 -16333 48028 -16322
rect 48031 -16333 48037 -16284
rect 48270 -16293 48278 -16285
rect 48370 -16293 48378 -16285
rect 48197 -16327 48267 -16293
rect 48269 -16327 48311 -16293
rect 48381 -16327 48423 -16293
rect 48912 -16317 48954 -16283
rect 49008 -16317 49050 -16283
rect 49104 -16317 49146 -16283
rect 49200 -16317 49242 -16283
rect 49296 -16317 49338 -16283
rect 50321 -16324 50363 -16290
rect 50366 -16324 50374 -16279
rect 48031 -16367 48073 -16333
rect 48624 -16336 48632 -16328
rect 48724 -16336 48732 -16328
rect 48020 -16417 48028 -16406
rect 48031 -16417 48037 -16367
rect 48225 -16410 48267 -16376
rect 48270 -16410 48278 -16365
rect 48370 -16376 48378 -16365
rect 48551 -16370 48621 -16336
rect 48623 -16370 48665 -16336
rect 48735 -16370 48777 -16336
rect 49460 -16360 49502 -16326
rect 49556 -16360 49598 -16326
rect 49652 -16360 49694 -16326
rect 49748 -16360 49790 -16326
rect 49844 -16360 49886 -16326
rect 49940 -16360 49982 -16326
rect 50036 -16360 50078 -16326
rect 48381 -16410 48423 -16376
rect 49014 -16379 49022 -16371
rect 49091 -16379 49097 -16363
rect 49114 -16379 49122 -16371
rect 49125 -16379 49131 -16363
rect 48031 -16451 48073 -16417
rect 48020 -16500 48028 -16489
rect 48031 -16500 48037 -16451
rect 48225 -16494 48267 -16460
rect 48270 -16494 48278 -16449
rect 48370 -16460 48378 -16449
rect 48579 -16453 48621 -16419
rect 48624 -16453 48632 -16408
rect 48724 -16419 48732 -16408
rect 48905 -16413 48947 -16379
rect 48969 -16413 49022 -16379
rect 49049 -16413 49097 -16379
rect 48735 -16453 48777 -16419
rect 48381 -16494 48423 -16460
rect 48031 -16534 48073 -16500
rect 48031 -16568 48037 -16534
rect 46681 -16740 46687 -16706
rect 46977 -16723 47019 -16689
rect 47022 -16723 47030 -16681
rect 44428 -16906 44470 -16872
rect 44500 -16906 44542 -16872
rect 44572 -16906 44614 -16872
rect 44885 -16913 44927 -16879
rect 44930 -16913 44938 -16868
rect 45030 -16879 45038 -16868
rect 45041 -16913 45083 -16879
rect 45625 -16895 45667 -16861
rect 45670 -16895 45678 -16853
rect 43519 -16959 44002 -16925
rect 44853 -16949 44895 -16915
rect 44925 -16949 44967 -16915
rect 45239 -16956 45281 -16922
rect 45284 -16956 45292 -16911
rect 45384 -16922 45392 -16911
rect 45812 -16913 45825 -16845
rect 45853 -16879 45859 -16811
rect 45898 -16843 45904 -16775
rect 45932 -16809 45938 -16743
rect 45942 -16793 45984 -16759
rect 46145 -16838 46187 -16804
rect 45912 -16861 45920 -16853
rect 45923 -16895 45965 -16861
rect 46145 -16906 46187 -16872
rect 45395 -16956 45437 -16922
rect 43519 -16985 43989 -16959
rect 43523 -16993 43731 -16985
rect 43539 -17003 43715 -16993
rect 43265 -17140 43447 -17114
rect 42772 -17174 42814 -17140
rect 42868 -17174 42910 -17140
rect 42964 -17174 43006 -17140
rect 43060 -17174 43102 -17140
rect 43156 -17174 43198 -17140
rect 43252 -17174 43447 -17140
rect 43265 -17200 43447 -17174
rect 43465 -17174 43573 -17050
rect 43724 -17062 43731 -17051
rect 43343 -17870 43385 -17200
rect 43465 -17228 43475 -17174
rect 43150 -17936 43302 -17924
rect 42818 -17970 43302 -17936
rect 43150 -17971 43302 -17970
rect 43331 -17971 43385 -17870
rect 43477 -17971 43519 -17174
rect 43523 -17971 43530 -17174
rect 43735 -17971 43777 -17062
rect 43869 -17971 43911 -16985
rect 44122 -17002 44164 -16968
rect 44218 -17002 44260 -16968
rect 44314 -17002 44356 -16968
rect 44410 -17002 44452 -16968
rect 44506 -17002 44548 -16968
rect 44602 -17002 44644 -16968
rect 44698 -17002 44740 -16968
rect 45207 -16992 45249 -16958
rect 45279 -16992 45321 -16958
rect 45625 -16995 45667 -16961
rect 45670 -16995 45678 -16950
rect 45812 -17001 45820 -16913
rect 46194 -16922 46200 -16788
rect 45912 -16961 45920 -16950
rect 46228 -16956 46234 -16762
rect 46268 -16778 46276 -16767
rect 46264 -16809 46276 -16778
rect 46590 -16796 46632 -16762
rect 45923 -16995 45965 -16961
rect 44860 -17045 44902 -17011
rect 44956 -17045 44998 -17011
rect 45052 -17045 45094 -17011
rect 45561 -17035 45603 -17001
rect 45633 -17035 45675 -17001
rect 45705 -17035 45747 -17001
rect 45777 -17029 45820 -17001
rect 46123 -17025 46165 -16991
rect 46168 -17025 46176 -16980
rect 46264 -16992 46270 -16809
rect 46298 -16995 46304 -16812
rect 45777 -17035 45819 -17029
rect 45214 -17088 45256 -17054
rect 45310 -17088 45352 -17054
rect 45406 -17088 45448 -17054
rect 46310 -17076 46318 -16809
rect 46647 -16812 46648 -16742
rect 46681 -16819 46682 -16740
rect 47164 -16741 47177 -16673
rect 47205 -16707 47211 -16639
rect 47250 -16671 47256 -16603
rect 47284 -16637 47290 -16571
rect 47294 -16621 47336 -16587
rect 47495 -16666 47537 -16632
rect 47264 -16689 47272 -16681
rect 47275 -16723 47317 -16689
rect 47495 -16734 47537 -16700
rect 47164 -16753 47172 -16741
rect 47544 -16750 47550 -16616
rect 46939 -16819 47333 -16753
rect 47578 -16784 47584 -16590
rect 47618 -16606 47626 -16595
rect 47614 -16637 47626 -16606
rect 47940 -16624 47982 -16590
rect 46326 -16860 46368 -16826
rect 46675 -16830 46693 -16819
rect 46675 -16832 46682 -16830
rect 46326 -16928 46368 -16894
rect 46378 -16995 46384 -16860
rect 46609 -16874 46682 -16832
rect 46737 -16874 47333 -16819
rect 47473 -16853 47515 -16819
rect 47518 -16853 47526 -16808
rect 47614 -16820 47620 -16637
rect 47648 -16823 47654 -16640
rect 46609 -16877 47333 -16874
rect 46412 -16980 46418 -16892
rect 46529 -16942 46571 -16908
rect 46574 -16942 46582 -16900
rect 46410 -16991 46418 -16980
rect 46412 -17025 46418 -16991
rect 46421 -17025 46463 -16991
rect 46529 -17042 46571 -17008
rect 46574 -17042 46582 -16997
rect 46422 -17078 46464 -17044
rect 46494 -17078 46536 -17044
rect 46566 -17078 46608 -17044
rect 45568 -17131 45610 -17097
rect 45664 -17131 45706 -17097
rect 45760 -17131 45802 -17097
rect 45856 -17131 45898 -17097
rect 45952 -17131 45994 -17097
rect 46609 -17114 46761 -16877
rect 46939 -16899 47333 -16877
rect 46863 -16925 47333 -16899
rect 47660 -16904 47668 -16637
rect 47997 -16640 47998 -16570
rect 47676 -16688 47718 -16654
rect 48031 -16674 48032 -16568
rect 48225 -16577 48267 -16543
rect 48270 -16577 48278 -16532
rect 48370 -16543 48378 -16532
rect 48579 -16537 48621 -16503
rect 48624 -16537 48632 -16492
rect 48724 -16503 48732 -16492
rect 48969 -16496 49011 -16462
rect 49014 -16496 49022 -16451
rect 48735 -16537 48777 -16503
rect 48381 -16577 48423 -16543
rect 47676 -16756 47718 -16722
rect 47728 -16823 47734 -16688
rect 48290 -16691 48332 -16657
rect 48342 -16718 48348 -16641
rect 47762 -16808 47768 -16720
rect 47879 -16770 47921 -16736
rect 47924 -16770 47932 -16728
rect 48024 -16740 48032 -16729
rect 48035 -16774 48077 -16740
rect 48376 -16752 48382 -16607
rect 48579 -16620 48621 -16586
rect 48624 -16620 48632 -16575
rect 48724 -16586 48732 -16575
rect 48969 -16580 49011 -16546
rect 49014 -16580 49022 -16535
rect 48735 -16620 48777 -16586
rect 48644 -16734 48686 -16700
rect 48696 -16761 48702 -16684
rect 47760 -16819 47768 -16808
rect 48229 -16813 48271 -16779
rect 48274 -16813 48282 -16771
rect 48374 -16779 48382 -16771
rect 48385 -16813 48427 -16779
rect 48730 -16795 48736 -16650
rect 48969 -16663 49011 -16629
rect 49014 -16663 49022 -16618
rect 49091 -16679 49097 -16413
rect 49125 -16413 49167 -16379
rect 49170 -16413 49178 -16371
rect 49114 -16462 49122 -16451
rect 49125 -16462 49131 -16413
rect 49125 -16496 49167 -16462
rect 49170 -16496 49178 -16451
rect 49114 -16546 49122 -16535
rect 49125 -16546 49131 -16496
rect 49125 -16580 49167 -16546
rect 49170 -16580 49178 -16535
rect 49114 -16629 49122 -16618
rect 49125 -16629 49131 -16580
rect 49125 -16663 49167 -16629
rect 49170 -16663 49178 -16618
rect 49114 -16697 49122 -16671
rect 49125 -16713 49131 -16663
rect 49034 -16777 49076 -16743
rect 49091 -16804 49092 -16727
rect 49125 -16809 49126 -16713
rect 47762 -16853 47768 -16819
rect 47771 -16853 47813 -16819
rect 47879 -16870 47921 -16836
rect 47924 -16870 47932 -16825
rect 48024 -16832 48032 -16821
rect 48035 -16866 48077 -16832
rect 48583 -16856 48625 -16822
rect 48628 -16856 48636 -16814
rect 48728 -16822 48736 -16814
rect 48739 -16856 48781 -16822
rect 49156 -16845 49164 -16697
rect 49179 -16713 49183 -16363
rect 49213 -16679 49217 -16363
rect 49270 -16379 49278 -16371
rect 49219 -16413 49261 -16379
rect 49281 -16413 49333 -16379
rect 49991 -16422 49997 -16406
rect 50014 -16422 50022 -16414
rect 50025 -16422 50031 -16406
rect 50321 -16408 50363 -16374
rect 50366 -16408 50374 -16363
rect 49270 -16462 49278 -16451
rect 49451 -16456 49493 -16422
rect 49523 -16456 49565 -16422
rect 49595 -16456 49637 -16422
rect 49739 -16456 49781 -16422
rect 49811 -16456 49925 -16422
rect 49955 -16456 49997 -16422
rect 49281 -16496 49323 -16462
rect 49270 -16546 49278 -16535
rect 49848 -16539 49890 -16505
rect 49281 -16580 49323 -16546
rect 49270 -16629 49278 -16618
rect 49281 -16663 49323 -16629
rect 49513 -16689 49555 -16655
rect 49558 -16689 49566 -16644
rect 49635 -16706 49641 -16588
rect 49658 -16655 49666 -16644
rect 49669 -16655 49675 -16622
rect 49705 -16655 49711 -16622
rect 49669 -16689 49711 -16655
rect 49714 -16689 49722 -16644
rect 49669 -16740 49675 -16689
rect 49705 -16740 49711 -16689
rect 49739 -16706 49745 -16589
rect 49836 -16630 49837 -16589
rect 49848 -16623 49890 -16589
rect 49848 -16706 49890 -16672
rect 49991 -16706 49997 -16456
rect 50025 -16456 50067 -16422
rect 50014 -16505 50022 -16494
rect 50025 -16505 50031 -16456
rect 50321 -16491 50363 -16457
rect 50366 -16491 50374 -16446
rect 50025 -16539 50067 -16505
rect 50014 -16589 50022 -16578
rect 50025 -16589 50031 -16539
rect 50175 -16565 50283 -16499
rect 50443 -16507 50449 -16241
rect 50477 -16241 50519 -16207
rect 50522 -16241 50530 -16199
rect 50466 -16290 50474 -16279
rect 50477 -16290 50483 -16241
rect 50477 -16324 50519 -16290
rect 50522 -16324 50530 -16279
rect 50466 -16374 50474 -16363
rect 50477 -16374 50483 -16324
rect 50477 -16408 50519 -16374
rect 50522 -16408 50530 -16363
rect 50466 -16457 50474 -16446
rect 50477 -16457 50483 -16408
rect 50477 -16491 50519 -16457
rect 50522 -16491 50530 -16446
rect 50466 -16525 50474 -16499
rect 50477 -16541 50483 -16491
rect 50025 -16623 50067 -16589
rect 50386 -16605 50428 -16571
rect 50014 -16672 50022 -16661
rect 50025 -16672 50031 -16623
rect 50443 -16632 50444 -16555
rect 50477 -16637 50478 -16541
rect 50025 -16706 50067 -16672
rect 50508 -16673 50516 -16525
rect 50531 -16541 50535 -16191
rect 50565 -16507 50569 -16191
rect 50622 -16207 50630 -16199
rect 50571 -16241 50613 -16207
rect 50633 -16241 50685 -16207
rect 51548 -16231 51590 -16197
rect 51644 -16231 51686 -16197
rect 51740 -16231 51782 -16197
rect 53711 -16207 53718 -16199
rect 51341 -16250 51347 -16234
rect 51364 -16250 51372 -16242
rect 51375 -16250 51381 -16234
rect 50622 -16290 50630 -16279
rect 50801 -16284 50843 -16250
rect 50873 -16284 50915 -16250
rect 50945 -16284 50987 -16250
rect 51089 -16284 51131 -16250
rect 51161 -16284 51275 -16250
rect 51305 -16284 51347 -16250
rect 50633 -16324 50675 -16290
rect 50622 -16374 50630 -16363
rect 51198 -16367 51240 -16333
rect 50633 -16408 50675 -16374
rect 50622 -16457 50630 -16446
rect 50633 -16491 50675 -16457
rect 50863 -16517 50905 -16483
rect 50908 -16517 50916 -16472
rect 50985 -16534 50991 -16416
rect 51008 -16483 51016 -16472
rect 51019 -16483 51025 -16450
rect 51055 -16483 51061 -16450
rect 51019 -16517 51061 -16483
rect 51064 -16517 51072 -16472
rect 51019 -16568 51025 -16517
rect 51055 -16568 51061 -16517
rect 51089 -16534 51095 -16417
rect 51186 -16458 51187 -16417
rect 51198 -16451 51240 -16417
rect 51198 -16534 51240 -16500
rect 51341 -16534 51347 -16284
rect 51375 -16284 51417 -16250
rect 51902 -16274 51944 -16240
rect 51998 -16274 52040 -16240
rect 52094 -16274 52136 -16240
rect 53602 -16241 53643 -16207
rect 53666 -16241 53718 -16207
rect 53746 -16241 53787 -16207
rect 51364 -16333 51372 -16322
rect 51375 -16333 51381 -16284
rect 51614 -16293 51622 -16285
rect 51714 -16293 51722 -16285
rect 51541 -16327 51611 -16293
rect 51613 -16327 51655 -16293
rect 51725 -16327 51767 -16293
rect 52256 -16317 52298 -16283
rect 52352 -16317 52394 -16283
rect 52448 -16317 52490 -16283
rect 52544 -16317 52586 -16283
rect 52640 -16317 52682 -16283
rect 53666 -16324 53707 -16290
rect 53711 -16324 53718 -16279
rect 51375 -16367 51417 -16333
rect 51968 -16336 51976 -16328
rect 52068 -16336 52076 -16328
rect 51364 -16417 51372 -16406
rect 51375 -16417 51381 -16367
rect 51569 -16410 51611 -16376
rect 51614 -16410 51622 -16365
rect 51714 -16376 51722 -16365
rect 51895 -16370 51965 -16336
rect 51967 -16370 52009 -16336
rect 52079 -16370 52121 -16336
rect 52804 -16360 52846 -16326
rect 52900 -16360 52942 -16326
rect 52996 -16360 53038 -16326
rect 53092 -16360 53134 -16326
rect 53188 -16360 53230 -16326
rect 53284 -16360 53326 -16326
rect 53380 -16360 53422 -16326
rect 51725 -16410 51767 -16376
rect 52358 -16379 52366 -16371
rect 52435 -16379 52441 -16363
rect 52458 -16379 52466 -16371
rect 52469 -16379 52475 -16363
rect 51375 -16451 51417 -16417
rect 51364 -16500 51372 -16489
rect 51375 -16500 51381 -16451
rect 51569 -16494 51611 -16460
rect 51614 -16494 51622 -16449
rect 51714 -16460 51722 -16449
rect 51923 -16453 51965 -16419
rect 51968 -16453 51976 -16408
rect 52068 -16419 52076 -16408
rect 52249 -16413 52291 -16379
rect 52313 -16413 52366 -16379
rect 52393 -16413 52441 -16379
rect 52079 -16453 52121 -16419
rect 51725 -16494 51767 -16460
rect 51375 -16534 51417 -16500
rect 51375 -16568 51381 -16534
rect 50025 -16740 50031 -16706
rect 50321 -16723 50363 -16689
rect 50366 -16723 50374 -16681
rect 47772 -16906 47814 -16872
rect 47844 -16906 47886 -16872
rect 47916 -16906 47958 -16872
rect 48229 -16913 48271 -16879
rect 48274 -16913 48282 -16868
rect 48374 -16879 48382 -16868
rect 48385 -16913 48427 -16879
rect 48969 -16895 49011 -16861
rect 49014 -16895 49022 -16853
rect 46863 -16959 47346 -16925
rect 48197 -16949 48239 -16915
rect 48269 -16949 48311 -16915
rect 48583 -16956 48625 -16922
rect 48628 -16956 48636 -16911
rect 48728 -16922 48736 -16911
rect 49156 -16913 49169 -16845
rect 49197 -16879 49203 -16811
rect 49242 -16843 49248 -16775
rect 49276 -16809 49282 -16743
rect 49286 -16793 49328 -16759
rect 49489 -16838 49531 -16804
rect 49256 -16861 49264 -16853
rect 49267 -16895 49309 -16861
rect 49489 -16906 49531 -16872
rect 48739 -16956 48781 -16922
rect 46863 -16985 47333 -16959
rect 46867 -16993 47075 -16985
rect 46883 -17003 47059 -16993
rect 46609 -17140 46791 -17114
rect 46116 -17174 46158 -17140
rect 46212 -17174 46254 -17140
rect 46308 -17174 46350 -17140
rect 46404 -17174 46446 -17140
rect 46500 -17174 46542 -17140
rect 46596 -17174 46791 -17140
rect 46609 -17200 46791 -17174
rect 46809 -17174 46917 -17050
rect 47068 -17062 47075 -17051
rect 46687 -17870 46729 -17200
rect 46809 -17228 46819 -17174
rect 46494 -17936 46646 -17924
rect 46162 -17970 46646 -17936
rect 46494 -17971 46646 -17970
rect 46675 -17971 46729 -17870
rect 46821 -17971 46863 -17174
rect 46867 -17971 46874 -17174
rect 47079 -17971 47121 -17062
rect 47213 -17971 47255 -16985
rect 47466 -17002 47508 -16968
rect 47562 -17002 47604 -16968
rect 47658 -17002 47700 -16968
rect 47754 -17002 47796 -16968
rect 47850 -17002 47892 -16968
rect 47946 -17002 47988 -16968
rect 48042 -17002 48084 -16968
rect 48551 -16992 48593 -16958
rect 48623 -16992 48665 -16958
rect 48969 -16995 49011 -16961
rect 49014 -16995 49022 -16950
rect 49156 -17001 49164 -16913
rect 49538 -16922 49544 -16788
rect 49256 -16961 49264 -16950
rect 49572 -16956 49578 -16762
rect 49612 -16778 49620 -16767
rect 49608 -16809 49620 -16778
rect 49934 -16796 49976 -16762
rect 49267 -16995 49309 -16961
rect 48204 -17045 48246 -17011
rect 48300 -17045 48342 -17011
rect 48396 -17045 48438 -17011
rect 48905 -17035 48947 -17001
rect 48977 -17035 49019 -17001
rect 49049 -17035 49091 -17001
rect 49121 -17029 49164 -17001
rect 49467 -17025 49509 -16991
rect 49512 -17025 49520 -16980
rect 49608 -16992 49614 -16809
rect 49642 -16995 49648 -16812
rect 49121 -17035 49163 -17029
rect 48558 -17088 48600 -17054
rect 48654 -17088 48696 -17054
rect 48750 -17088 48792 -17054
rect 49654 -17076 49662 -16809
rect 49991 -16812 49992 -16742
rect 50025 -16819 50026 -16740
rect 50508 -16741 50521 -16673
rect 50549 -16707 50555 -16639
rect 50594 -16671 50600 -16603
rect 50628 -16637 50634 -16571
rect 50638 -16621 50680 -16587
rect 50839 -16666 50881 -16632
rect 50608 -16689 50616 -16681
rect 50619 -16723 50661 -16689
rect 50839 -16734 50881 -16700
rect 50508 -16753 50516 -16741
rect 50888 -16750 50894 -16616
rect 50283 -16819 50677 -16753
rect 50922 -16784 50928 -16590
rect 50962 -16606 50970 -16595
rect 50958 -16637 50970 -16606
rect 51284 -16624 51326 -16590
rect 49670 -16860 49712 -16826
rect 50019 -16830 50037 -16819
rect 50019 -16832 50026 -16830
rect 49670 -16928 49712 -16894
rect 49722 -16995 49728 -16860
rect 49953 -16874 50026 -16832
rect 50081 -16874 50677 -16819
rect 50817 -16853 50859 -16819
rect 50862 -16853 50870 -16808
rect 50958 -16820 50964 -16637
rect 50992 -16823 50998 -16640
rect 49953 -16877 50677 -16874
rect 49756 -16980 49762 -16892
rect 49873 -16942 49915 -16908
rect 49918 -16942 49926 -16900
rect 49754 -16991 49762 -16980
rect 49756 -17025 49762 -16991
rect 49765 -17025 49807 -16991
rect 49873 -17042 49915 -17008
rect 49918 -17042 49926 -16997
rect 49766 -17078 49808 -17044
rect 49838 -17078 49880 -17044
rect 49910 -17078 49952 -17044
rect 48912 -17131 48954 -17097
rect 49008 -17131 49050 -17097
rect 49104 -17131 49146 -17097
rect 49200 -17131 49242 -17097
rect 49296 -17131 49338 -17097
rect 49953 -17114 50105 -16877
rect 50283 -16899 50677 -16877
rect 50207 -16925 50677 -16899
rect 51004 -16904 51012 -16637
rect 51341 -16640 51342 -16570
rect 51020 -16688 51062 -16654
rect 51375 -16674 51376 -16568
rect 51569 -16577 51611 -16543
rect 51614 -16577 51622 -16532
rect 51714 -16543 51722 -16532
rect 51923 -16537 51965 -16503
rect 51968 -16537 51976 -16492
rect 52068 -16503 52076 -16492
rect 52313 -16496 52355 -16462
rect 52358 -16496 52366 -16451
rect 52079 -16537 52121 -16503
rect 51725 -16577 51767 -16543
rect 51020 -16756 51062 -16722
rect 51072 -16823 51078 -16688
rect 51634 -16691 51676 -16657
rect 51686 -16718 51692 -16641
rect 51106 -16808 51112 -16720
rect 51223 -16770 51265 -16736
rect 51268 -16770 51276 -16728
rect 51368 -16740 51376 -16729
rect 51379 -16774 51421 -16740
rect 51720 -16752 51726 -16607
rect 51923 -16620 51965 -16586
rect 51968 -16620 51976 -16575
rect 52068 -16586 52076 -16575
rect 52313 -16580 52355 -16546
rect 52358 -16580 52366 -16535
rect 52079 -16620 52121 -16586
rect 51988 -16734 52030 -16700
rect 52040 -16761 52046 -16684
rect 51104 -16819 51112 -16808
rect 51573 -16813 51615 -16779
rect 51618 -16813 51626 -16771
rect 51718 -16779 51726 -16771
rect 51729 -16813 51771 -16779
rect 52074 -16795 52080 -16650
rect 52313 -16663 52355 -16629
rect 52358 -16663 52366 -16618
rect 52435 -16679 52441 -16413
rect 52469 -16413 52511 -16379
rect 52514 -16413 52522 -16371
rect 52458 -16462 52466 -16451
rect 52469 -16462 52475 -16413
rect 52469 -16496 52511 -16462
rect 52514 -16496 52522 -16451
rect 52458 -16546 52466 -16535
rect 52469 -16546 52475 -16496
rect 52469 -16580 52511 -16546
rect 52514 -16580 52522 -16535
rect 52458 -16629 52466 -16618
rect 52469 -16629 52475 -16580
rect 52469 -16663 52511 -16629
rect 52514 -16663 52522 -16618
rect 52458 -16697 52466 -16671
rect 52469 -16713 52475 -16663
rect 52378 -16777 52420 -16743
rect 52435 -16804 52436 -16727
rect 52469 -16809 52470 -16713
rect 51106 -16853 51112 -16819
rect 51115 -16853 51157 -16819
rect 51223 -16870 51265 -16836
rect 51268 -16870 51276 -16825
rect 51368 -16832 51376 -16821
rect 51379 -16866 51421 -16832
rect 51927 -16856 51969 -16822
rect 51972 -16856 51980 -16814
rect 52072 -16822 52080 -16814
rect 52083 -16856 52125 -16822
rect 52500 -16845 52508 -16697
rect 52523 -16713 52527 -16363
rect 52557 -16679 52561 -16363
rect 52614 -16379 52622 -16371
rect 52563 -16413 52605 -16379
rect 52625 -16413 52677 -16379
rect 53335 -16422 53341 -16406
rect 53358 -16422 53366 -16414
rect 53369 -16422 53375 -16406
rect 53666 -16408 53707 -16374
rect 53711 -16408 53718 -16363
rect 52614 -16462 52622 -16451
rect 52795 -16456 52837 -16422
rect 52867 -16456 52909 -16422
rect 52939 -16456 52981 -16422
rect 53083 -16456 53125 -16422
rect 53155 -16456 53269 -16422
rect 53299 -16456 53341 -16422
rect 52625 -16496 52667 -16462
rect 52614 -16546 52622 -16535
rect 53192 -16539 53234 -16505
rect 52625 -16580 52667 -16546
rect 52614 -16629 52622 -16618
rect 52625 -16663 52667 -16629
rect 52857 -16689 52899 -16655
rect 52902 -16689 52910 -16644
rect 52979 -16706 52985 -16588
rect 53002 -16655 53010 -16644
rect 53013 -16655 53019 -16622
rect 53049 -16655 53055 -16622
rect 53013 -16689 53055 -16655
rect 53058 -16689 53066 -16644
rect 53013 -16740 53019 -16689
rect 53049 -16740 53055 -16689
rect 53083 -16706 53089 -16589
rect 53180 -16630 53181 -16589
rect 53192 -16623 53234 -16589
rect 53192 -16706 53234 -16672
rect 53335 -16706 53341 -16456
rect 53369 -16456 53411 -16422
rect 53358 -16505 53366 -16494
rect 53369 -16505 53375 -16456
rect 53666 -16491 53707 -16457
rect 53711 -16491 53718 -16446
rect 53369 -16539 53411 -16505
rect 53358 -16589 53366 -16578
rect 53369 -16589 53375 -16539
rect 53519 -16565 53628 -16499
rect 53788 -16507 53793 -16191
rect 53811 -16207 53818 -16199
rect 53822 -16207 53827 -16191
rect 53822 -16241 53863 -16207
rect 53867 -16241 53874 -16199
rect 53811 -16290 53818 -16279
rect 53822 -16290 53827 -16241
rect 53822 -16324 53863 -16290
rect 53867 -16324 53874 -16279
rect 53811 -16374 53818 -16363
rect 53822 -16374 53827 -16324
rect 53822 -16408 53863 -16374
rect 53867 -16408 53874 -16363
rect 53811 -16457 53818 -16446
rect 53822 -16457 53827 -16408
rect 53822 -16491 53863 -16457
rect 53867 -16491 53874 -16446
rect 53811 -16525 53818 -16499
rect 53822 -16541 53827 -16491
rect 53369 -16623 53411 -16589
rect 53731 -16605 53772 -16571
rect 53358 -16672 53366 -16661
rect 53369 -16672 53375 -16623
rect 53369 -16706 53411 -16672
rect 53853 -16673 53860 -16525
rect 53876 -16541 53879 -16191
rect 53910 -16507 53913 -16191
rect 53967 -16207 53974 -16199
rect 53916 -16241 53957 -16207
rect 53978 -16241 54029 -16207
rect 54893 -16231 54934 -16197
rect 54989 -16231 55030 -16197
rect 55085 -16231 55126 -16197
rect 57055 -16207 57062 -16199
rect 54686 -16250 54691 -16234
rect 54709 -16250 54716 -16242
rect 54720 -16250 54725 -16234
rect 53967 -16290 53974 -16279
rect 54146 -16284 54187 -16250
rect 54218 -16284 54259 -16250
rect 54290 -16284 54331 -16250
rect 54434 -16284 54475 -16250
rect 54506 -16284 54619 -16250
rect 54650 -16284 54691 -16250
rect 53978 -16324 54019 -16290
rect 53967 -16374 53974 -16363
rect 54543 -16367 54584 -16333
rect 53978 -16408 54019 -16374
rect 53967 -16457 53974 -16446
rect 53978 -16491 54019 -16457
rect 54208 -16517 54249 -16483
rect 54253 -16517 54260 -16472
rect 54330 -16534 54335 -16416
rect 54353 -16483 54360 -16472
rect 54364 -16483 54369 -16450
rect 54400 -16483 54405 -16450
rect 54364 -16517 54405 -16483
rect 54409 -16517 54416 -16472
rect 54364 -16568 54369 -16517
rect 54400 -16568 54405 -16517
rect 54434 -16534 54439 -16417
rect 54543 -16451 54584 -16417
rect 54543 -16534 54584 -16500
rect 54686 -16534 54691 -16284
rect 54720 -16284 54761 -16250
rect 55247 -16274 55288 -16240
rect 55343 -16274 55384 -16240
rect 55439 -16274 55480 -16240
rect 56946 -16241 56987 -16207
rect 57010 -16241 57062 -16207
rect 57090 -16241 57131 -16207
rect 54709 -16333 54716 -16322
rect 54720 -16333 54725 -16284
rect 54959 -16293 54966 -16285
rect 55059 -16293 55066 -16285
rect 54886 -16327 54955 -16293
rect 54958 -16327 54999 -16293
rect 55070 -16327 55111 -16293
rect 55601 -16317 55642 -16283
rect 55697 -16317 55738 -16283
rect 55793 -16317 55834 -16283
rect 55889 -16317 55930 -16283
rect 55985 -16317 56026 -16283
rect 57010 -16324 57051 -16290
rect 57055 -16324 57062 -16279
rect 54720 -16367 54761 -16333
rect 55313 -16336 55320 -16328
rect 55413 -16336 55420 -16328
rect 54709 -16417 54716 -16406
rect 54720 -16417 54725 -16367
rect 54914 -16410 54955 -16376
rect 54959 -16410 54966 -16365
rect 55059 -16376 55066 -16365
rect 55240 -16370 55309 -16336
rect 55312 -16370 55353 -16336
rect 55424 -16370 55465 -16336
rect 56149 -16360 56190 -16326
rect 56245 -16360 56286 -16326
rect 56341 -16360 56382 -16326
rect 56437 -16360 56478 -16326
rect 56533 -16360 56574 -16326
rect 56629 -16360 56670 -16326
rect 56725 -16360 56766 -16326
rect 55070 -16410 55111 -16376
rect 55703 -16379 55710 -16371
rect 54720 -16451 54761 -16417
rect 54709 -16500 54716 -16489
rect 54720 -16500 54725 -16451
rect 54914 -16494 54955 -16460
rect 54959 -16494 54966 -16449
rect 55059 -16460 55066 -16449
rect 55268 -16453 55309 -16419
rect 55313 -16453 55320 -16408
rect 55413 -16419 55420 -16408
rect 55594 -16413 55635 -16379
rect 55658 -16413 55710 -16379
rect 55738 -16413 55779 -16379
rect 55424 -16453 55465 -16419
rect 55070 -16494 55111 -16460
rect 54720 -16534 54761 -16500
rect 54720 -16568 54725 -16534
rect 53369 -16740 53375 -16706
rect 53666 -16723 53707 -16689
rect 53711 -16723 53718 -16681
rect 51116 -16906 51158 -16872
rect 51188 -16906 51230 -16872
rect 51260 -16906 51302 -16872
rect 51573 -16913 51615 -16879
rect 51618 -16913 51626 -16868
rect 51718 -16879 51726 -16868
rect 51729 -16913 51771 -16879
rect 52313 -16895 52355 -16861
rect 52358 -16895 52366 -16853
rect 50207 -16959 50690 -16925
rect 51541 -16949 51583 -16915
rect 51613 -16949 51655 -16915
rect 51927 -16956 51969 -16922
rect 51972 -16956 51980 -16911
rect 52072 -16922 52080 -16911
rect 52500 -16913 52513 -16845
rect 52541 -16879 52547 -16811
rect 52586 -16843 52592 -16775
rect 52620 -16809 52626 -16743
rect 52630 -16793 52672 -16759
rect 52833 -16838 52875 -16804
rect 52600 -16861 52608 -16853
rect 52611 -16895 52653 -16861
rect 52833 -16906 52875 -16872
rect 52083 -16956 52125 -16922
rect 50207 -16985 50677 -16959
rect 50211 -16993 50419 -16985
rect 50227 -17003 50403 -16993
rect 49953 -17140 50135 -17114
rect 49460 -17174 49502 -17140
rect 49556 -17174 49598 -17140
rect 49652 -17174 49694 -17140
rect 49748 -17174 49790 -17140
rect 49844 -17174 49886 -17140
rect 49940 -17174 50135 -17140
rect 49953 -17200 50135 -17174
rect 50153 -17174 50261 -17050
rect 50412 -17062 50419 -17051
rect 50031 -17870 50073 -17200
rect 50153 -17228 50163 -17174
rect 49838 -17936 49990 -17924
rect 49506 -17970 49990 -17936
rect 49838 -17971 49990 -17970
rect 50019 -17971 50073 -17870
rect 50165 -17971 50207 -17174
rect 50211 -17971 50218 -17174
rect 50423 -17971 50465 -17062
rect 50557 -17971 50599 -16985
rect 50810 -17002 50852 -16968
rect 50906 -17002 50948 -16968
rect 51002 -17002 51044 -16968
rect 51098 -17002 51140 -16968
rect 51194 -17002 51236 -16968
rect 51290 -17002 51332 -16968
rect 51386 -17002 51428 -16968
rect 51895 -16992 51937 -16958
rect 51967 -16992 52009 -16958
rect 52313 -16995 52355 -16961
rect 52358 -16995 52366 -16950
rect 52500 -17001 52508 -16913
rect 52882 -16922 52888 -16788
rect 52600 -16961 52608 -16950
rect 52916 -16956 52922 -16762
rect 52956 -16778 52964 -16767
rect 52952 -16809 52964 -16778
rect 53278 -16796 53320 -16762
rect 52611 -16995 52653 -16961
rect 51548 -17045 51590 -17011
rect 51644 -17045 51686 -17011
rect 51740 -17045 51782 -17011
rect 52249 -17035 52291 -17001
rect 52321 -17035 52363 -17001
rect 52393 -17035 52435 -17001
rect 52465 -17029 52508 -17001
rect 52811 -17025 52853 -16991
rect 52856 -17025 52864 -16980
rect 52952 -16992 52958 -16809
rect 52986 -16995 52992 -16812
rect 52465 -17035 52507 -17029
rect 51902 -17088 51944 -17054
rect 51998 -17088 52040 -17054
rect 52094 -17088 52136 -17054
rect 52998 -17076 53006 -16809
rect 53335 -16812 53336 -16742
rect 53369 -16819 53370 -16740
rect 53853 -16741 53865 -16673
rect 53894 -16707 53899 -16639
rect 53939 -16671 53944 -16603
rect 53973 -16637 53978 -16571
rect 54914 -16577 54955 -16543
rect 54959 -16577 54966 -16532
rect 55059 -16543 55066 -16532
rect 55268 -16537 55309 -16503
rect 55313 -16537 55320 -16492
rect 55413 -16503 55420 -16492
rect 55658 -16496 55699 -16462
rect 55703 -16496 55710 -16451
rect 55424 -16537 55465 -16503
rect 55070 -16577 55111 -16543
rect 53983 -16621 54024 -16587
rect 54184 -16666 54225 -16632
rect 53953 -16689 53960 -16681
rect 53964 -16723 54005 -16689
rect 54184 -16734 54225 -16700
rect 53853 -16753 53860 -16741
rect 54233 -16750 54238 -16616
rect 53628 -16819 54021 -16753
rect 54267 -16784 54272 -16590
rect 54307 -16606 54314 -16595
rect 54303 -16637 54314 -16606
rect 54629 -16624 54670 -16590
rect 53014 -16860 53056 -16826
rect 53363 -16830 53381 -16819
rect 53363 -16832 53370 -16830
rect 53014 -16928 53056 -16894
rect 53066 -16995 53072 -16860
rect 53297 -16874 53370 -16832
rect 53426 -16874 54021 -16819
rect 54162 -16853 54203 -16819
rect 54207 -16853 54214 -16808
rect 54303 -16820 54308 -16637
rect 54337 -16823 54342 -16640
rect 53297 -16877 54021 -16874
rect 53100 -16980 53106 -16892
rect 53217 -16942 53259 -16908
rect 53262 -16942 53270 -16900
rect 53098 -16991 53106 -16980
rect 53100 -17025 53106 -16991
rect 53109 -17025 53151 -16991
rect 53217 -17042 53259 -17008
rect 53262 -17042 53270 -16997
rect 53110 -17078 53152 -17044
rect 53182 -17078 53224 -17044
rect 53254 -17078 53296 -17044
rect 52256 -17131 52298 -17097
rect 52352 -17131 52394 -17097
rect 52448 -17131 52490 -17097
rect 52544 -17131 52586 -17097
rect 52640 -17131 52682 -17097
rect 53297 -17114 53449 -16877
rect 53628 -16899 54021 -16877
rect 53552 -16925 54021 -16899
rect 54349 -16904 54356 -16637
rect 54365 -16688 54406 -16654
rect 54365 -16756 54406 -16722
rect 54417 -16823 54422 -16688
rect 54979 -16691 55020 -16657
rect 55031 -16718 55036 -16641
rect 54451 -16808 54456 -16720
rect 54568 -16770 54609 -16736
rect 54613 -16770 54620 -16728
rect 54713 -16740 54720 -16729
rect 54724 -16774 54765 -16740
rect 55065 -16752 55070 -16607
rect 55268 -16620 55309 -16586
rect 55313 -16620 55320 -16575
rect 55413 -16586 55420 -16575
rect 55658 -16580 55699 -16546
rect 55703 -16580 55710 -16535
rect 55424 -16620 55465 -16586
rect 55333 -16734 55374 -16700
rect 55385 -16761 55390 -16684
rect 54449 -16819 54456 -16808
rect 54918 -16813 54959 -16779
rect 54963 -16813 54970 -16771
rect 55063 -16779 55070 -16771
rect 55074 -16813 55115 -16779
rect 55419 -16795 55424 -16650
rect 55658 -16663 55699 -16629
rect 55703 -16663 55710 -16618
rect 55780 -16679 55785 -16363
rect 55803 -16379 55810 -16371
rect 55814 -16379 55819 -16363
rect 55814 -16413 55855 -16379
rect 55859 -16413 55866 -16371
rect 55803 -16462 55810 -16451
rect 55814 -16462 55819 -16413
rect 55814 -16496 55855 -16462
rect 55859 -16496 55866 -16451
rect 55803 -16546 55810 -16535
rect 55814 -16546 55819 -16496
rect 55814 -16580 55855 -16546
rect 55859 -16580 55866 -16535
rect 55803 -16629 55810 -16618
rect 55814 -16629 55819 -16580
rect 55814 -16663 55855 -16629
rect 55859 -16663 55866 -16618
rect 55803 -16697 55810 -16671
rect 55814 -16713 55819 -16663
rect 55723 -16777 55764 -16743
rect 54451 -16853 54456 -16819
rect 54460 -16853 54501 -16819
rect 54568 -16870 54609 -16836
rect 54613 -16870 54620 -16825
rect 54713 -16832 54720 -16821
rect 54724 -16866 54765 -16832
rect 55272 -16856 55313 -16822
rect 55317 -16856 55324 -16814
rect 55417 -16822 55424 -16814
rect 55428 -16856 55469 -16822
rect 55845 -16845 55852 -16697
rect 55868 -16713 55871 -16363
rect 55902 -16679 55905 -16363
rect 55959 -16379 55966 -16371
rect 55908 -16413 55949 -16379
rect 55970 -16413 56021 -16379
rect 56680 -16422 56685 -16406
rect 56703 -16422 56710 -16414
rect 56714 -16422 56719 -16406
rect 57010 -16408 57051 -16374
rect 57055 -16408 57062 -16363
rect 55959 -16462 55966 -16451
rect 56140 -16456 56181 -16422
rect 56212 -16456 56253 -16422
rect 56284 -16456 56325 -16422
rect 56428 -16456 56469 -16422
rect 56500 -16456 56613 -16422
rect 56644 -16456 56685 -16422
rect 55970 -16496 56011 -16462
rect 55959 -16546 55966 -16535
rect 56537 -16539 56578 -16505
rect 55970 -16580 56011 -16546
rect 55959 -16629 55966 -16618
rect 55970 -16663 56011 -16629
rect 56202 -16689 56243 -16655
rect 56247 -16689 56254 -16644
rect 56324 -16706 56329 -16588
rect 56347 -16655 56354 -16644
rect 56358 -16655 56363 -16622
rect 56394 -16655 56399 -16622
rect 56358 -16689 56399 -16655
rect 56403 -16689 56410 -16644
rect 56358 -16740 56363 -16689
rect 56394 -16740 56399 -16689
rect 56428 -16706 56433 -16589
rect 56537 -16623 56578 -16589
rect 56537 -16706 56578 -16672
rect 56680 -16706 56685 -16456
rect 56714 -16456 56755 -16422
rect 56703 -16505 56710 -16494
rect 56714 -16505 56719 -16456
rect 57010 -16491 57051 -16457
rect 57055 -16491 57062 -16446
rect 56714 -16539 56755 -16505
rect 56703 -16589 56710 -16578
rect 56714 -16589 56719 -16539
rect 56863 -16565 56972 -16499
rect 57132 -16507 57137 -16191
rect 57155 -16207 57162 -16199
rect 57166 -16207 57171 -16191
rect 57166 -16241 57207 -16207
rect 57211 -16241 57218 -16199
rect 57155 -16290 57162 -16279
rect 57166 -16290 57171 -16241
rect 57166 -16324 57207 -16290
rect 57211 -16324 57218 -16279
rect 57155 -16374 57162 -16363
rect 57166 -16374 57171 -16324
rect 57166 -16408 57207 -16374
rect 57211 -16408 57218 -16363
rect 57155 -16457 57162 -16446
rect 57166 -16457 57171 -16408
rect 57166 -16491 57207 -16457
rect 57211 -16491 57218 -16446
rect 57155 -16525 57162 -16499
rect 57166 -16541 57171 -16491
rect 56714 -16623 56755 -16589
rect 57075 -16605 57116 -16571
rect 56703 -16672 56710 -16661
rect 56714 -16672 56719 -16623
rect 56714 -16706 56755 -16672
rect 57197 -16673 57204 -16525
rect 57220 -16541 57223 -16191
rect 57254 -16507 57257 -16191
rect 57311 -16207 57318 -16199
rect 57260 -16241 57301 -16207
rect 57322 -16241 57373 -16207
rect 58237 -16231 58278 -16197
rect 58333 -16231 58374 -16197
rect 58429 -16231 58470 -16197
rect 60399 -16207 60406 -16199
rect 58030 -16250 58035 -16234
rect 58053 -16250 58060 -16242
rect 58064 -16250 58069 -16234
rect 57311 -16290 57318 -16279
rect 57490 -16284 57531 -16250
rect 57562 -16284 57603 -16250
rect 57634 -16284 57675 -16250
rect 57778 -16284 57819 -16250
rect 57850 -16284 57963 -16250
rect 57994 -16284 58035 -16250
rect 57322 -16324 57363 -16290
rect 57311 -16374 57318 -16363
rect 57887 -16367 57928 -16333
rect 57322 -16408 57363 -16374
rect 57311 -16457 57318 -16446
rect 57322 -16491 57363 -16457
rect 57552 -16517 57593 -16483
rect 57597 -16517 57604 -16472
rect 57674 -16534 57679 -16416
rect 57697 -16483 57704 -16472
rect 57708 -16483 57713 -16450
rect 57744 -16483 57749 -16450
rect 57708 -16517 57749 -16483
rect 57753 -16517 57760 -16472
rect 57708 -16568 57713 -16517
rect 57744 -16568 57749 -16517
rect 57778 -16534 57783 -16417
rect 57887 -16451 57928 -16417
rect 57887 -16534 57928 -16500
rect 58030 -16534 58035 -16284
rect 58064 -16284 58105 -16250
rect 58591 -16274 58632 -16240
rect 58687 -16274 58728 -16240
rect 58783 -16274 58824 -16240
rect 60290 -16241 60331 -16207
rect 60354 -16241 60406 -16207
rect 60434 -16241 60475 -16207
rect 58053 -16333 58060 -16322
rect 58064 -16333 58069 -16284
rect 58303 -16293 58310 -16285
rect 58403 -16293 58410 -16285
rect 58230 -16327 58299 -16293
rect 58302 -16327 58343 -16293
rect 58414 -16327 58455 -16293
rect 58945 -16317 58986 -16283
rect 59041 -16317 59082 -16283
rect 59137 -16317 59178 -16283
rect 59233 -16317 59274 -16283
rect 59329 -16317 59370 -16283
rect 60354 -16324 60395 -16290
rect 60399 -16324 60406 -16279
rect 58064 -16367 58105 -16333
rect 58657 -16336 58664 -16328
rect 58757 -16336 58764 -16328
rect 58053 -16417 58060 -16406
rect 58064 -16417 58069 -16367
rect 58258 -16410 58299 -16376
rect 58303 -16410 58310 -16365
rect 58403 -16376 58410 -16365
rect 58584 -16370 58653 -16336
rect 58656 -16370 58697 -16336
rect 58768 -16370 58809 -16336
rect 59493 -16360 59534 -16326
rect 59589 -16360 59630 -16326
rect 59685 -16360 59726 -16326
rect 59781 -16360 59822 -16326
rect 59877 -16360 59918 -16326
rect 59973 -16360 60014 -16326
rect 60069 -16360 60110 -16326
rect 58414 -16410 58455 -16376
rect 59047 -16379 59054 -16371
rect 58064 -16451 58105 -16417
rect 58053 -16500 58060 -16489
rect 58064 -16500 58069 -16451
rect 58258 -16494 58299 -16460
rect 58303 -16494 58310 -16449
rect 58403 -16460 58410 -16449
rect 58612 -16453 58653 -16419
rect 58657 -16453 58664 -16408
rect 58757 -16419 58764 -16408
rect 58938 -16413 58979 -16379
rect 59002 -16413 59054 -16379
rect 59082 -16413 59123 -16379
rect 58768 -16453 58809 -16419
rect 58414 -16494 58455 -16460
rect 58064 -16534 58105 -16500
rect 58064 -16568 58069 -16534
rect 56714 -16740 56719 -16706
rect 57010 -16723 57051 -16689
rect 57055 -16723 57062 -16681
rect 57197 -16741 57209 -16673
rect 57238 -16707 57243 -16639
rect 57283 -16671 57288 -16603
rect 57317 -16637 57322 -16571
rect 58258 -16577 58299 -16543
rect 58303 -16577 58310 -16532
rect 58403 -16543 58410 -16532
rect 58612 -16537 58653 -16503
rect 58657 -16537 58664 -16492
rect 58757 -16503 58764 -16492
rect 59002 -16496 59043 -16462
rect 59047 -16496 59054 -16451
rect 58768 -16537 58809 -16503
rect 58414 -16577 58455 -16543
rect 57327 -16621 57368 -16587
rect 57528 -16666 57569 -16632
rect 57297 -16689 57304 -16681
rect 57308 -16723 57349 -16689
rect 57528 -16734 57569 -16700
rect 54461 -16906 54502 -16872
rect 54533 -16906 54574 -16872
rect 54605 -16906 54646 -16872
rect 54918 -16913 54959 -16879
rect 54963 -16913 54970 -16868
rect 55063 -16879 55070 -16868
rect 55074 -16913 55115 -16879
rect 55658 -16895 55699 -16861
rect 55703 -16895 55710 -16853
rect 53552 -16959 54034 -16925
rect 54886 -16949 54927 -16915
rect 54958 -16949 54999 -16915
rect 55272 -16956 55313 -16922
rect 55317 -16956 55324 -16911
rect 55417 -16922 55424 -16911
rect 55845 -16913 55857 -16845
rect 55886 -16879 55891 -16811
rect 55931 -16843 55936 -16775
rect 55965 -16809 55970 -16743
rect 57197 -16753 57204 -16741
rect 57577 -16750 57582 -16616
rect 55975 -16793 56016 -16759
rect 56178 -16838 56219 -16804
rect 55945 -16861 55952 -16853
rect 55956 -16895 55997 -16861
rect 56178 -16906 56219 -16872
rect 55428 -16956 55469 -16922
rect 53552 -16985 54021 -16959
rect 53555 -16993 53763 -16985
rect 53571 -17003 53747 -16993
rect 53297 -17140 53479 -17114
rect 52804 -17174 52846 -17140
rect 52900 -17174 52942 -17140
rect 52996 -17174 53038 -17140
rect 53092 -17174 53134 -17140
rect 53188 -17174 53230 -17140
rect 53284 -17174 53479 -17140
rect 53297 -17200 53479 -17174
rect 53497 -17174 53605 -17050
rect 53756 -17062 53763 -17051
rect 53375 -17870 53417 -17200
rect 53497 -17228 53507 -17174
rect 53182 -17936 53334 -17924
rect 52850 -17970 53334 -17936
rect 53182 -17971 53334 -17970
rect 53363 -17971 53417 -17870
rect 53509 -17971 53551 -17174
rect 53555 -17971 53562 -17174
rect 53767 -17971 53809 -17062
rect 53901 -17971 53943 -16985
rect 54155 -17002 54196 -16968
rect 54251 -17002 54292 -16968
rect 54347 -17002 54388 -16968
rect 54443 -17002 54484 -16968
rect 54539 -17002 54580 -16968
rect 54635 -17002 54676 -16968
rect 54731 -17002 54772 -16968
rect 55240 -16992 55281 -16958
rect 55312 -16992 55353 -16958
rect 55658 -16995 55699 -16961
rect 55703 -16995 55710 -16950
rect 55845 -17001 55852 -16913
rect 56227 -16922 56232 -16788
rect 55945 -16961 55952 -16950
rect 56261 -16956 56266 -16762
rect 56301 -16778 56308 -16767
rect 56297 -16809 56308 -16778
rect 56623 -16796 56664 -16762
rect 55956 -16995 55997 -16961
rect 54893 -17045 54934 -17011
rect 54989 -17045 55030 -17011
rect 55085 -17045 55126 -17011
rect 55594 -17035 55635 -17001
rect 55666 -17035 55707 -17001
rect 55738 -17035 55779 -17001
rect 55810 -17029 55852 -17001
rect 56156 -17025 56197 -16991
rect 56201 -17025 56208 -16980
rect 56297 -16992 56302 -16809
rect 56331 -16995 56336 -16812
rect 55810 -17035 55851 -17029
rect 55247 -17088 55288 -17054
rect 55343 -17088 55384 -17054
rect 55439 -17088 55480 -17054
rect 56343 -17076 56350 -16809
rect 56972 -16819 57365 -16753
rect 57611 -16784 57616 -16590
rect 57651 -16606 57658 -16595
rect 57647 -16637 57658 -16606
rect 57973 -16624 58014 -16590
rect 56359 -16860 56400 -16826
rect 56708 -16830 56725 -16819
rect 56708 -16832 56714 -16830
rect 56359 -16928 56400 -16894
rect 56411 -16995 56416 -16860
rect 56642 -16874 56714 -16832
rect 56770 -16874 57365 -16819
rect 57506 -16853 57547 -16819
rect 57551 -16853 57558 -16808
rect 57647 -16820 57652 -16637
rect 57681 -16823 57686 -16640
rect 56642 -16877 57365 -16874
rect 56445 -16980 56450 -16892
rect 56562 -16942 56603 -16908
rect 56607 -16942 56614 -16900
rect 56443 -16991 56450 -16980
rect 56445 -17025 56450 -16991
rect 56454 -17025 56495 -16991
rect 56562 -17042 56603 -17008
rect 56607 -17042 56614 -16997
rect 56455 -17078 56496 -17044
rect 56527 -17078 56568 -17044
rect 56599 -17078 56640 -17044
rect 55601 -17131 55642 -17097
rect 55697 -17131 55738 -17097
rect 55793 -17131 55834 -17097
rect 55889 -17131 55930 -17097
rect 55985 -17131 56026 -17097
rect 56642 -17114 56793 -16877
rect 56972 -16899 57365 -16877
rect 56896 -16925 57365 -16899
rect 57693 -16904 57700 -16637
rect 57709 -16688 57750 -16654
rect 57709 -16756 57750 -16722
rect 57761 -16823 57766 -16688
rect 58323 -16691 58364 -16657
rect 58375 -16718 58380 -16641
rect 57795 -16808 57800 -16720
rect 57912 -16770 57953 -16736
rect 57957 -16770 57964 -16728
rect 58057 -16740 58064 -16729
rect 58068 -16774 58109 -16740
rect 58409 -16752 58414 -16607
rect 58612 -16620 58653 -16586
rect 58657 -16620 58664 -16575
rect 58757 -16586 58764 -16575
rect 59002 -16580 59043 -16546
rect 59047 -16580 59054 -16535
rect 58768 -16620 58809 -16586
rect 58677 -16734 58718 -16700
rect 58729 -16761 58734 -16684
rect 57793 -16819 57800 -16808
rect 58262 -16813 58303 -16779
rect 58307 -16813 58314 -16771
rect 58407 -16779 58414 -16771
rect 58418 -16813 58459 -16779
rect 58763 -16795 58768 -16650
rect 59002 -16663 59043 -16629
rect 59047 -16663 59054 -16618
rect 59124 -16679 59129 -16363
rect 59147 -16379 59154 -16371
rect 59158 -16379 59163 -16363
rect 59158 -16413 59199 -16379
rect 59203 -16413 59210 -16371
rect 59147 -16462 59154 -16451
rect 59158 -16462 59163 -16413
rect 59158 -16496 59199 -16462
rect 59203 -16496 59210 -16451
rect 59147 -16546 59154 -16535
rect 59158 -16546 59163 -16496
rect 59158 -16580 59199 -16546
rect 59203 -16580 59210 -16535
rect 59147 -16629 59154 -16618
rect 59158 -16629 59163 -16580
rect 59158 -16663 59199 -16629
rect 59203 -16663 59210 -16618
rect 59147 -16697 59154 -16671
rect 59158 -16713 59163 -16663
rect 59067 -16777 59108 -16743
rect 57795 -16853 57800 -16819
rect 57804 -16853 57845 -16819
rect 57912 -16870 57953 -16836
rect 57957 -16870 57964 -16825
rect 58057 -16832 58064 -16821
rect 58068 -16866 58109 -16832
rect 58616 -16856 58657 -16822
rect 58661 -16856 58668 -16814
rect 58761 -16822 58768 -16814
rect 58772 -16856 58813 -16822
rect 59189 -16845 59196 -16697
rect 59212 -16713 59215 -16363
rect 59246 -16679 59249 -16363
rect 59303 -16379 59310 -16371
rect 59252 -16413 59293 -16379
rect 59314 -16413 59365 -16379
rect 60024 -16422 60029 -16406
rect 60047 -16422 60054 -16414
rect 60058 -16422 60063 -16406
rect 60354 -16408 60395 -16374
rect 60399 -16408 60406 -16363
rect 59303 -16462 59310 -16451
rect 59484 -16456 59525 -16422
rect 59556 -16456 59597 -16422
rect 59628 -16456 59669 -16422
rect 59772 -16456 59813 -16422
rect 59844 -16456 59957 -16422
rect 59988 -16456 60029 -16422
rect 59314 -16496 59355 -16462
rect 59303 -16546 59310 -16535
rect 59881 -16539 59922 -16505
rect 59314 -16580 59355 -16546
rect 59303 -16629 59310 -16618
rect 59314 -16663 59355 -16629
rect 59546 -16689 59587 -16655
rect 59591 -16689 59598 -16644
rect 59668 -16706 59673 -16588
rect 59691 -16655 59698 -16644
rect 59702 -16655 59707 -16622
rect 59738 -16655 59743 -16622
rect 59702 -16689 59743 -16655
rect 59747 -16689 59754 -16644
rect 59702 -16740 59707 -16689
rect 59738 -16740 59743 -16689
rect 59772 -16706 59777 -16589
rect 59881 -16623 59922 -16589
rect 59881 -16706 59922 -16672
rect 60024 -16706 60029 -16456
rect 60058 -16456 60099 -16422
rect 60047 -16505 60054 -16494
rect 60058 -16505 60063 -16456
rect 60354 -16491 60395 -16457
rect 60399 -16491 60406 -16446
rect 60058 -16539 60099 -16505
rect 60047 -16589 60054 -16578
rect 60058 -16589 60063 -16539
rect 60207 -16565 60316 -16499
rect 60476 -16507 60481 -16191
rect 60499 -16207 60506 -16199
rect 60510 -16207 60515 -16191
rect 60510 -16241 60551 -16207
rect 60555 -16241 60562 -16199
rect 60499 -16290 60506 -16279
rect 60510 -16290 60515 -16241
rect 60510 -16324 60551 -16290
rect 60555 -16324 60562 -16279
rect 60499 -16374 60506 -16363
rect 60510 -16374 60515 -16324
rect 60510 -16408 60551 -16374
rect 60555 -16408 60562 -16363
rect 60499 -16457 60506 -16446
rect 60510 -16457 60515 -16408
rect 60510 -16491 60551 -16457
rect 60555 -16491 60562 -16446
rect 60499 -16525 60506 -16499
rect 60510 -16541 60515 -16491
rect 60058 -16623 60099 -16589
rect 60419 -16605 60460 -16571
rect 60047 -16672 60054 -16661
rect 60058 -16672 60063 -16623
rect 60058 -16706 60099 -16672
rect 60541 -16673 60548 -16525
rect 60564 -16541 60567 -16191
rect 60598 -16507 60601 -16191
rect 60655 -16207 60662 -16199
rect 60604 -16241 60645 -16207
rect 60666 -16241 60717 -16207
rect 61581 -16231 61622 -16197
rect 61677 -16231 61718 -16197
rect 61773 -16231 61814 -16197
rect 63743 -16207 63750 -16199
rect 61374 -16250 61379 -16234
rect 61397 -16250 61404 -16242
rect 61408 -16250 61413 -16234
rect 60655 -16290 60662 -16279
rect 60834 -16284 60875 -16250
rect 60906 -16284 60947 -16250
rect 60978 -16284 61019 -16250
rect 61122 -16284 61163 -16250
rect 61194 -16284 61307 -16250
rect 61338 -16284 61379 -16250
rect 60666 -16324 60707 -16290
rect 60655 -16374 60662 -16363
rect 61231 -16367 61272 -16333
rect 60666 -16408 60707 -16374
rect 60655 -16457 60662 -16446
rect 60666 -16491 60707 -16457
rect 60896 -16517 60937 -16483
rect 60941 -16517 60948 -16472
rect 61018 -16534 61023 -16416
rect 61041 -16483 61048 -16472
rect 61052 -16483 61057 -16450
rect 61088 -16483 61093 -16450
rect 61052 -16517 61093 -16483
rect 61097 -16517 61104 -16472
rect 61052 -16568 61057 -16517
rect 61088 -16568 61093 -16517
rect 61122 -16534 61127 -16417
rect 61231 -16451 61272 -16417
rect 61231 -16534 61272 -16500
rect 61374 -16534 61379 -16284
rect 61408 -16284 61449 -16250
rect 61935 -16274 61976 -16240
rect 62031 -16274 62072 -16240
rect 62127 -16274 62168 -16240
rect 63634 -16241 63675 -16207
rect 63698 -16241 63750 -16207
rect 63778 -16241 63819 -16207
rect 61397 -16333 61404 -16322
rect 61408 -16333 61413 -16284
rect 61647 -16293 61654 -16285
rect 61747 -16293 61754 -16285
rect 61574 -16327 61643 -16293
rect 61646 -16327 61687 -16293
rect 61758 -16327 61799 -16293
rect 62289 -16317 62330 -16283
rect 62385 -16317 62426 -16283
rect 62481 -16317 62522 -16283
rect 62577 -16317 62618 -16283
rect 62673 -16317 62714 -16283
rect 63698 -16324 63739 -16290
rect 63743 -16324 63750 -16279
rect 61408 -16367 61449 -16333
rect 62001 -16336 62008 -16328
rect 62101 -16336 62108 -16328
rect 61397 -16417 61404 -16406
rect 61408 -16417 61413 -16367
rect 61602 -16410 61643 -16376
rect 61647 -16410 61654 -16365
rect 61747 -16376 61754 -16365
rect 61928 -16370 61997 -16336
rect 62000 -16370 62041 -16336
rect 62112 -16370 62153 -16336
rect 62837 -16360 62878 -16326
rect 62933 -16360 62974 -16326
rect 63029 -16360 63070 -16326
rect 63125 -16360 63166 -16326
rect 63221 -16360 63262 -16326
rect 63317 -16360 63358 -16326
rect 63413 -16360 63454 -16326
rect 61758 -16410 61799 -16376
rect 62391 -16379 62398 -16371
rect 61408 -16451 61449 -16417
rect 61397 -16500 61404 -16489
rect 61408 -16500 61413 -16451
rect 61602 -16494 61643 -16460
rect 61647 -16494 61654 -16449
rect 61747 -16460 61754 -16449
rect 61956 -16453 61997 -16419
rect 62001 -16453 62008 -16408
rect 62101 -16419 62108 -16408
rect 62282 -16413 62323 -16379
rect 62346 -16413 62398 -16379
rect 62426 -16413 62467 -16379
rect 62112 -16453 62153 -16419
rect 61758 -16494 61799 -16460
rect 61408 -16534 61449 -16500
rect 61408 -16568 61413 -16534
rect 60058 -16740 60063 -16706
rect 60354 -16723 60395 -16689
rect 60399 -16723 60406 -16681
rect 60541 -16741 60553 -16673
rect 60582 -16707 60587 -16639
rect 60627 -16671 60632 -16603
rect 60661 -16637 60666 -16571
rect 61602 -16577 61643 -16543
rect 61647 -16577 61654 -16532
rect 61747 -16543 61754 -16532
rect 61956 -16537 61997 -16503
rect 62001 -16537 62008 -16492
rect 62101 -16503 62108 -16492
rect 62346 -16496 62387 -16462
rect 62391 -16496 62398 -16451
rect 62112 -16537 62153 -16503
rect 61758 -16577 61799 -16543
rect 60671 -16621 60712 -16587
rect 60872 -16666 60913 -16632
rect 60641 -16689 60648 -16681
rect 60652 -16723 60693 -16689
rect 60872 -16734 60913 -16700
rect 57805 -16906 57846 -16872
rect 57877 -16906 57918 -16872
rect 57949 -16906 57990 -16872
rect 58262 -16913 58303 -16879
rect 58307 -16913 58314 -16868
rect 58407 -16879 58414 -16868
rect 58418 -16913 58459 -16879
rect 59002 -16895 59043 -16861
rect 59047 -16895 59054 -16853
rect 56896 -16959 57378 -16925
rect 58230 -16949 58271 -16915
rect 58302 -16949 58343 -16915
rect 58616 -16956 58657 -16922
rect 58661 -16956 58668 -16911
rect 58761 -16922 58768 -16911
rect 59189 -16913 59201 -16845
rect 59230 -16879 59235 -16811
rect 59275 -16843 59280 -16775
rect 59309 -16809 59314 -16743
rect 60541 -16753 60548 -16741
rect 60921 -16750 60926 -16616
rect 59319 -16793 59360 -16759
rect 59522 -16838 59563 -16804
rect 59289 -16861 59296 -16853
rect 59300 -16895 59341 -16861
rect 59522 -16906 59563 -16872
rect 58772 -16956 58813 -16922
rect 56896 -16985 57365 -16959
rect 56900 -16993 57107 -16985
rect 56916 -17003 57091 -16993
rect 56642 -17140 56823 -17114
rect 56149 -17174 56190 -17140
rect 56245 -17174 56286 -17140
rect 56341 -17174 56382 -17140
rect 56437 -17174 56478 -17140
rect 56533 -17174 56574 -17140
rect 56629 -17174 56823 -17140
rect 56642 -17200 56823 -17174
rect 56842 -17174 56949 -17050
rect 57101 -17062 57107 -17051
rect 56720 -17870 56761 -17200
rect 56842 -17228 56851 -17174
rect 56527 -17936 56678 -17924
rect 56195 -17970 56678 -17936
rect 56527 -17971 56678 -17970
rect 56708 -17971 56761 -17870
rect 56854 -17971 56895 -17174
rect 56900 -17971 56906 -17174
rect 57112 -17971 57153 -17062
rect 57246 -17971 57287 -16985
rect 57499 -17002 57540 -16968
rect 57595 -17002 57636 -16968
rect 57691 -17002 57732 -16968
rect 57787 -17002 57828 -16968
rect 57883 -17002 57924 -16968
rect 57979 -17002 58020 -16968
rect 58075 -17002 58116 -16968
rect 58584 -16992 58625 -16958
rect 58656 -16992 58697 -16958
rect 59002 -16995 59043 -16961
rect 59047 -16995 59054 -16950
rect 59189 -17001 59196 -16913
rect 59571 -16922 59576 -16788
rect 59289 -16961 59296 -16950
rect 59605 -16956 59610 -16762
rect 59645 -16778 59652 -16767
rect 59641 -16809 59652 -16778
rect 59967 -16796 60008 -16762
rect 59300 -16995 59341 -16961
rect 58237 -17045 58278 -17011
rect 58333 -17045 58374 -17011
rect 58429 -17045 58470 -17011
rect 58938 -17035 58979 -17001
rect 59010 -17035 59051 -17001
rect 59082 -17035 59123 -17001
rect 59154 -17029 59196 -17001
rect 59500 -17025 59541 -16991
rect 59545 -17025 59552 -16980
rect 59641 -16992 59646 -16809
rect 59675 -16995 59680 -16812
rect 59154 -17035 59195 -17029
rect 58591 -17088 58632 -17054
rect 58687 -17088 58728 -17054
rect 58783 -17088 58824 -17054
rect 59687 -17076 59694 -16809
rect 60316 -16819 60709 -16753
rect 60955 -16784 60960 -16590
rect 60995 -16606 61002 -16595
rect 60991 -16637 61002 -16606
rect 61317 -16624 61358 -16590
rect 59703 -16860 59744 -16826
rect 60052 -16830 60069 -16819
rect 60052 -16832 60058 -16830
rect 59703 -16928 59744 -16894
rect 59755 -16995 59760 -16860
rect 59986 -16874 60058 -16832
rect 60114 -16874 60709 -16819
rect 60850 -16853 60891 -16819
rect 60895 -16853 60902 -16808
rect 60991 -16820 60996 -16637
rect 61025 -16823 61030 -16640
rect 59986 -16877 60709 -16874
rect 59789 -16980 59794 -16892
rect 59906 -16942 59947 -16908
rect 59951 -16942 59958 -16900
rect 59787 -16991 59794 -16980
rect 59789 -17025 59794 -16991
rect 59798 -17025 59839 -16991
rect 59906 -17042 59947 -17008
rect 59951 -17042 59958 -16997
rect 59799 -17078 59840 -17044
rect 59871 -17078 59912 -17044
rect 59943 -17078 59984 -17044
rect 58945 -17131 58986 -17097
rect 59041 -17131 59082 -17097
rect 59137 -17131 59178 -17097
rect 59233 -17131 59274 -17097
rect 59329 -17131 59370 -17097
rect 59986 -17114 60137 -16877
rect 60316 -16899 60709 -16877
rect 60240 -16925 60709 -16899
rect 61037 -16904 61044 -16637
rect 61053 -16688 61094 -16654
rect 61053 -16756 61094 -16722
rect 61105 -16823 61110 -16688
rect 61667 -16691 61708 -16657
rect 61719 -16718 61724 -16641
rect 61139 -16808 61144 -16720
rect 61256 -16770 61297 -16736
rect 61301 -16770 61308 -16728
rect 61401 -16740 61408 -16729
rect 61412 -16774 61453 -16740
rect 61753 -16752 61758 -16607
rect 61956 -16620 61997 -16586
rect 62001 -16620 62008 -16575
rect 62101 -16586 62108 -16575
rect 62346 -16580 62387 -16546
rect 62391 -16580 62398 -16535
rect 62112 -16620 62153 -16586
rect 62021 -16734 62062 -16700
rect 62073 -16761 62078 -16684
rect 61137 -16819 61144 -16808
rect 61606 -16813 61647 -16779
rect 61651 -16813 61658 -16771
rect 61751 -16779 61758 -16771
rect 61762 -16813 61803 -16779
rect 62107 -16795 62112 -16650
rect 62346 -16663 62387 -16629
rect 62391 -16663 62398 -16618
rect 62468 -16679 62473 -16363
rect 62491 -16379 62498 -16371
rect 62502 -16379 62507 -16363
rect 62502 -16413 62543 -16379
rect 62547 -16413 62554 -16371
rect 62491 -16462 62498 -16451
rect 62502 -16462 62507 -16413
rect 62502 -16496 62543 -16462
rect 62547 -16496 62554 -16451
rect 62491 -16546 62498 -16535
rect 62502 -16546 62507 -16496
rect 62502 -16580 62543 -16546
rect 62547 -16580 62554 -16535
rect 62491 -16629 62498 -16618
rect 62502 -16629 62507 -16580
rect 62502 -16663 62543 -16629
rect 62547 -16663 62554 -16618
rect 62491 -16697 62498 -16671
rect 62502 -16713 62507 -16663
rect 62411 -16777 62452 -16743
rect 61139 -16853 61144 -16819
rect 61148 -16853 61189 -16819
rect 61256 -16870 61297 -16836
rect 61301 -16870 61308 -16825
rect 61401 -16832 61408 -16821
rect 61412 -16866 61453 -16832
rect 61960 -16856 62001 -16822
rect 62005 -16856 62012 -16814
rect 62105 -16822 62112 -16814
rect 62116 -16856 62157 -16822
rect 62533 -16845 62540 -16697
rect 62556 -16713 62559 -16363
rect 62590 -16679 62593 -16363
rect 62647 -16379 62654 -16371
rect 62596 -16413 62637 -16379
rect 62658 -16413 62709 -16379
rect 63368 -16422 63373 -16406
rect 63391 -16422 63398 -16414
rect 63402 -16422 63407 -16406
rect 63698 -16408 63739 -16374
rect 63743 -16408 63750 -16363
rect 62647 -16462 62654 -16451
rect 62828 -16456 62869 -16422
rect 62900 -16456 62941 -16422
rect 62972 -16456 63013 -16422
rect 63116 -16456 63157 -16422
rect 63188 -16456 63301 -16422
rect 63332 -16456 63373 -16422
rect 62658 -16496 62699 -16462
rect 62647 -16546 62654 -16535
rect 63225 -16539 63266 -16505
rect 62658 -16580 62699 -16546
rect 62647 -16629 62654 -16618
rect 62658 -16663 62699 -16629
rect 62890 -16689 62931 -16655
rect 62935 -16689 62942 -16644
rect 63012 -16706 63017 -16588
rect 63035 -16655 63042 -16644
rect 63046 -16655 63051 -16622
rect 63082 -16655 63087 -16622
rect 63046 -16689 63087 -16655
rect 63091 -16689 63098 -16644
rect 63046 -16740 63051 -16689
rect 63082 -16740 63087 -16689
rect 63116 -16706 63121 -16589
rect 63225 -16623 63266 -16589
rect 63225 -16706 63266 -16672
rect 63368 -16706 63373 -16456
rect 63402 -16456 63443 -16422
rect 63391 -16505 63398 -16494
rect 63402 -16505 63407 -16456
rect 63698 -16491 63739 -16457
rect 63743 -16491 63750 -16446
rect 63402 -16539 63443 -16505
rect 63391 -16589 63398 -16578
rect 63402 -16589 63407 -16539
rect 63551 -16565 63660 -16499
rect 63820 -16507 63825 -16191
rect 63843 -16207 63850 -16199
rect 63854 -16207 63859 -16191
rect 63854 -16241 63895 -16207
rect 63899 -16241 63906 -16199
rect 63843 -16290 63850 -16279
rect 63854 -16290 63859 -16241
rect 63854 -16324 63895 -16290
rect 63899 -16324 63906 -16279
rect 63843 -16374 63850 -16363
rect 63854 -16374 63859 -16324
rect 63854 -16408 63895 -16374
rect 63899 -16408 63906 -16363
rect 63843 -16457 63850 -16446
rect 63854 -16457 63859 -16408
rect 63854 -16491 63895 -16457
rect 63899 -16491 63906 -16446
rect 63843 -16525 63850 -16499
rect 63854 -16541 63859 -16491
rect 63402 -16623 63443 -16589
rect 63763 -16605 63804 -16571
rect 63391 -16672 63398 -16661
rect 63402 -16672 63407 -16623
rect 63402 -16706 63443 -16672
rect 63885 -16673 63892 -16525
rect 63908 -16541 63911 -16191
rect 63942 -16507 63945 -16191
rect 63999 -16207 64006 -16199
rect 63948 -16241 63989 -16207
rect 64010 -16241 64061 -16207
rect 64925 -16231 64966 -16197
rect 65021 -16231 65062 -16197
rect 65117 -16231 65158 -16197
rect 67087 -16207 67094 -16199
rect 64718 -16250 64723 -16234
rect 64741 -16250 64748 -16242
rect 64752 -16250 64757 -16234
rect 63999 -16290 64006 -16279
rect 64178 -16284 64219 -16250
rect 64250 -16284 64291 -16250
rect 64322 -16284 64363 -16250
rect 64466 -16284 64507 -16250
rect 64538 -16284 64651 -16250
rect 64682 -16284 64723 -16250
rect 64010 -16324 64051 -16290
rect 63999 -16374 64006 -16363
rect 64575 -16367 64616 -16333
rect 64010 -16408 64051 -16374
rect 63999 -16457 64006 -16446
rect 64010 -16491 64051 -16457
rect 64240 -16517 64281 -16483
rect 64285 -16517 64292 -16472
rect 64362 -16534 64367 -16416
rect 64385 -16483 64392 -16472
rect 64396 -16483 64401 -16450
rect 64432 -16483 64437 -16450
rect 64396 -16517 64437 -16483
rect 64441 -16517 64448 -16472
rect 64396 -16568 64401 -16517
rect 64432 -16568 64437 -16517
rect 64466 -16534 64471 -16417
rect 64575 -16451 64616 -16417
rect 64575 -16534 64616 -16500
rect 64718 -16534 64723 -16284
rect 64752 -16284 64793 -16250
rect 65279 -16274 65320 -16240
rect 65375 -16274 65416 -16240
rect 65471 -16274 65512 -16240
rect 66978 -16241 67019 -16207
rect 67042 -16241 67094 -16207
rect 67122 -16241 67163 -16207
rect 64741 -16333 64748 -16322
rect 64752 -16333 64757 -16284
rect 64991 -16293 64998 -16285
rect 65091 -16293 65098 -16285
rect 64918 -16327 64987 -16293
rect 64990 -16327 65031 -16293
rect 65102 -16327 65143 -16293
rect 65633 -16317 65674 -16283
rect 65729 -16317 65770 -16283
rect 65825 -16317 65866 -16283
rect 65921 -16317 65962 -16283
rect 66017 -16317 66058 -16283
rect 67042 -16324 67083 -16290
rect 67087 -16324 67094 -16279
rect 64752 -16367 64793 -16333
rect 65345 -16336 65352 -16328
rect 65445 -16336 65452 -16328
rect 64741 -16417 64748 -16406
rect 64752 -16417 64757 -16367
rect 64946 -16410 64987 -16376
rect 64991 -16410 64998 -16365
rect 65091 -16376 65098 -16365
rect 65272 -16370 65341 -16336
rect 65344 -16370 65385 -16336
rect 65456 -16370 65497 -16336
rect 66181 -16360 66222 -16326
rect 66277 -16360 66318 -16326
rect 66373 -16360 66414 -16326
rect 66469 -16360 66510 -16326
rect 66565 -16360 66606 -16326
rect 66661 -16360 66702 -16326
rect 66757 -16360 66798 -16326
rect 65102 -16410 65143 -16376
rect 65735 -16379 65742 -16371
rect 64752 -16451 64793 -16417
rect 64741 -16500 64748 -16489
rect 64752 -16500 64757 -16451
rect 64946 -16494 64987 -16460
rect 64991 -16494 64998 -16449
rect 65091 -16460 65098 -16449
rect 65300 -16453 65341 -16419
rect 65345 -16453 65352 -16408
rect 65445 -16419 65452 -16408
rect 65626 -16413 65667 -16379
rect 65690 -16413 65742 -16379
rect 65770 -16413 65811 -16379
rect 65456 -16453 65497 -16419
rect 65102 -16494 65143 -16460
rect 64752 -16534 64793 -16500
rect 64752 -16568 64757 -16534
rect 63402 -16740 63407 -16706
rect 63698 -16723 63739 -16689
rect 63743 -16723 63750 -16681
rect 63885 -16741 63897 -16673
rect 63926 -16707 63931 -16639
rect 63971 -16671 63976 -16603
rect 64005 -16637 64010 -16571
rect 64946 -16577 64987 -16543
rect 64991 -16577 64998 -16532
rect 65091 -16543 65098 -16532
rect 65300 -16537 65341 -16503
rect 65345 -16537 65352 -16492
rect 65445 -16503 65452 -16492
rect 65690 -16496 65731 -16462
rect 65735 -16496 65742 -16451
rect 65456 -16537 65497 -16503
rect 65102 -16577 65143 -16543
rect 64015 -16621 64056 -16587
rect 64216 -16666 64257 -16632
rect 63985 -16689 63992 -16681
rect 63996 -16723 64037 -16689
rect 64216 -16734 64257 -16700
rect 61149 -16906 61190 -16872
rect 61221 -16906 61262 -16872
rect 61293 -16906 61334 -16872
rect 61606 -16913 61647 -16879
rect 61651 -16913 61658 -16868
rect 61751 -16879 61758 -16868
rect 61762 -16913 61803 -16879
rect 62346 -16895 62387 -16861
rect 62391 -16895 62398 -16853
rect 60240 -16959 60722 -16925
rect 61574 -16949 61615 -16915
rect 61646 -16949 61687 -16915
rect 61960 -16956 62001 -16922
rect 62005 -16956 62012 -16911
rect 62105 -16922 62112 -16911
rect 62533 -16913 62545 -16845
rect 62574 -16879 62579 -16811
rect 62619 -16843 62624 -16775
rect 62653 -16809 62658 -16743
rect 63885 -16753 63892 -16741
rect 64265 -16750 64270 -16616
rect 62663 -16793 62704 -16759
rect 62866 -16838 62907 -16804
rect 62633 -16861 62640 -16853
rect 62644 -16895 62685 -16861
rect 62866 -16906 62907 -16872
rect 62116 -16956 62157 -16922
rect 60240 -16985 60709 -16959
rect 60244 -16993 60451 -16985
rect 60260 -17003 60435 -16993
rect 59986 -17140 60167 -17114
rect 59493 -17174 59534 -17140
rect 59589 -17174 59630 -17140
rect 59685 -17174 59726 -17140
rect 59781 -17174 59822 -17140
rect 59877 -17174 59918 -17140
rect 59973 -17174 60167 -17140
rect 59986 -17200 60167 -17174
rect 60186 -17174 60293 -17050
rect 60445 -17062 60451 -17051
rect 60064 -17870 60105 -17200
rect 60186 -17228 60195 -17174
rect 59871 -17936 60022 -17924
rect 59539 -17970 60022 -17936
rect 59871 -17971 60022 -17970
rect 60052 -17971 60105 -17870
rect 60198 -17971 60239 -17174
rect 60244 -17971 60250 -17174
rect 60456 -17971 60497 -17062
rect 60590 -17971 60631 -16985
rect 60843 -17002 60884 -16968
rect 60939 -17002 60980 -16968
rect 61035 -17002 61076 -16968
rect 61131 -17002 61172 -16968
rect 61227 -17002 61268 -16968
rect 61323 -17002 61364 -16968
rect 61419 -17002 61460 -16968
rect 61928 -16992 61969 -16958
rect 62000 -16992 62041 -16958
rect 62346 -16995 62387 -16961
rect 62391 -16995 62398 -16950
rect 62533 -17001 62540 -16913
rect 62915 -16922 62920 -16788
rect 62633 -16961 62640 -16950
rect 62949 -16956 62954 -16762
rect 62989 -16778 62996 -16767
rect 62985 -16809 62996 -16778
rect 63311 -16796 63352 -16762
rect 62644 -16995 62685 -16961
rect 61581 -17045 61622 -17011
rect 61677 -17045 61718 -17011
rect 61773 -17045 61814 -17011
rect 62282 -17035 62323 -17001
rect 62354 -17035 62395 -17001
rect 62426 -17035 62467 -17001
rect 62498 -17029 62540 -17001
rect 62844 -17025 62885 -16991
rect 62889 -17025 62896 -16980
rect 62985 -16992 62990 -16809
rect 63019 -16995 63024 -16812
rect 62498 -17035 62539 -17029
rect 61935 -17088 61976 -17054
rect 62031 -17088 62072 -17054
rect 62127 -17088 62168 -17054
rect 63031 -17076 63038 -16809
rect 63660 -16819 64053 -16753
rect 64299 -16784 64304 -16590
rect 64339 -16606 64346 -16595
rect 64335 -16637 64346 -16606
rect 64661 -16624 64702 -16590
rect 63047 -16860 63088 -16826
rect 63396 -16830 63413 -16819
rect 63396 -16832 63402 -16830
rect 63047 -16928 63088 -16894
rect 63099 -16995 63104 -16860
rect 63330 -16874 63402 -16832
rect 63458 -16874 64053 -16819
rect 64194 -16853 64235 -16819
rect 64239 -16853 64246 -16808
rect 64335 -16820 64340 -16637
rect 64369 -16823 64374 -16640
rect 63330 -16877 64053 -16874
rect 63133 -16980 63138 -16892
rect 63250 -16942 63291 -16908
rect 63295 -16942 63302 -16900
rect 63131 -16991 63138 -16980
rect 63133 -17025 63138 -16991
rect 63142 -17025 63183 -16991
rect 63250 -17042 63291 -17008
rect 63295 -17042 63302 -16997
rect 63143 -17078 63184 -17044
rect 63215 -17078 63256 -17044
rect 63287 -17078 63328 -17044
rect 62289 -17131 62330 -17097
rect 62385 -17131 62426 -17097
rect 62481 -17131 62522 -17097
rect 62577 -17131 62618 -17097
rect 62673 -17131 62714 -17097
rect 63330 -17114 63481 -16877
rect 63660 -16899 64053 -16877
rect 63584 -16925 64053 -16899
rect 64381 -16904 64388 -16637
rect 64397 -16688 64438 -16654
rect 64397 -16756 64438 -16722
rect 64449 -16823 64454 -16688
rect 65011 -16691 65052 -16657
rect 65063 -16718 65068 -16641
rect 64483 -16808 64488 -16720
rect 64600 -16770 64641 -16736
rect 64645 -16770 64652 -16728
rect 64745 -16740 64752 -16729
rect 64756 -16774 64797 -16740
rect 65097 -16752 65102 -16607
rect 65300 -16620 65341 -16586
rect 65345 -16620 65352 -16575
rect 65445 -16586 65452 -16575
rect 65690 -16580 65731 -16546
rect 65735 -16580 65742 -16535
rect 65456 -16620 65497 -16586
rect 65365 -16734 65406 -16700
rect 65417 -16761 65422 -16684
rect 64481 -16819 64488 -16808
rect 64950 -16813 64991 -16779
rect 64995 -16813 65002 -16771
rect 65095 -16779 65102 -16771
rect 65106 -16813 65147 -16779
rect 65451 -16795 65456 -16650
rect 65690 -16663 65731 -16629
rect 65735 -16663 65742 -16618
rect 65812 -16679 65817 -16363
rect 65835 -16379 65842 -16371
rect 65846 -16379 65851 -16363
rect 65846 -16413 65887 -16379
rect 65891 -16413 65898 -16371
rect 65835 -16462 65842 -16451
rect 65846 -16462 65851 -16413
rect 65846 -16496 65887 -16462
rect 65891 -16496 65898 -16451
rect 65835 -16546 65842 -16535
rect 65846 -16546 65851 -16496
rect 65846 -16580 65887 -16546
rect 65891 -16580 65898 -16535
rect 65835 -16629 65842 -16618
rect 65846 -16629 65851 -16580
rect 65846 -16663 65887 -16629
rect 65891 -16663 65898 -16618
rect 65835 -16697 65842 -16671
rect 65846 -16713 65851 -16663
rect 65755 -16777 65796 -16743
rect 64483 -16853 64488 -16819
rect 64492 -16853 64533 -16819
rect 64600 -16870 64641 -16836
rect 64645 -16870 64652 -16825
rect 64745 -16832 64752 -16821
rect 64756 -16866 64797 -16832
rect 65304 -16856 65345 -16822
rect 65349 -16856 65356 -16814
rect 65449 -16822 65456 -16814
rect 65460 -16856 65501 -16822
rect 65877 -16845 65884 -16697
rect 65900 -16713 65903 -16363
rect 65934 -16679 65937 -16363
rect 65991 -16379 65998 -16371
rect 65940 -16413 65981 -16379
rect 66002 -16413 66053 -16379
rect 66712 -16422 66717 -16406
rect 66735 -16422 66742 -16414
rect 66746 -16422 66751 -16406
rect 67042 -16408 67083 -16374
rect 67087 -16408 67094 -16363
rect 65991 -16462 65998 -16451
rect 66172 -16456 66213 -16422
rect 66244 -16456 66285 -16422
rect 66316 -16456 66357 -16422
rect 66460 -16456 66501 -16422
rect 66532 -16456 66645 -16422
rect 66676 -16456 66717 -16422
rect 66002 -16496 66043 -16462
rect 65991 -16546 65998 -16535
rect 66569 -16539 66610 -16505
rect 66002 -16580 66043 -16546
rect 65991 -16629 65998 -16618
rect 66002 -16663 66043 -16629
rect 66234 -16689 66275 -16655
rect 66279 -16689 66286 -16644
rect 66356 -16706 66361 -16588
rect 66379 -16655 66386 -16644
rect 66390 -16655 66395 -16622
rect 66426 -16655 66431 -16622
rect 66390 -16689 66431 -16655
rect 66435 -16689 66442 -16644
rect 66390 -16740 66395 -16689
rect 66426 -16740 66431 -16689
rect 66460 -16706 66465 -16589
rect 66569 -16623 66610 -16589
rect 66569 -16706 66610 -16672
rect 66712 -16706 66717 -16456
rect 66746 -16456 66787 -16422
rect 66735 -16505 66742 -16494
rect 66746 -16505 66751 -16456
rect 67042 -16491 67083 -16457
rect 67087 -16491 67094 -16446
rect 66746 -16539 66787 -16505
rect 66735 -16589 66742 -16578
rect 66746 -16589 66751 -16539
rect 66895 -16565 67004 -16499
rect 67164 -16507 67169 -16191
rect 67187 -16207 67194 -16199
rect 67198 -16207 67203 -16191
rect 67198 -16241 67239 -16207
rect 67243 -16241 67250 -16199
rect 67187 -16290 67194 -16279
rect 67198 -16290 67203 -16241
rect 67198 -16324 67239 -16290
rect 67243 -16324 67250 -16279
rect 67187 -16374 67194 -16363
rect 67198 -16374 67203 -16324
rect 67198 -16408 67239 -16374
rect 67243 -16408 67250 -16363
rect 67187 -16457 67194 -16446
rect 67198 -16457 67203 -16408
rect 67198 -16491 67239 -16457
rect 67243 -16491 67250 -16446
rect 67187 -16525 67194 -16499
rect 67198 -16541 67203 -16491
rect 66746 -16623 66787 -16589
rect 67107 -16605 67148 -16571
rect 66735 -16672 66742 -16661
rect 66746 -16672 66751 -16623
rect 66746 -16706 66787 -16672
rect 67229 -16673 67236 -16525
rect 67252 -16541 67255 -16191
rect 67286 -16507 67289 -16191
rect 67343 -16207 67350 -16199
rect 67292 -16241 67333 -16207
rect 67354 -16241 67405 -16207
rect 68269 -16231 68310 -16197
rect 68365 -16231 68406 -16197
rect 68461 -16231 68502 -16197
rect 70431 -16207 70438 -16199
rect 68062 -16250 68067 -16234
rect 68085 -16250 68092 -16242
rect 68096 -16250 68101 -16234
rect 67343 -16290 67350 -16279
rect 67522 -16284 67563 -16250
rect 67594 -16284 67635 -16250
rect 67666 -16284 67707 -16250
rect 67810 -16284 67851 -16250
rect 67882 -16284 67995 -16250
rect 68026 -16284 68067 -16250
rect 67354 -16324 67395 -16290
rect 67343 -16374 67350 -16363
rect 67919 -16367 67960 -16333
rect 67354 -16408 67395 -16374
rect 67343 -16457 67350 -16446
rect 67354 -16491 67395 -16457
rect 67584 -16517 67625 -16483
rect 67629 -16517 67636 -16472
rect 67706 -16534 67711 -16416
rect 67729 -16483 67736 -16472
rect 67740 -16483 67745 -16450
rect 67776 -16483 67781 -16450
rect 67740 -16517 67781 -16483
rect 67785 -16517 67792 -16472
rect 67740 -16568 67745 -16517
rect 67776 -16568 67781 -16517
rect 67810 -16534 67815 -16417
rect 67919 -16451 67960 -16417
rect 67919 -16534 67960 -16500
rect 68062 -16534 68067 -16284
rect 68096 -16284 68137 -16250
rect 68623 -16274 68664 -16240
rect 68719 -16274 68760 -16240
rect 68815 -16274 68856 -16240
rect 70322 -16241 70363 -16207
rect 70386 -16241 70438 -16207
rect 70466 -16241 70507 -16207
rect 68085 -16333 68092 -16322
rect 68096 -16333 68101 -16284
rect 68335 -16293 68342 -16285
rect 68435 -16293 68442 -16285
rect 68262 -16327 68331 -16293
rect 68334 -16327 68375 -16293
rect 68446 -16327 68487 -16293
rect 68977 -16317 69018 -16283
rect 69073 -16317 69114 -16283
rect 69169 -16317 69210 -16283
rect 69265 -16317 69306 -16283
rect 69361 -16317 69402 -16283
rect 70386 -16324 70427 -16290
rect 70431 -16324 70438 -16279
rect 68096 -16367 68137 -16333
rect 68689 -16336 68696 -16328
rect 68789 -16336 68796 -16328
rect 68085 -16417 68092 -16406
rect 68096 -16417 68101 -16367
rect 68290 -16410 68331 -16376
rect 68335 -16410 68342 -16365
rect 68435 -16376 68442 -16365
rect 68616 -16370 68685 -16336
rect 68688 -16370 68729 -16336
rect 68800 -16370 68841 -16336
rect 69525 -16360 69566 -16326
rect 69621 -16360 69662 -16326
rect 69717 -16360 69758 -16326
rect 69813 -16360 69854 -16326
rect 69909 -16360 69950 -16326
rect 70005 -16360 70046 -16326
rect 70101 -16360 70142 -16326
rect 68446 -16410 68487 -16376
rect 69079 -16379 69086 -16371
rect 68096 -16451 68137 -16417
rect 68085 -16500 68092 -16489
rect 68096 -16500 68101 -16451
rect 68290 -16494 68331 -16460
rect 68335 -16494 68342 -16449
rect 68435 -16460 68442 -16449
rect 68644 -16453 68685 -16419
rect 68689 -16453 68696 -16408
rect 68789 -16419 68796 -16408
rect 68970 -16413 69011 -16379
rect 69034 -16413 69086 -16379
rect 69114 -16413 69155 -16379
rect 68800 -16453 68841 -16419
rect 68446 -16494 68487 -16460
rect 68096 -16534 68137 -16500
rect 68096 -16568 68101 -16534
rect 66746 -16740 66751 -16706
rect 67042 -16723 67083 -16689
rect 67087 -16723 67094 -16681
rect 67229 -16741 67241 -16673
rect 67270 -16707 67275 -16639
rect 67315 -16671 67320 -16603
rect 67349 -16637 67354 -16571
rect 68290 -16577 68331 -16543
rect 68335 -16577 68342 -16532
rect 68435 -16543 68442 -16532
rect 68644 -16537 68685 -16503
rect 68689 -16537 68696 -16492
rect 68789 -16503 68796 -16492
rect 69034 -16496 69075 -16462
rect 69079 -16496 69086 -16451
rect 68800 -16537 68841 -16503
rect 68446 -16577 68487 -16543
rect 67359 -16621 67400 -16587
rect 67560 -16666 67601 -16632
rect 67329 -16689 67336 -16681
rect 67340 -16723 67381 -16689
rect 67560 -16734 67601 -16700
rect 64493 -16906 64534 -16872
rect 64565 -16906 64606 -16872
rect 64637 -16906 64678 -16872
rect 64950 -16913 64991 -16879
rect 64995 -16913 65002 -16868
rect 65095 -16879 65102 -16868
rect 65106 -16913 65147 -16879
rect 65690 -16895 65731 -16861
rect 65735 -16895 65742 -16853
rect 63584 -16959 64066 -16925
rect 64918 -16949 64959 -16915
rect 64990 -16949 65031 -16915
rect 65304 -16956 65345 -16922
rect 65349 -16956 65356 -16911
rect 65449 -16922 65456 -16911
rect 65877 -16913 65889 -16845
rect 65918 -16879 65923 -16811
rect 65963 -16843 65968 -16775
rect 65997 -16809 66002 -16743
rect 67229 -16753 67236 -16741
rect 67609 -16750 67614 -16616
rect 66007 -16793 66048 -16759
rect 66210 -16838 66251 -16804
rect 65977 -16861 65984 -16853
rect 65988 -16895 66029 -16861
rect 66210 -16906 66251 -16872
rect 65460 -16956 65501 -16922
rect 63584 -16985 64053 -16959
rect 63588 -16993 63795 -16985
rect 63604 -17003 63779 -16993
rect 63330 -17140 63511 -17114
rect 62837 -17174 62878 -17140
rect 62933 -17174 62974 -17140
rect 63029 -17174 63070 -17140
rect 63125 -17174 63166 -17140
rect 63221 -17174 63262 -17140
rect 63317 -17174 63511 -17140
rect 63330 -17200 63511 -17174
rect 63530 -17174 63637 -17050
rect 63789 -17062 63795 -17051
rect 63408 -17870 63449 -17200
rect 63530 -17228 63539 -17174
rect 63215 -17936 63366 -17924
rect 62883 -17970 63366 -17936
rect 63215 -17971 63366 -17970
rect 63396 -17971 63449 -17870
rect 63542 -17971 63583 -17174
rect 63588 -17971 63594 -17174
rect 63800 -17971 63841 -17062
rect 63934 -17971 63975 -16985
rect 64187 -17002 64228 -16968
rect 64283 -17002 64324 -16968
rect 64379 -17002 64420 -16968
rect 64475 -17002 64516 -16968
rect 64571 -17002 64612 -16968
rect 64667 -17002 64708 -16968
rect 64763 -17002 64804 -16968
rect 65272 -16992 65313 -16958
rect 65344 -16992 65385 -16958
rect 65690 -16995 65731 -16961
rect 65735 -16995 65742 -16950
rect 65877 -17001 65884 -16913
rect 66259 -16922 66264 -16788
rect 65977 -16961 65984 -16950
rect 66293 -16956 66298 -16762
rect 66333 -16778 66340 -16767
rect 66329 -16809 66340 -16778
rect 66655 -16796 66696 -16762
rect 65988 -16995 66029 -16961
rect 64925 -17045 64966 -17011
rect 65021 -17045 65062 -17011
rect 65117 -17045 65158 -17011
rect 65626 -17035 65667 -17001
rect 65698 -17035 65739 -17001
rect 65770 -17035 65811 -17001
rect 65842 -17029 65884 -17001
rect 66188 -17025 66229 -16991
rect 66233 -17025 66240 -16980
rect 66329 -16992 66334 -16809
rect 66363 -16995 66368 -16812
rect 65842 -17035 65883 -17029
rect 65279 -17088 65320 -17054
rect 65375 -17088 65416 -17054
rect 65471 -17088 65512 -17054
rect 66375 -17076 66382 -16809
rect 67004 -16819 67397 -16753
rect 67643 -16784 67648 -16590
rect 67683 -16606 67690 -16595
rect 67679 -16637 67690 -16606
rect 68005 -16624 68046 -16590
rect 66391 -16860 66432 -16826
rect 66740 -16830 66757 -16819
rect 66740 -16832 66746 -16830
rect 66391 -16928 66432 -16894
rect 66443 -16995 66448 -16860
rect 66674 -16874 66746 -16832
rect 66802 -16874 67397 -16819
rect 67538 -16853 67579 -16819
rect 67583 -16853 67590 -16808
rect 67679 -16820 67684 -16637
rect 67713 -16823 67718 -16640
rect 66674 -16877 67397 -16874
rect 66477 -16980 66482 -16892
rect 66594 -16942 66635 -16908
rect 66639 -16942 66646 -16900
rect 66475 -16991 66482 -16980
rect 66477 -17025 66482 -16991
rect 66486 -17025 66527 -16991
rect 66594 -17042 66635 -17008
rect 66639 -17042 66646 -16997
rect 66487 -17078 66528 -17044
rect 66559 -17078 66600 -17044
rect 66631 -17078 66672 -17044
rect 65633 -17131 65674 -17097
rect 65729 -17131 65770 -17097
rect 65825 -17131 65866 -17097
rect 65921 -17131 65962 -17097
rect 66017 -17131 66058 -17097
rect 66674 -17114 66825 -16877
rect 67004 -16899 67397 -16877
rect 66928 -16925 67397 -16899
rect 67725 -16904 67732 -16637
rect 67741 -16688 67782 -16654
rect 67741 -16756 67782 -16722
rect 67793 -16823 67798 -16688
rect 68355 -16691 68396 -16657
rect 68407 -16718 68412 -16641
rect 67827 -16808 67832 -16720
rect 67944 -16770 67985 -16736
rect 67989 -16770 67996 -16728
rect 68089 -16740 68096 -16729
rect 68100 -16774 68141 -16740
rect 68441 -16752 68446 -16607
rect 68644 -16620 68685 -16586
rect 68689 -16620 68696 -16575
rect 68789 -16586 68796 -16575
rect 69034 -16580 69075 -16546
rect 69079 -16580 69086 -16535
rect 68800 -16620 68841 -16586
rect 68709 -16734 68750 -16700
rect 68761 -16761 68766 -16684
rect 67825 -16819 67832 -16808
rect 68294 -16813 68335 -16779
rect 68339 -16813 68346 -16771
rect 68439 -16779 68446 -16771
rect 68450 -16813 68491 -16779
rect 68795 -16795 68800 -16650
rect 69034 -16663 69075 -16629
rect 69079 -16663 69086 -16618
rect 69156 -16679 69161 -16363
rect 69179 -16379 69186 -16371
rect 69190 -16379 69195 -16363
rect 69190 -16413 69231 -16379
rect 69235 -16413 69242 -16371
rect 69179 -16462 69186 -16451
rect 69190 -16462 69195 -16413
rect 69190 -16496 69231 -16462
rect 69235 -16496 69242 -16451
rect 69179 -16546 69186 -16535
rect 69190 -16546 69195 -16496
rect 69190 -16580 69231 -16546
rect 69235 -16580 69242 -16535
rect 69179 -16629 69186 -16618
rect 69190 -16629 69195 -16580
rect 69190 -16663 69231 -16629
rect 69235 -16663 69242 -16618
rect 69179 -16697 69186 -16671
rect 69190 -16713 69195 -16663
rect 69099 -16777 69140 -16743
rect 67827 -16853 67832 -16819
rect 67836 -16853 67877 -16819
rect 67944 -16870 67985 -16836
rect 67989 -16870 67996 -16825
rect 68089 -16832 68096 -16821
rect 68100 -16866 68141 -16832
rect 68648 -16856 68689 -16822
rect 68693 -16856 68700 -16814
rect 68793 -16822 68800 -16814
rect 68804 -16856 68845 -16822
rect 69221 -16845 69228 -16697
rect 69244 -16713 69247 -16363
rect 69278 -16679 69281 -16363
rect 69335 -16379 69342 -16371
rect 69284 -16413 69325 -16379
rect 69346 -16413 69397 -16379
rect 70056 -16422 70061 -16406
rect 70079 -16422 70086 -16414
rect 70090 -16422 70095 -16406
rect 70386 -16408 70427 -16374
rect 70431 -16408 70438 -16363
rect 69335 -16462 69342 -16451
rect 69516 -16456 69557 -16422
rect 69588 -16456 69629 -16422
rect 69660 -16456 69701 -16422
rect 69804 -16456 69845 -16422
rect 69876 -16456 69989 -16422
rect 70020 -16456 70061 -16422
rect 69346 -16496 69387 -16462
rect 69335 -16546 69342 -16535
rect 69913 -16539 69954 -16505
rect 69346 -16580 69387 -16546
rect 69335 -16629 69342 -16618
rect 69346 -16663 69387 -16629
rect 69578 -16689 69619 -16655
rect 69623 -16689 69630 -16644
rect 69700 -16706 69705 -16588
rect 69723 -16655 69730 -16644
rect 69734 -16655 69739 -16622
rect 69770 -16655 69775 -16622
rect 69734 -16689 69775 -16655
rect 69779 -16689 69786 -16644
rect 69734 -16740 69739 -16689
rect 69770 -16740 69775 -16689
rect 69804 -16706 69809 -16589
rect 69913 -16623 69954 -16589
rect 69913 -16706 69954 -16672
rect 70056 -16706 70061 -16456
rect 70090 -16456 70131 -16422
rect 70079 -16505 70086 -16494
rect 70090 -16505 70095 -16456
rect 70386 -16491 70427 -16457
rect 70431 -16491 70438 -16446
rect 70090 -16539 70131 -16505
rect 70079 -16589 70086 -16578
rect 70090 -16589 70095 -16539
rect 70239 -16565 70348 -16499
rect 70508 -16507 70513 -16191
rect 70531 -16207 70538 -16199
rect 70542 -16207 70547 -16191
rect 70542 -16241 70583 -16207
rect 70587 -16241 70594 -16199
rect 70531 -16290 70538 -16279
rect 70542 -16290 70547 -16241
rect 70542 -16324 70583 -16290
rect 70587 -16324 70594 -16279
rect 70531 -16374 70538 -16363
rect 70542 -16374 70547 -16324
rect 70542 -16408 70583 -16374
rect 70587 -16408 70594 -16363
rect 70531 -16457 70538 -16446
rect 70542 -16457 70547 -16408
rect 70542 -16491 70583 -16457
rect 70587 -16491 70594 -16446
rect 70531 -16525 70538 -16499
rect 70542 -16541 70547 -16491
rect 70090 -16623 70131 -16589
rect 70451 -16605 70492 -16571
rect 70079 -16672 70086 -16661
rect 70090 -16672 70095 -16623
rect 70090 -16706 70131 -16672
rect 70573 -16673 70580 -16525
rect 70596 -16541 70599 -16191
rect 70630 -16507 70633 -16191
rect 70687 -16207 70694 -16199
rect 70636 -16241 70677 -16207
rect 70698 -16241 70749 -16207
rect 71613 -16231 71654 -16197
rect 71709 -16231 71750 -16197
rect 71805 -16231 71846 -16197
rect 73775 -16207 73782 -16199
rect 71406 -16250 71411 -16234
rect 71429 -16250 71436 -16242
rect 71440 -16250 71445 -16234
rect 70687 -16290 70694 -16279
rect 70866 -16284 70907 -16250
rect 70938 -16284 70979 -16250
rect 71010 -16284 71051 -16250
rect 71154 -16284 71195 -16250
rect 71226 -16284 71339 -16250
rect 71370 -16284 71411 -16250
rect 70698 -16324 70739 -16290
rect 70687 -16374 70694 -16363
rect 71263 -16367 71304 -16333
rect 70698 -16408 70739 -16374
rect 70687 -16457 70694 -16446
rect 70698 -16491 70739 -16457
rect 70928 -16517 70969 -16483
rect 70973 -16517 70980 -16472
rect 71050 -16534 71055 -16416
rect 71073 -16483 71080 -16472
rect 71084 -16483 71089 -16450
rect 71120 -16483 71125 -16450
rect 71084 -16517 71125 -16483
rect 71129 -16517 71136 -16472
rect 71084 -16568 71089 -16517
rect 71120 -16568 71125 -16517
rect 71154 -16534 71159 -16417
rect 71263 -16451 71304 -16417
rect 71263 -16534 71304 -16500
rect 71406 -16534 71411 -16284
rect 71440 -16284 71481 -16250
rect 71967 -16274 72008 -16240
rect 72063 -16274 72104 -16240
rect 72159 -16274 72200 -16240
rect 73666 -16241 73707 -16207
rect 73730 -16241 73782 -16207
rect 73810 -16241 73851 -16207
rect 71429 -16333 71436 -16322
rect 71440 -16333 71445 -16284
rect 71679 -16293 71686 -16285
rect 71779 -16293 71786 -16285
rect 71606 -16327 71675 -16293
rect 71678 -16327 71719 -16293
rect 71790 -16327 71831 -16293
rect 72321 -16317 72362 -16283
rect 72417 -16317 72458 -16283
rect 72513 -16317 72554 -16283
rect 72609 -16317 72650 -16283
rect 72705 -16317 72746 -16283
rect 73730 -16324 73771 -16290
rect 73775 -16324 73782 -16279
rect 71440 -16367 71481 -16333
rect 72033 -16336 72040 -16328
rect 72133 -16336 72140 -16328
rect 71429 -16417 71436 -16406
rect 71440 -16417 71445 -16367
rect 71634 -16410 71675 -16376
rect 71679 -16410 71686 -16365
rect 71779 -16376 71786 -16365
rect 71960 -16370 72029 -16336
rect 72032 -16370 72073 -16336
rect 72144 -16370 72185 -16336
rect 72869 -16360 72910 -16326
rect 72965 -16360 73006 -16326
rect 73061 -16360 73102 -16326
rect 73157 -16360 73198 -16326
rect 73253 -16360 73294 -16326
rect 73349 -16360 73390 -16326
rect 73445 -16360 73486 -16326
rect 71790 -16410 71831 -16376
rect 72423 -16379 72430 -16371
rect 71440 -16451 71481 -16417
rect 71429 -16500 71436 -16489
rect 71440 -16500 71445 -16451
rect 71634 -16494 71675 -16460
rect 71679 -16494 71686 -16449
rect 71779 -16460 71786 -16449
rect 71988 -16453 72029 -16419
rect 72033 -16453 72040 -16408
rect 72133 -16419 72140 -16408
rect 72314 -16413 72355 -16379
rect 72378 -16413 72430 -16379
rect 72458 -16413 72499 -16379
rect 72144 -16453 72185 -16419
rect 71790 -16494 71831 -16460
rect 71440 -16534 71481 -16500
rect 71440 -16568 71445 -16534
rect 70090 -16740 70095 -16706
rect 70386 -16723 70427 -16689
rect 70431 -16723 70438 -16681
rect 70573 -16741 70585 -16673
rect 70614 -16707 70619 -16639
rect 70659 -16671 70664 -16603
rect 70693 -16637 70698 -16571
rect 71634 -16577 71675 -16543
rect 71679 -16577 71686 -16532
rect 71779 -16543 71786 -16532
rect 71988 -16537 72029 -16503
rect 72033 -16537 72040 -16492
rect 72133 -16503 72140 -16492
rect 72378 -16496 72419 -16462
rect 72423 -16496 72430 -16451
rect 72144 -16537 72185 -16503
rect 71790 -16577 71831 -16543
rect 70703 -16621 70744 -16587
rect 70904 -16666 70945 -16632
rect 70673 -16689 70680 -16681
rect 70684 -16723 70725 -16689
rect 70904 -16734 70945 -16700
rect 67837 -16906 67878 -16872
rect 67909 -16906 67950 -16872
rect 67981 -16906 68022 -16872
rect 68294 -16913 68335 -16879
rect 68339 -16913 68346 -16868
rect 68439 -16879 68446 -16868
rect 68450 -16913 68491 -16879
rect 69034 -16895 69075 -16861
rect 69079 -16895 69086 -16853
rect 66928 -16959 67410 -16925
rect 68262 -16949 68303 -16915
rect 68334 -16949 68375 -16915
rect 68648 -16956 68689 -16922
rect 68693 -16956 68700 -16911
rect 68793 -16922 68800 -16911
rect 69221 -16913 69233 -16845
rect 69262 -16879 69267 -16811
rect 69307 -16843 69312 -16775
rect 69341 -16809 69346 -16743
rect 70573 -16753 70580 -16741
rect 70953 -16750 70958 -16616
rect 69351 -16793 69392 -16759
rect 69554 -16838 69595 -16804
rect 69321 -16861 69328 -16853
rect 69332 -16895 69373 -16861
rect 69554 -16906 69595 -16872
rect 68804 -16956 68845 -16922
rect 66928 -16985 67397 -16959
rect 66932 -16993 67139 -16985
rect 66948 -17003 67123 -16993
rect 66674 -17140 66855 -17114
rect 66181 -17174 66222 -17140
rect 66277 -17174 66318 -17140
rect 66373 -17174 66414 -17140
rect 66469 -17174 66510 -17140
rect 66565 -17174 66606 -17140
rect 66661 -17174 66855 -17140
rect 66674 -17200 66855 -17174
rect 66874 -17174 66981 -17050
rect 67133 -17062 67139 -17051
rect 66752 -17870 66793 -17200
rect 66874 -17228 66883 -17174
rect 66559 -17936 66710 -17924
rect 66227 -17970 66710 -17936
rect 66559 -17971 66710 -17970
rect 66740 -17971 66793 -17870
rect 66886 -17971 66927 -17174
rect 66932 -17971 66938 -17174
rect 67144 -17971 67185 -17062
rect 67278 -17971 67319 -16985
rect 67531 -17002 67572 -16968
rect 67627 -17002 67668 -16968
rect 67723 -17002 67764 -16968
rect 67819 -17002 67860 -16968
rect 67915 -17002 67956 -16968
rect 68011 -17002 68052 -16968
rect 68107 -17002 68148 -16968
rect 68616 -16992 68657 -16958
rect 68688 -16992 68729 -16958
rect 69034 -16995 69075 -16961
rect 69079 -16995 69086 -16950
rect 69221 -17001 69228 -16913
rect 69603 -16922 69608 -16788
rect 69321 -16961 69328 -16950
rect 69637 -16956 69642 -16762
rect 69677 -16778 69684 -16767
rect 69673 -16809 69684 -16778
rect 69999 -16796 70040 -16762
rect 69332 -16995 69373 -16961
rect 68269 -17045 68310 -17011
rect 68365 -17045 68406 -17011
rect 68461 -17045 68502 -17011
rect 68970 -17035 69011 -17001
rect 69042 -17035 69083 -17001
rect 69114 -17035 69155 -17001
rect 69186 -17029 69228 -17001
rect 69532 -17025 69573 -16991
rect 69577 -17025 69584 -16980
rect 69673 -16992 69678 -16809
rect 69707 -16995 69712 -16812
rect 69186 -17035 69227 -17029
rect 68623 -17088 68664 -17054
rect 68719 -17088 68760 -17054
rect 68815 -17088 68856 -17054
rect 69719 -17076 69726 -16809
rect 70348 -16819 70741 -16753
rect 70987 -16784 70992 -16590
rect 71027 -16606 71034 -16595
rect 71023 -16637 71034 -16606
rect 71349 -16624 71390 -16590
rect 69735 -16860 69776 -16826
rect 70084 -16830 70101 -16819
rect 70084 -16832 70090 -16830
rect 69735 -16928 69776 -16894
rect 69787 -16995 69792 -16860
rect 70018 -16874 70090 -16832
rect 70146 -16874 70741 -16819
rect 70882 -16853 70923 -16819
rect 70927 -16853 70934 -16808
rect 71023 -16820 71028 -16637
rect 71057 -16823 71062 -16640
rect 70018 -16877 70741 -16874
rect 69821 -16980 69826 -16892
rect 69938 -16942 69979 -16908
rect 69983 -16942 69990 -16900
rect 69819 -16991 69826 -16980
rect 69821 -17025 69826 -16991
rect 69830 -17025 69871 -16991
rect 69938 -17042 69979 -17008
rect 69983 -17042 69990 -16997
rect 69831 -17078 69872 -17044
rect 69903 -17078 69944 -17044
rect 69975 -17078 70016 -17044
rect 68977 -17131 69018 -17097
rect 69073 -17131 69114 -17097
rect 69169 -17131 69210 -17097
rect 69265 -17131 69306 -17097
rect 69361 -17131 69402 -17097
rect 70018 -17114 70169 -16877
rect 70348 -16899 70741 -16877
rect 70272 -16925 70741 -16899
rect 71069 -16904 71076 -16637
rect 71085 -16688 71126 -16654
rect 71085 -16756 71126 -16722
rect 71137 -16823 71142 -16688
rect 71699 -16691 71740 -16657
rect 71751 -16718 71756 -16641
rect 71171 -16808 71176 -16720
rect 71288 -16770 71329 -16736
rect 71333 -16770 71340 -16728
rect 71433 -16740 71440 -16729
rect 71444 -16774 71485 -16740
rect 71785 -16752 71790 -16607
rect 71988 -16620 72029 -16586
rect 72033 -16620 72040 -16575
rect 72133 -16586 72140 -16575
rect 72378 -16580 72419 -16546
rect 72423 -16580 72430 -16535
rect 72144 -16620 72185 -16586
rect 72053 -16734 72094 -16700
rect 72105 -16761 72110 -16684
rect 71169 -16819 71176 -16808
rect 71638 -16813 71679 -16779
rect 71683 -16813 71690 -16771
rect 71783 -16779 71790 -16771
rect 71794 -16813 71835 -16779
rect 72139 -16795 72144 -16650
rect 72378 -16663 72419 -16629
rect 72423 -16663 72430 -16618
rect 72500 -16679 72505 -16363
rect 72523 -16379 72530 -16371
rect 72534 -16379 72539 -16363
rect 72534 -16413 72575 -16379
rect 72579 -16413 72586 -16371
rect 72523 -16462 72530 -16451
rect 72534 -16462 72539 -16413
rect 72534 -16496 72575 -16462
rect 72579 -16496 72586 -16451
rect 72523 -16546 72530 -16535
rect 72534 -16546 72539 -16496
rect 72534 -16580 72575 -16546
rect 72579 -16580 72586 -16535
rect 72523 -16629 72530 -16618
rect 72534 -16629 72539 -16580
rect 72534 -16663 72575 -16629
rect 72579 -16663 72586 -16618
rect 72523 -16697 72530 -16671
rect 72534 -16713 72539 -16663
rect 72443 -16777 72484 -16743
rect 71171 -16853 71176 -16819
rect 71180 -16853 71221 -16819
rect 71288 -16870 71329 -16836
rect 71333 -16870 71340 -16825
rect 71433 -16832 71440 -16821
rect 71444 -16866 71485 -16832
rect 71992 -16856 72033 -16822
rect 72037 -16856 72044 -16814
rect 72137 -16822 72144 -16814
rect 72148 -16856 72189 -16822
rect 72565 -16845 72572 -16697
rect 72588 -16713 72591 -16363
rect 72622 -16679 72625 -16363
rect 72679 -16379 72686 -16371
rect 72628 -16413 72669 -16379
rect 72690 -16413 72741 -16379
rect 73400 -16422 73405 -16406
rect 73423 -16422 73430 -16414
rect 73434 -16422 73439 -16406
rect 73730 -16408 73771 -16374
rect 73775 -16408 73782 -16363
rect 72679 -16462 72686 -16451
rect 72860 -16456 72901 -16422
rect 72932 -16456 72973 -16422
rect 73004 -16456 73045 -16422
rect 73148 -16456 73189 -16422
rect 73220 -16456 73333 -16422
rect 73364 -16456 73405 -16422
rect 72690 -16496 72731 -16462
rect 72679 -16546 72686 -16535
rect 73257 -16539 73298 -16505
rect 72690 -16580 72731 -16546
rect 72679 -16629 72686 -16618
rect 72690 -16663 72731 -16629
rect 72922 -16689 72963 -16655
rect 72967 -16689 72974 -16644
rect 73044 -16706 73049 -16588
rect 73067 -16655 73074 -16644
rect 73078 -16655 73083 -16622
rect 73114 -16655 73119 -16622
rect 73078 -16689 73119 -16655
rect 73123 -16689 73130 -16644
rect 73078 -16740 73083 -16689
rect 73114 -16740 73119 -16689
rect 73148 -16706 73153 -16589
rect 73257 -16623 73298 -16589
rect 73257 -16706 73298 -16672
rect 73400 -16706 73405 -16456
rect 73434 -16456 73475 -16422
rect 73423 -16505 73430 -16494
rect 73434 -16505 73439 -16456
rect 73730 -16491 73771 -16457
rect 73775 -16491 73782 -16446
rect 73434 -16539 73475 -16505
rect 73423 -16589 73430 -16578
rect 73434 -16589 73439 -16539
rect 73583 -16565 73692 -16499
rect 73852 -16507 73857 -16191
rect 73875 -16207 73882 -16199
rect 73886 -16207 73891 -16191
rect 73886 -16241 73927 -16207
rect 73931 -16241 73938 -16199
rect 73875 -16290 73882 -16279
rect 73886 -16290 73891 -16241
rect 73886 -16324 73927 -16290
rect 73931 -16324 73938 -16279
rect 73875 -16374 73882 -16363
rect 73886 -16374 73891 -16324
rect 73886 -16408 73927 -16374
rect 73931 -16408 73938 -16363
rect 73875 -16457 73882 -16446
rect 73886 -16457 73891 -16408
rect 73886 -16491 73927 -16457
rect 73931 -16491 73938 -16446
rect 73875 -16525 73882 -16499
rect 73886 -16541 73891 -16491
rect 73434 -16623 73475 -16589
rect 73795 -16605 73836 -16571
rect 73423 -16672 73430 -16661
rect 73434 -16672 73439 -16623
rect 73434 -16706 73475 -16672
rect 73917 -16673 73924 -16525
rect 73940 -16541 73943 -16191
rect 73974 -16507 73977 -16191
rect 74031 -16207 74038 -16199
rect 73980 -16241 74021 -16207
rect 74042 -16241 74093 -16207
rect 74957 -16231 74998 -16197
rect 75053 -16231 75094 -16197
rect 75149 -16231 75190 -16197
rect 77119 -16207 77126 -16199
rect 74750 -16250 74755 -16234
rect 74773 -16250 74780 -16242
rect 74784 -16250 74789 -16234
rect 74031 -16290 74038 -16279
rect 74210 -16284 74251 -16250
rect 74282 -16284 74323 -16250
rect 74354 -16284 74395 -16250
rect 74498 -16284 74539 -16250
rect 74570 -16284 74683 -16250
rect 74714 -16284 74755 -16250
rect 74042 -16324 74083 -16290
rect 74031 -16374 74038 -16363
rect 74607 -16367 74648 -16333
rect 74042 -16408 74083 -16374
rect 74031 -16457 74038 -16446
rect 74042 -16491 74083 -16457
rect 74272 -16517 74313 -16483
rect 74317 -16517 74324 -16472
rect 74394 -16534 74399 -16416
rect 74417 -16483 74424 -16472
rect 74428 -16483 74433 -16450
rect 74464 -16483 74469 -16450
rect 74428 -16517 74469 -16483
rect 74473 -16517 74480 -16472
rect 74428 -16568 74433 -16517
rect 74464 -16568 74469 -16517
rect 74498 -16534 74503 -16417
rect 74607 -16451 74648 -16417
rect 74607 -16534 74648 -16500
rect 74750 -16534 74755 -16284
rect 74784 -16284 74825 -16250
rect 75311 -16274 75352 -16240
rect 75407 -16274 75448 -16240
rect 75503 -16274 75544 -16240
rect 77010 -16241 77051 -16207
rect 77074 -16241 77126 -16207
rect 77154 -16241 77195 -16207
rect 74773 -16333 74780 -16322
rect 74784 -16333 74789 -16284
rect 75023 -16293 75030 -16285
rect 75123 -16293 75130 -16285
rect 74950 -16327 75019 -16293
rect 75022 -16327 75063 -16293
rect 75134 -16327 75175 -16293
rect 75665 -16317 75706 -16283
rect 75761 -16317 75802 -16283
rect 75857 -16317 75898 -16283
rect 75953 -16317 75994 -16283
rect 76049 -16317 76090 -16283
rect 77074 -16324 77115 -16290
rect 77119 -16324 77126 -16279
rect 74784 -16367 74825 -16333
rect 75377 -16336 75384 -16328
rect 75477 -16336 75484 -16328
rect 74773 -16417 74780 -16406
rect 74784 -16417 74789 -16367
rect 74978 -16410 75019 -16376
rect 75023 -16410 75030 -16365
rect 75123 -16376 75130 -16365
rect 75304 -16370 75373 -16336
rect 75376 -16370 75417 -16336
rect 75488 -16370 75529 -16336
rect 76213 -16360 76254 -16326
rect 76309 -16360 76350 -16326
rect 76405 -16360 76446 -16326
rect 76501 -16360 76542 -16326
rect 76597 -16360 76638 -16326
rect 76693 -16360 76734 -16326
rect 76789 -16360 76830 -16326
rect 75134 -16410 75175 -16376
rect 75767 -16379 75774 -16371
rect 74784 -16451 74825 -16417
rect 74773 -16500 74780 -16489
rect 74784 -16500 74789 -16451
rect 74978 -16494 75019 -16460
rect 75023 -16494 75030 -16449
rect 75123 -16460 75130 -16449
rect 75332 -16453 75373 -16419
rect 75377 -16453 75384 -16408
rect 75477 -16419 75484 -16408
rect 75658 -16413 75699 -16379
rect 75722 -16413 75774 -16379
rect 75802 -16413 75843 -16379
rect 75488 -16453 75529 -16419
rect 75134 -16494 75175 -16460
rect 74784 -16534 74825 -16500
rect 74784 -16568 74789 -16534
rect 73434 -16740 73439 -16706
rect 73730 -16723 73771 -16689
rect 73775 -16723 73782 -16681
rect 73917 -16741 73929 -16673
rect 73958 -16707 73963 -16639
rect 74003 -16671 74008 -16603
rect 74037 -16637 74042 -16571
rect 74978 -16577 75019 -16543
rect 75023 -16577 75030 -16532
rect 75123 -16543 75130 -16532
rect 75332 -16537 75373 -16503
rect 75377 -16537 75384 -16492
rect 75477 -16503 75484 -16492
rect 75722 -16496 75763 -16462
rect 75767 -16496 75774 -16451
rect 75488 -16537 75529 -16503
rect 75134 -16577 75175 -16543
rect 74047 -16621 74088 -16587
rect 74248 -16666 74289 -16632
rect 74017 -16689 74024 -16681
rect 74028 -16723 74069 -16689
rect 74248 -16734 74289 -16700
rect 71181 -16906 71222 -16872
rect 71253 -16906 71294 -16872
rect 71325 -16906 71366 -16872
rect 71638 -16913 71679 -16879
rect 71683 -16913 71690 -16868
rect 71783 -16879 71790 -16868
rect 71794 -16913 71835 -16879
rect 72378 -16895 72419 -16861
rect 72423 -16895 72430 -16853
rect 70272 -16959 70754 -16925
rect 71606 -16949 71647 -16915
rect 71678 -16949 71719 -16915
rect 71992 -16956 72033 -16922
rect 72037 -16956 72044 -16911
rect 72137 -16922 72144 -16911
rect 72565 -16913 72577 -16845
rect 72606 -16879 72611 -16811
rect 72651 -16843 72656 -16775
rect 72685 -16809 72690 -16743
rect 73917 -16753 73924 -16741
rect 74297 -16750 74302 -16616
rect 72695 -16793 72736 -16759
rect 72898 -16838 72939 -16804
rect 72665 -16861 72672 -16853
rect 72676 -16895 72717 -16861
rect 72898 -16906 72939 -16872
rect 72148 -16956 72189 -16922
rect 70272 -16985 70741 -16959
rect 70276 -16993 70483 -16985
rect 70292 -17003 70467 -16993
rect 70018 -17140 70199 -17114
rect 69525 -17174 69566 -17140
rect 69621 -17174 69662 -17140
rect 69717 -17174 69758 -17140
rect 69813 -17174 69854 -17140
rect 69909 -17174 69950 -17140
rect 70005 -17174 70199 -17140
rect 70018 -17200 70199 -17174
rect 70218 -17174 70325 -17050
rect 70477 -17062 70483 -17051
rect 70096 -17870 70137 -17200
rect 70218 -17228 70227 -17174
rect 69903 -17936 70054 -17924
rect 69571 -17970 70054 -17936
rect 69903 -17971 70054 -17970
rect 70084 -17971 70137 -17870
rect 70230 -17971 70271 -17174
rect 70276 -17971 70282 -17174
rect 70488 -17971 70529 -17062
rect 70622 -17971 70663 -16985
rect 70875 -17002 70916 -16968
rect 70971 -17002 71012 -16968
rect 71067 -17002 71108 -16968
rect 71163 -17002 71204 -16968
rect 71259 -17002 71300 -16968
rect 71355 -17002 71396 -16968
rect 71451 -17002 71492 -16968
rect 71960 -16992 72001 -16958
rect 72032 -16992 72073 -16958
rect 72378 -16995 72419 -16961
rect 72423 -16995 72430 -16950
rect 72565 -17001 72572 -16913
rect 72947 -16922 72952 -16788
rect 72665 -16961 72672 -16950
rect 72981 -16956 72986 -16762
rect 73021 -16778 73028 -16767
rect 73017 -16809 73028 -16778
rect 73343 -16796 73384 -16762
rect 72676 -16995 72717 -16961
rect 71613 -17045 71654 -17011
rect 71709 -17045 71750 -17011
rect 71805 -17045 71846 -17011
rect 72314 -17035 72355 -17001
rect 72386 -17035 72427 -17001
rect 72458 -17035 72499 -17001
rect 72530 -17029 72572 -17001
rect 72876 -17025 72917 -16991
rect 72921 -17025 72928 -16980
rect 73017 -16992 73022 -16809
rect 73051 -16995 73056 -16812
rect 72530 -17035 72571 -17029
rect 71967 -17088 72008 -17054
rect 72063 -17088 72104 -17054
rect 72159 -17088 72200 -17054
rect 73063 -17076 73070 -16809
rect 73692 -16819 74085 -16753
rect 74331 -16784 74336 -16590
rect 74371 -16606 74378 -16595
rect 74367 -16637 74378 -16606
rect 74693 -16624 74734 -16590
rect 73079 -16860 73120 -16826
rect 73428 -16830 73445 -16819
rect 73428 -16832 73434 -16830
rect 73079 -16928 73120 -16894
rect 73131 -16995 73136 -16860
rect 73362 -16874 73434 -16832
rect 73490 -16874 74085 -16819
rect 74226 -16853 74267 -16819
rect 74271 -16853 74278 -16808
rect 74367 -16820 74372 -16637
rect 74401 -16823 74406 -16640
rect 73362 -16877 74085 -16874
rect 73165 -16980 73170 -16892
rect 73282 -16942 73323 -16908
rect 73327 -16942 73334 -16900
rect 73163 -16991 73170 -16980
rect 73165 -17025 73170 -16991
rect 73174 -17025 73215 -16991
rect 73282 -17042 73323 -17008
rect 73327 -17042 73334 -16997
rect 73175 -17078 73216 -17044
rect 73247 -17078 73288 -17044
rect 73319 -17078 73360 -17044
rect 72321 -17131 72362 -17097
rect 72417 -17131 72458 -17097
rect 72513 -17131 72554 -17097
rect 72609 -17131 72650 -17097
rect 72705 -17131 72746 -17097
rect 73362 -17114 73513 -16877
rect 73692 -16899 74085 -16877
rect 73616 -16925 74085 -16899
rect 74413 -16904 74420 -16637
rect 74429 -16688 74470 -16654
rect 74429 -16756 74470 -16722
rect 74481 -16823 74486 -16688
rect 75043 -16691 75084 -16657
rect 75095 -16718 75100 -16641
rect 74515 -16808 74520 -16720
rect 74632 -16770 74673 -16736
rect 74677 -16770 74684 -16728
rect 74777 -16740 74784 -16729
rect 74788 -16774 74829 -16740
rect 75129 -16752 75134 -16607
rect 75332 -16620 75373 -16586
rect 75377 -16620 75384 -16575
rect 75477 -16586 75484 -16575
rect 75722 -16580 75763 -16546
rect 75767 -16580 75774 -16535
rect 75488 -16620 75529 -16586
rect 75397 -16734 75438 -16700
rect 75449 -16761 75454 -16684
rect 74513 -16819 74520 -16808
rect 74982 -16813 75023 -16779
rect 75027 -16813 75034 -16771
rect 75127 -16779 75134 -16771
rect 75138 -16813 75179 -16779
rect 75483 -16795 75488 -16650
rect 75722 -16663 75763 -16629
rect 75767 -16663 75774 -16618
rect 75844 -16679 75849 -16363
rect 75867 -16379 75874 -16371
rect 75878 -16379 75883 -16363
rect 75878 -16413 75919 -16379
rect 75923 -16413 75930 -16371
rect 75867 -16462 75874 -16451
rect 75878 -16462 75883 -16413
rect 75878 -16496 75919 -16462
rect 75923 -16496 75930 -16451
rect 75867 -16546 75874 -16535
rect 75878 -16546 75883 -16496
rect 75878 -16580 75919 -16546
rect 75923 -16580 75930 -16535
rect 75867 -16629 75874 -16618
rect 75878 -16629 75883 -16580
rect 75878 -16663 75919 -16629
rect 75923 -16663 75930 -16618
rect 75867 -16697 75874 -16671
rect 75878 -16713 75883 -16663
rect 75787 -16777 75828 -16743
rect 74515 -16853 74520 -16819
rect 74524 -16853 74565 -16819
rect 74632 -16870 74673 -16836
rect 74677 -16870 74684 -16825
rect 74777 -16832 74784 -16821
rect 74788 -16866 74829 -16832
rect 75336 -16856 75377 -16822
rect 75381 -16856 75388 -16814
rect 75481 -16822 75488 -16814
rect 75492 -16856 75533 -16822
rect 75909 -16845 75916 -16697
rect 75932 -16713 75935 -16363
rect 75966 -16679 75969 -16363
rect 76023 -16379 76030 -16371
rect 75972 -16413 76013 -16379
rect 76034 -16413 76085 -16379
rect 76744 -16422 76749 -16406
rect 76767 -16422 76774 -16414
rect 76778 -16422 76783 -16406
rect 77074 -16408 77115 -16374
rect 77119 -16408 77126 -16363
rect 76023 -16462 76030 -16451
rect 76204 -16456 76245 -16422
rect 76276 -16456 76317 -16422
rect 76348 -16456 76389 -16422
rect 76492 -16456 76533 -16422
rect 76564 -16456 76677 -16422
rect 76708 -16456 76749 -16422
rect 76034 -16496 76075 -16462
rect 76023 -16546 76030 -16535
rect 76601 -16539 76642 -16505
rect 76034 -16580 76075 -16546
rect 76023 -16629 76030 -16618
rect 76034 -16663 76075 -16629
rect 76266 -16689 76307 -16655
rect 76311 -16689 76318 -16644
rect 76388 -16706 76393 -16588
rect 76411 -16655 76418 -16644
rect 76422 -16655 76427 -16622
rect 76458 -16655 76463 -16622
rect 76422 -16689 76463 -16655
rect 76467 -16689 76474 -16644
rect 76422 -16740 76427 -16689
rect 76458 -16740 76463 -16689
rect 76492 -16706 76497 -16589
rect 76601 -16623 76642 -16589
rect 76601 -16706 76642 -16672
rect 76744 -16706 76749 -16456
rect 76778 -16456 76819 -16422
rect 76767 -16505 76774 -16494
rect 76778 -16505 76783 -16456
rect 77074 -16491 77115 -16457
rect 77119 -16491 77126 -16446
rect 76778 -16539 76819 -16505
rect 76767 -16589 76774 -16578
rect 76778 -16589 76783 -16539
rect 76927 -16565 77036 -16499
rect 77196 -16507 77201 -16191
rect 77219 -16207 77226 -16199
rect 77230 -16207 77235 -16191
rect 77230 -16241 77271 -16207
rect 77275 -16241 77282 -16199
rect 77219 -16290 77226 -16279
rect 77230 -16290 77235 -16241
rect 77230 -16324 77271 -16290
rect 77275 -16324 77282 -16279
rect 77219 -16374 77226 -16363
rect 77230 -16374 77235 -16324
rect 77230 -16408 77271 -16374
rect 77275 -16408 77282 -16363
rect 77219 -16457 77226 -16446
rect 77230 -16457 77235 -16408
rect 77230 -16491 77271 -16457
rect 77275 -16491 77282 -16446
rect 77219 -16525 77226 -16499
rect 77230 -16541 77235 -16491
rect 76778 -16623 76819 -16589
rect 77139 -16605 77180 -16571
rect 76767 -16672 76774 -16661
rect 76778 -16672 76783 -16623
rect 76778 -16706 76819 -16672
rect 77261 -16673 77268 -16525
rect 77284 -16541 77287 -16191
rect 77318 -16507 77321 -16191
rect 77375 -16207 77382 -16199
rect 77324 -16241 77365 -16207
rect 77386 -16241 77437 -16207
rect 78301 -16231 78342 -16197
rect 78397 -16231 78438 -16197
rect 78493 -16231 78534 -16197
rect 80463 -16207 80470 -16199
rect 78094 -16250 78099 -16234
rect 78117 -16250 78124 -16242
rect 78128 -16250 78133 -16234
rect 77375 -16290 77382 -16279
rect 77554 -16284 77595 -16250
rect 77626 -16284 77667 -16250
rect 77698 -16284 77739 -16250
rect 77842 -16284 77883 -16250
rect 77914 -16284 78027 -16250
rect 78058 -16284 78099 -16250
rect 77386 -16324 77427 -16290
rect 77375 -16374 77382 -16363
rect 77951 -16367 77992 -16333
rect 77386 -16408 77427 -16374
rect 77375 -16457 77382 -16446
rect 77386 -16491 77427 -16457
rect 77616 -16517 77657 -16483
rect 77661 -16517 77668 -16472
rect 77738 -16534 77743 -16416
rect 77761 -16483 77768 -16472
rect 77772 -16483 77777 -16450
rect 77808 -16483 77813 -16450
rect 77772 -16517 77813 -16483
rect 77817 -16517 77824 -16472
rect 77772 -16568 77777 -16517
rect 77808 -16568 77813 -16517
rect 77842 -16534 77847 -16417
rect 77951 -16451 77992 -16417
rect 77951 -16534 77992 -16500
rect 78094 -16534 78099 -16284
rect 78128 -16284 78169 -16250
rect 78655 -16274 78696 -16240
rect 78751 -16274 78792 -16240
rect 78847 -16274 78888 -16240
rect 80354 -16241 80395 -16207
rect 80418 -16241 80470 -16207
rect 80498 -16241 80539 -16207
rect 78117 -16333 78124 -16322
rect 78128 -16333 78133 -16284
rect 78367 -16293 78374 -16285
rect 78467 -16293 78474 -16285
rect 78294 -16327 78363 -16293
rect 78366 -16327 78407 -16293
rect 78478 -16327 78519 -16293
rect 79009 -16317 79050 -16283
rect 79105 -16317 79146 -16283
rect 79201 -16317 79242 -16283
rect 79297 -16317 79338 -16283
rect 79393 -16317 79434 -16283
rect 80418 -16324 80459 -16290
rect 80463 -16324 80470 -16279
rect 78128 -16367 78169 -16333
rect 78721 -16336 78728 -16328
rect 78821 -16336 78828 -16328
rect 78117 -16417 78124 -16406
rect 78128 -16417 78133 -16367
rect 78322 -16410 78363 -16376
rect 78367 -16410 78374 -16365
rect 78467 -16376 78474 -16365
rect 78648 -16370 78717 -16336
rect 78720 -16370 78761 -16336
rect 78832 -16370 78873 -16336
rect 79557 -16360 79598 -16326
rect 79653 -16360 79694 -16326
rect 79749 -16360 79790 -16326
rect 79845 -16360 79886 -16326
rect 79941 -16360 79982 -16326
rect 80037 -16360 80078 -16326
rect 80133 -16360 80174 -16326
rect 78478 -16410 78519 -16376
rect 79111 -16379 79118 -16371
rect 78128 -16451 78169 -16417
rect 78117 -16500 78124 -16489
rect 78128 -16500 78133 -16451
rect 78322 -16494 78363 -16460
rect 78367 -16494 78374 -16449
rect 78467 -16460 78474 -16449
rect 78676 -16453 78717 -16419
rect 78721 -16453 78728 -16408
rect 78821 -16419 78828 -16408
rect 79002 -16413 79043 -16379
rect 79066 -16413 79118 -16379
rect 79146 -16413 79187 -16379
rect 78832 -16453 78873 -16419
rect 78478 -16494 78519 -16460
rect 78128 -16534 78169 -16500
rect 78128 -16568 78133 -16534
rect 76778 -16740 76783 -16706
rect 77074 -16723 77115 -16689
rect 77119 -16723 77126 -16681
rect 77261 -16741 77273 -16673
rect 77302 -16707 77307 -16639
rect 77347 -16671 77352 -16603
rect 77381 -16637 77386 -16571
rect 78322 -16577 78363 -16543
rect 78367 -16577 78374 -16532
rect 78467 -16543 78474 -16532
rect 78676 -16537 78717 -16503
rect 78721 -16537 78728 -16492
rect 78821 -16503 78828 -16492
rect 79066 -16496 79107 -16462
rect 79111 -16496 79118 -16451
rect 78832 -16537 78873 -16503
rect 78478 -16577 78519 -16543
rect 77391 -16621 77432 -16587
rect 77592 -16666 77633 -16632
rect 77361 -16689 77368 -16681
rect 77372 -16723 77413 -16689
rect 77592 -16734 77633 -16700
rect 74525 -16906 74566 -16872
rect 74597 -16906 74638 -16872
rect 74669 -16906 74710 -16872
rect 74982 -16913 75023 -16879
rect 75027 -16913 75034 -16868
rect 75127 -16879 75134 -16868
rect 75138 -16913 75179 -16879
rect 75722 -16895 75763 -16861
rect 75767 -16895 75774 -16853
rect 73616 -16959 74098 -16925
rect 74950 -16949 74991 -16915
rect 75022 -16949 75063 -16915
rect 75336 -16956 75377 -16922
rect 75381 -16956 75388 -16911
rect 75481 -16922 75488 -16911
rect 75909 -16913 75921 -16845
rect 75950 -16879 75955 -16811
rect 75995 -16843 76000 -16775
rect 76029 -16809 76034 -16743
rect 77261 -16753 77268 -16741
rect 77641 -16750 77646 -16616
rect 76039 -16793 76080 -16759
rect 76242 -16838 76283 -16804
rect 76009 -16861 76016 -16853
rect 76020 -16895 76061 -16861
rect 76242 -16906 76283 -16872
rect 75492 -16956 75533 -16922
rect 73616 -16985 74085 -16959
rect 73620 -16993 73827 -16985
rect 73636 -17003 73811 -16993
rect 73362 -17140 73543 -17114
rect 72869 -17174 72910 -17140
rect 72965 -17174 73006 -17140
rect 73061 -17174 73102 -17140
rect 73157 -17174 73198 -17140
rect 73253 -17174 73294 -17140
rect 73349 -17174 73543 -17140
rect 73362 -17200 73543 -17174
rect 73562 -17174 73669 -17050
rect 73821 -17062 73827 -17051
rect 73440 -17870 73481 -17200
rect 73562 -17228 73571 -17174
rect 73247 -17936 73398 -17924
rect 72915 -17970 73398 -17936
rect 73247 -17971 73398 -17970
rect 73428 -17971 73481 -17870
rect 73574 -17971 73615 -17174
rect 73620 -17971 73626 -17174
rect 73832 -17971 73873 -17062
rect 73966 -17971 74007 -16985
rect 74219 -17002 74260 -16968
rect 74315 -17002 74356 -16968
rect 74411 -17002 74452 -16968
rect 74507 -17002 74548 -16968
rect 74603 -17002 74644 -16968
rect 74699 -17002 74740 -16968
rect 74795 -17002 74836 -16968
rect 75304 -16992 75345 -16958
rect 75376 -16992 75417 -16958
rect 75722 -16995 75763 -16961
rect 75767 -16995 75774 -16950
rect 75909 -17001 75916 -16913
rect 76291 -16922 76296 -16788
rect 76009 -16961 76016 -16950
rect 76325 -16956 76330 -16762
rect 76365 -16778 76372 -16767
rect 76361 -16809 76372 -16778
rect 76687 -16796 76728 -16762
rect 76020 -16995 76061 -16961
rect 74957 -17045 74998 -17011
rect 75053 -17045 75094 -17011
rect 75149 -17045 75190 -17011
rect 75658 -17035 75699 -17001
rect 75730 -17035 75771 -17001
rect 75802 -17035 75843 -17001
rect 75874 -17029 75916 -17001
rect 76220 -17025 76261 -16991
rect 76265 -17025 76272 -16980
rect 76361 -16992 76366 -16809
rect 76395 -16995 76400 -16812
rect 75874 -17035 75915 -17029
rect 75311 -17088 75352 -17054
rect 75407 -17088 75448 -17054
rect 75503 -17088 75544 -17054
rect 76407 -17076 76414 -16809
rect 77036 -16819 77429 -16753
rect 77675 -16784 77680 -16590
rect 77715 -16606 77722 -16595
rect 77711 -16637 77722 -16606
rect 78037 -16624 78078 -16590
rect 76423 -16860 76464 -16826
rect 76772 -16830 76789 -16819
rect 76772 -16832 76778 -16830
rect 76423 -16928 76464 -16894
rect 76475 -16995 76480 -16860
rect 76706 -16874 76778 -16832
rect 76834 -16874 77429 -16819
rect 77570 -16853 77611 -16819
rect 77615 -16853 77622 -16808
rect 77711 -16820 77716 -16637
rect 77745 -16823 77750 -16640
rect 76706 -16877 77429 -16874
rect 76509 -16980 76514 -16892
rect 76626 -16942 76667 -16908
rect 76671 -16942 76678 -16900
rect 76507 -16991 76514 -16980
rect 76509 -17025 76514 -16991
rect 76518 -17025 76559 -16991
rect 76626 -17042 76667 -17008
rect 76671 -17042 76678 -16997
rect 76519 -17078 76560 -17044
rect 76591 -17078 76632 -17044
rect 76663 -17078 76704 -17044
rect 75665 -17131 75706 -17097
rect 75761 -17131 75802 -17097
rect 75857 -17131 75898 -17097
rect 75953 -17131 75994 -17097
rect 76049 -17131 76090 -17097
rect 76706 -17114 76857 -16877
rect 77036 -16899 77429 -16877
rect 76960 -16925 77429 -16899
rect 77757 -16904 77764 -16637
rect 77773 -16688 77814 -16654
rect 77773 -16756 77814 -16722
rect 77825 -16823 77830 -16688
rect 78387 -16691 78428 -16657
rect 78439 -16718 78444 -16641
rect 77859 -16808 77864 -16720
rect 77976 -16770 78017 -16736
rect 78021 -16770 78028 -16728
rect 78121 -16740 78128 -16729
rect 78132 -16774 78173 -16740
rect 78473 -16752 78478 -16607
rect 78676 -16620 78717 -16586
rect 78721 -16620 78728 -16575
rect 78821 -16586 78828 -16575
rect 79066 -16580 79107 -16546
rect 79111 -16580 79118 -16535
rect 78832 -16620 78873 -16586
rect 78741 -16734 78782 -16700
rect 78793 -16761 78798 -16684
rect 77857 -16819 77864 -16808
rect 78326 -16813 78367 -16779
rect 78371 -16813 78378 -16771
rect 78471 -16779 78478 -16771
rect 78482 -16813 78523 -16779
rect 78827 -16795 78832 -16650
rect 79066 -16663 79107 -16629
rect 79111 -16663 79118 -16618
rect 79188 -16679 79193 -16363
rect 79211 -16379 79218 -16371
rect 79222 -16379 79227 -16363
rect 79222 -16413 79263 -16379
rect 79267 -16413 79274 -16371
rect 79211 -16462 79218 -16451
rect 79222 -16462 79227 -16413
rect 79222 -16496 79263 -16462
rect 79267 -16496 79274 -16451
rect 79211 -16546 79218 -16535
rect 79222 -16546 79227 -16496
rect 79222 -16580 79263 -16546
rect 79267 -16580 79274 -16535
rect 79211 -16629 79218 -16618
rect 79222 -16629 79227 -16580
rect 79222 -16663 79263 -16629
rect 79267 -16663 79274 -16618
rect 79211 -16697 79218 -16671
rect 79222 -16713 79227 -16663
rect 79131 -16777 79172 -16743
rect 77859 -16853 77864 -16819
rect 77868 -16853 77909 -16819
rect 77976 -16870 78017 -16836
rect 78021 -16870 78028 -16825
rect 78121 -16832 78128 -16821
rect 78132 -16866 78173 -16832
rect 78680 -16856 78721 -16822
rect 78725 -16856 78732 -16814
rect 78825 -16822 78832 -16814
rect 78836 -16856 78877 -16822
rect 79253 -16845 79260 -16697
rect 79276 -16713 79279 -16363
rect 79310 -16679 79313 -16363
rect 79367 -16379 79374 -16371
rect 79316 -16413 79357 -16379
rect 79378 -16413 79429 -16379
rect 80088 -16422 80093 -16406
rect 80111 -16422 80118 -16414
rect 80122 -16422 80127 -16406
rect 80418 -16408 80459 -16374
rect 80463 -16408 80470 -16363
rect 79367 -16462 79374 -16451
rect 79548 -16456 79589 -16422
rect 79620 -16456 79661 -16422
rect 79692 -16456 79733 -16422
rect 79836 -16456 79877 -16422
rect 79908 -16456 80021 -16422
rect 80052 -16456 80093 -16422
rect 79378 -16496 79419 -16462
rect 79367 -16546 79374 -16535
rect 79945 -16539 79986 -16505
rect 79378 -16580 79419 -16546
rect 79367 -16629 79374 -16618
rect 79378 -16663 79419 -16629
rect 79610 -16689 79651 -16655
rect 79655 -16689 79662 -16644
rect 79732 -16706 79737 -16588
rect 79755 -16655 79762 -16644
rect 79766 -16655 79771 -16622
rect 79802 -16655 79807 -16622
rect 79766 -16689 79807 -16655
rect 79811 -16689 79818 -16644
rect 79766 -16740 79771 -16689
rect 79802 -16740 79807 -16689
rect 79836 -16706 79841 -16589
rect 79945 -16623 79986 -16589
rect 79945 -16706 79986 -16672
rect 80088 -16706 80093 -16456
rect 80122 -16456 80163 -16422
rect 80111 -16505 80118 -16494
rect 80122 -16505 80127 -16456
rect 80418 -16491 80459 -16457
rect 80463 -16491 80470 -16446
rect 80122 -16539 80163 -16505
rect 80111 -16589 80118 -16578
rect 80122 -16589 80127 -16539
rect 80271 -16565 80380 -16499
rect 80540 -16507 80545 -16191
rect 80563 -16207 80570 -16199
rect 80574 -16207 80579 -16191
rect 80574 -16241 80615 -16207
rect 80619 -16241 80626 -16199
rect 80563 -16290 80570 -16279
rect 80574 -16290 80579 -16241
rect 80574 -16324 80615 -16290
rect 80619 -16324 80626 -16279
rect 80563 -16374 80570 -16363
rect 80574 -16374 80579 -16324
rect 80574 -16408 80615 -16374
rect 80619 -16408 80626 -16363
rect 80563 -16457 80570 -16446
rect 80574 -16457 80579 -16408
rect 80574 -16491 80615 -16457
rect 80619 -16491 80626 -16446
rect 80563 -16525 80570 -16499
rect 80574 -16541 80579 -16491
rect 80122 -16623 80163 -16589
rect 80483 -16605 80524 -16571
rect 80111 -16672 80118 -16661
rect 80122 -16672 80127 -16623
rect 80122 -16706 80163 -16672
rect 80605 -16673 80612 -16525
rect 80628 -16541 80631 -16191
rect 80662 -16507 80665 -16191
rect 80719 -16207 80726 -16199
rect 80668 -16241 80709 -16207
rect 80730 -16241 80781 -16207
rect 81645 -16231 81686 -16197
rect 81741 -16231 81782 -16197
rect 81837 -16231 81878 -16197
rect 83807 -16207 83814 -16199
rect 81438 -16250 81443 -16234
rect 81461 -16250 81468 -16242
rect 81472 -16250 81477 -16234
rect 80719 -16290 80726 -16279
rect 80898 -16284 80939 -16250
rect 80970 -16284 81011 -16250
rect 81042 -16284 81083 -16250
rect 81186 -16284 81227 -16250
rect 81258 -16284 81371 -16250
rect 81402 -16284 81443 -16250
rect 80730 -16324 80771 -16290
rect 80719 -16374 80726 -16363
rect 81295 -16367 81336 -16333
rect 80730 -16408 80771 -16374
rect 80719 -16457 80726 -16446
rect 80730 -16491 80771 -16457
rect 80960 -16517 81001 -16483
rect 81005 -16517 81012 -16472
rect 81082 -16534 81087 -16416
rect 81105 -16483 81112 -16472
rect 81116 -16483 81121 -16450
rect 81152 -16483 81157 -16450
rect 81116 -16517 81157 -16483
rect 81161 -16517 81168 -16472
rect 81116 -16568 81121 -16517
rect 81152 -16568 81157 -16517
rect 81186 -16534 81191 -16417
rect 81295 -16451 81336 -16417
rect 81295 -16534 81336 -16500
rect 81438 -16534 81443 -16284
rect 81472 -16284 81513 -16250
rect 81999 -16274 82040 -16240
rect 82095 -16274 82136 -16240
rect 82191 -16274 82232 -16240
rect 83698 -16241 83739 -16207
rect 83762 -16241 83814 -16207
rect 83842 -16241 83883 -16207
rect 81461 -16333 81468 -16322
rect 81472 -16333 81477 -16284
rect 81711 -16293 81718 -16285
rect 81811 -16293 81818 -16285
rect 81638 -16327 81707 -16293
rect 81710 -16327 81751 -16293
rect 81822 -16327 81863 -16293
rect 82353 -16317 82394 -16283
rect 82449 -16317 82490 -16283
rect 82545 -16317 82586 -16283
rect 82641 -16317 82682 -16283
rect 82737 -16317 82778 -16283
rect 83762 -16324 83803 -16290
rect 83807 -16324 83814 -16279
rect 81472 -16367 81513 -16333
rect 82065 -16336 82072 -16328
rect 82165 -16336 82172 -16328
rect 81461 -16417 81468 -16406
rect 81472 -16417 81477 -16367
rect 81666 -16410 81707 -16376
rect 81711 -16410 81718 -16365
rect 81811 -16376 81818 -16365
rect 81992 -16370 82061 -16336
rect 82064 -16370 82105 -16336
rect 82176 -16370 82217 -16336
rect 82901 -16360 82942 -16326
rect 82997 -16360 83038 -16326
rect 83093 -16360 83134 -16326
rect 83189 -16360 83230 -16326
rect 83285 -16360 83326 -16326
rect 83381 -16360 83422 -16326
rect 83477 -16360 83518 -16326
rect 81822 -16410 81863 -16376
rect 82455 -16379 82462 -16371
rect 81472 -16451 81513 -16417
rect 81461 -16500 81468 -16489
rect 81472 -16500 81477 -16451
rect 81666 -16494 81707 -16460
rect 81711 -16494 81718 -16449
rect 81811 -16460 81818 -16449
rect 82020 -16453 82061 -16419
rect 82065 -16453 82072 -16408
rect 82165 -16419 82172 -16408
rect 82346 -16413 82387 -16379
rect 82410 -16413 82462 -16379
rect 82490 -16413 82531 -16379
rect 82176 -16453 82217 -16419
rect 81822 -16494 81863 -16460
rect 81472 -16534 81513 -16500
rect 81472 -16568 81477 -16534
rect 80122 -16740 80127 -16706
rect 80418 -16723 80459 -16689
rect 80463 -16723 80470 -16681
rect 80605 -16741 80617 -16673
rect 80646 -16707 80651 -16639
rect 80691 -16671 80696 -16603
rect 80725 -16637 80730 -16571
rect 81666 -16577 81707 -16543
rect 81711 -16577 81718 -16532
rect 81811 -16543 81818 -16532
rect 82020 -16537 82061 -16503
rect 82065 -16537 82072 -16492
rect 82165 -16503 82172 -16492
rect 82410 -16496 82451 -16462
rect 82455 -16496 82462 -16451
rect 82176 -16537 82217 -16503
rect 81822 -16577 81863 -16543
rect 80735 -16621 80776 -16587
rect 80936 -16666 80977 -16632
rect 80705 -16689 80712 -16681
rect 80716 -16723 80757 -16689
rect 80936 -16734 80977 -16700
rect 77869 -16906 77910 -16872
rect 77941 -16906 77982 -16872
rect 78013 -16906 78054 -16872
rect 78326 -16913 78367 -16879
rect 78371 -16913 78378 -16868
rect 78471 -16879 78478 -16868
rect 78482 -16913 78523 -16879
rect 79066 -16895 79107 -16861
rect 79111 -16895 79118 -16853
rect 76960 -16959 77442 -16925
rect 78294 -16949 78335 -16915
rect 78366 -16949 78407 -16915
rect 78680 -16956 78721 -16922
rect 78725 -16956 78732 -16911
rect 78825 -16922 78832 -16911
rect 79253 -16913 79265 -16845
rect 79294 -16879 79299 -16811
rect 79339 -16843 79344 -16775
rect 79373 -16809 79378 -16743
rect 80605 -16753 80612 -16741
rect 80985 -16750 80990 -16616
rect 79383 -16793 79424 -16759
rect 79586 -16838 79627 -16804
rect 79353 -16861 79360 -16853
rect 79364 -16895 79405 -16861
rect 79586 -16906 79627 -16872
rect 78836 -16956 78877 -16922
rect 76960 -16985 77429 -16959
rect 76964 -16993 77171 -16985
rect 76980 -17003 77155 -16993
rect 76706 -17140 76887 -17114
rect 76213 -17174 76254 -17140
rect 76309 -17174 76350 -17140
rect 76405 -17174 76446 -17140
rect 76501 -17174 76542 -17140
rect 76597 -17174 76638 -17140
rect 76693 -17174 76887 -17140
rect 76706 -17200 76887 -17174
rect 76906 -17174 77013 -17050
rect 77165 -17062 77171 -17051
rect 76784 -17870 76825 -17200
rect 76906 -17228 76915 -17174
rect 76591 -17936 76742 -17924
rect 76259 -17970 76742 -17936
rect 76591 -17971 76742 -17970
rect 76772 -17971 76825 -17870
rect 76918 -17971 76959 -17174
rect 76964 -17971 76970 -17174
rect 77176 -17971 77217 -17062
rect 77310 -17971 77351 -16985
rect 77563 -17002 77604 -16968
rect 77659 -17002 77700 -16968
rect 77755 -17002 77796 -16968
rect 77851 -17002 77892 -16968
rect 77947 -17002 77988 -16968
rect 78043 -17002 78084 -16968
rect 78139 -17002 78180 -16968
rect 78648 -16992 78689 -16958
rect 78720 -16992 78761 -16958
rect 79066 -16995 79107 -16961
rect 79111 -16995 79118 -16950
rect 79253 -17001 79260 -16913
rect 79635 -16922 79640 -16788
rect 79353 -16961 79360 -16950
rect 79669 -16956 79674 -16762
rect 79709 -16778 79716 -16767
rect 79705 -16809 79716 -16778
rect 80031 -16796 80072 -16762
rect 79364 -16995 79405 -16961
rect 78301 -17045 78342 -17011
rect 78397 -17045 78438 -17011
rect 78493 -17045 78534 -17011
rect 79002 -17035 79043 -17001
rect 79074 -17035 79115 -17001
rect 79146 -17035 79187 -17001
rect 79218 -17029 79260 -17001
rect 79564 -17025 79605 -16991
rect 79609 -17025 79616 -16980
rect 79705 -16992 79710 -16809
rect 79739 -16995 79744 -16812
rect 79218 -17035 79259 -17029
rect 78655 -17088 78696 -17054
rect 78751 -17088 78792 -17054
rect 78847 -17088 78888 -17054
rect 79751 -17076 79758 -16809
rect 80380 -16819 80773 -16753
rect 81019 -16784 81024 -16590
rect 81059 -16606 81066 -16595
rect 81055 -16637 81066 -16606
rect 81381 -16624 81422 -16590
rect 79767 -16860 79808 -16826
rect 80116 -16830 80133 -16819
rect 80116 -16832 80122 -16830
rect 79767 -16928 79808 -16894
rect 79819 -16995 79824 -16860
rect 80050 -16874 80122 -16832
rect 80178 -16874 80773 -16819
rect 80914 -16853 80955 -16819
rect 80959 -16853 80966 -16808
rect 81055 -16820 81060 -16637
rect 81089 -16823 81094 -16640
rect 80050 -16877 80773 -16874
rect 79853 -16980 79858 -16892
rect 79970 -16942 80011 -16908
rect 80015 -16942 80022 -16900
rect 79851 -16991 79858 -16980
rect 79853 -17025 79858 -16991
rect 79862 -17025 79903 -16991
rect 79970 -17042 80011 -17008
rect 80015 -17042 80022 -16997
rect 79863 -17078 79904 -17044
rect 79935 -17078 79976 -17044
rect 80007 -17078 80048 -17044
rect 79009 -17131 79050 -17097
rect 79105 -17131 79146 -17097
rect 79201 -17131 79242 -17097
rect 79297 -17131 79338 -17097
rect 79393 -17131 79434 -17097
rect 80050 -17114 80201 -16877
rect 80380 -16899 80773 -16877
rect 80304 -16925 80773 -16899
rect 81101 -16904 81108 -16637
rect 81117 -16688 81158 -16654
rect 81117 -16756 81158 -16722
rect 81169 -16823 81174 -16688
rect 81731 -16691 81772 -16657
rect 81783 -16718 81788 -16641
rect 81203 -16808 81208 -16720
rect 81320 -16770 81361 -16736
rect 81365 -16770 81372 -16728
rect 81465 -16740 81472 -16729
rect 81476 -16774 81517 -16740
rect 81817 -16752 81822 -16607
rect 82020 -16620 82061 -16586
rect 82065 -16620 82072 -16575
rect 82165 -16586 82172 -16575
rect 82410 -16580 82451 -16546
rect 82455 -16580 82462 -16535
rect 82176 -16620 82217 -16586
rect 82085 -16734 82126 -16700
rect 82137 -16761 82142 -16684
rect 81201 -16819 81208 -16808
rect 81670 -16813 81711 -16779
rect 81715 -16813 81722 -16771
rect 81815 -16779 81822 -16771
rect 81826 -16813 81867 -16779
rect 82171 -16795 82176 -16650
rect 82410 -16663 82451 -16629
rect 82455 -16663 82462 -16618
rect 82532 -16679 82537 -16363
rect 82555 -16379 82562 -16371
rect 82566 -16379 82571 -16363
rect 82566 -16413 82607 -16379
rect 82611 -16413 82618 -16371
rect 82555 -16462 82562 -16451
rect 82566 -16462 82571 -16413
rect 82566 -16496 82607 -16462
rect 82611 -16496 82618 -16451
rect 82555 -16546 82562 -16535
rect 82566 -16546 82571 -16496
rect 82566 -16580 82607 -16546
rect 82611 -16580 82618 -16535
rect 82555 -16629 82562 -16618
rect 82566 -16629 82571 -16580
rect 82566 -16663 82607 -16629
rect 82611 -16663 82618 -16618
rect 82555 -16697 82562 -16671
rect 82566 -16713 82571 -16663
rect 82475 -16777 82516 -16743
rect 81203 -16853 81208 -16819
rect 81212 -16853 81253 -16819
rect 81320 -16870 81361 -16836
rect 81365 -16870 81372 -16825
rect 81465 -16832 81472 -16821
rect 81476 -16866 81517 -16832
rect 82024 -16856 82065 -16822
rect 82069 -16856 82076 -16814
rect 82169 -16822 82176 -16814
rect 82180 -16856 82221 -16822
rect 82597 -16845 82604 -16697
rect 82620 -16713 82623 -16363
rect 82654 -16679 82657 -16363
rect 82711 -16379 82718 -16371
rect 82660 -16413 82701 -16379
rect 82722 -16413 82773 -16379
rect 83432 -16422 83437 -16406
rect 83455 -16422 83462 -16414
rect 83466 -16422 83471 -16406
rect 83762 -16408 83803 -16374
rect 83807 -16408 83814 -16363
rect 82711 -16462 82718 -16451
rect 82892 -16456 82933 -16422
rect 82964 -16456 83005 -16422
rect 83036 -16456 83077 -16422
rect 83180 -16456 83221 -16422
rect 83252 -16456 83365 -16422
rect 83396 -16456 83437 -16422
rect 82722 -16496 82763 -16462
rect 82711 -16546 82718 -16535
rect 83289 -16539 83330 -16505
rect 82722 -16580 82763 -16546
rect 82711 -16629 82718 -16618
rect 82722 -16663 82763 -16629
rect 82954 -16689 82995 -16655
rect 82999 -16689 83006 -16644
rect 83076 -16706 83081 -16588
rect 83099 -16655 83106 -16644
rect 83110 -16655 83115 -16622
rect 83146 -16655 83151 -16622
rect 83110 -16689 83151 -16655
rect 83155 -16689 83162 -16644
rect 83110 -16740 83115 -16689
rect 83146 -16740 83151 -16689
rect 83180 -16706 83185 -16589
rect 83289 -16623 83330 -16589
rect 83289 -16706 83330 -16672
rect 83432 -16706 83437 -16456
rect 83466 -16456 83507 -16422
rect 83455 -16505 83462 -16494
rect 83466 -16505 83471 -16456
rect 83762 -16491 83803 -16457
rect 83807 -16491 83814 -16446
rect 83466 -16539 83507 -16505
rect 83455 -16589 83462 -16578
rect 83466 -16589 83471 -16539
rect 83615 -16565 83724 -16499
rect 83884 -16507 83889 -16191
rect 83907 -16207 83914 -16199
rect 83918 -16207 83923 -16191
rect 83918 -16241 83959 -16207
rect 83963 -16241 83970 -16199
rect 83907 -16290 83914 -16279
rect 83918 -16290 83923 -16241
rect 83918 -16324 83959 -16290
rect 83963 -16324 83970 -16279
rect 83907 -16374 83914 -16363
rect 83918 -16374 83923 -16324
rect 83918 -16408 83959 -16374
rect 83963 -16408 83970 -16363
rect 83907 -16457 83914 -16446
rect 83918 -16457 83923 -16408
rect 83918 -16491 83959 -16457
rect 83963 -16491 83970 -16446
rect 83907 -16525 83914 -16499
rect 83918 -16541 83923 -16491
rect 83466 -16623 83507 -16589
rect 83827 -16605 83868 -16571
rect 83455 -16672 83462 -16661
rect 83466 -16672 83471 -16623
rect 83466 -16706 83507 -16672
rect 83949 -16673 83956 -16525
rect 83972 -16541 83975 -16191
rect 84006 -16507 84009 -16191
rect 84063 -16207 84070 -16199
rect 84012 -16241 84053 -16207
rect 84074 -16241 84125 -16207
rect 84989 -16231 85030 -16197
rect 85085 -16231 85126 -16197
rect 85181 -16231 85222 -16197
rect 87151 -16207 87158 -16199
rect 84782 -16250 84787 -16234
rect 84805 -16250 84812 -16242
rect 84816 -16250 84821 -16234
rect 84063 -16290 84070 -16279
rect 84242 -16284 84283 -16250
rect 84314 -16284 84355 -16250
rect 84386 -16284 84427 -16250
rect 84530 -16284 84571 -16250
rect 84602 -16284 84715 -16250
rect 84746 -16284 84787 -16250
rect 84074 -16324 84115 -16290
rect 84063 -16374 84070 -16363
rect 84639 -16367 84680 -16333
rect 84074 -16408 84115 -16374
rect 84063 -16457 84070 -16446
rect 84074 -16491 84115 -16457
rect 84304 -16517 84345 -16483
rect 84349 -16517 84356 -16472
rect 84426 -16534 84431 -16416
rect 84449 -16483 84456 -16472
rect 84460 -16483 84465 -16450
rect 84496 -16483 84501 -16450
rect 84460 -16517 84501 -16483
rect 84505 -16517 84512 -16472
rect 84460 -16568 84465 -16517
rect 84496 -16568 84501 -16517
rect 84530 -16534 84535 -16417
rect 84639 -16451 84680 -16417
rect 84639 -16534 84680 -16500
rect 84782 -16534 84787 -16284
rect 84816 -16284 84857 -16250
rect 85343 -16274 85384 -16240
rect 85439 -16274 85480 -16240
rect 85535 -16274 85576 -16240
rect 87042 -16241 87083 -16207
rect 87106 -16241 87158 -16207
rect 87186 -16241 87227 -16207
rect 84805 -16333 84812 -16322
rect 84816 -16333 84821 -16284
rect 85055 -16293 85062 -16285
rect 85155 -16293 85162 -16285
rect 84982 -16327 85051 -16293
rect 85054 -16327 85095 -16293
rect 85166 -16327 85207 -16293
rect 85697 -16317 85738 -16283
rect 85793 -16317 85834 -16283
rect 85889 -16317 85930 -16283
rect 85985 -16317 86026 -16283
rect 86081 -16317 86122 -16283
rect 87106 -16324 87147 -16290
rect 87151 -16324 87158 -16279
rect 84816 -16367 84857 -16333
rect 85409 -16336 85416 -16328
rect 85509 -16336 85516 -16328
rect 84805 -16417 84812 -16406
rect 84816 -16417 84821 -16367
rect 85010 -16410 85051 -16376
rect 85055 -16410 85062 -16365
rect 85155 -16376 85162 -16365
rect 85336 -16370 85405 -16336
rect 85408 -16370 85449 -16336
rect 85520 -16370 85561 -16336
rect 86245 -16360 86286 -16326
rect 86341 -16360 86382 -16326
rect 86437 -16360 86478 -16326
rect 86533 -16360 86574 -16326
rect 86629 -16360 86670 -16326
rect 86725 -16360 86766 -16326
rect 86821 -16360 86862 -16326
rect 85166 -16410 85207 -16376
rect 85799 -16379 85806 -16371
rect 84816 -16451 84857 -16417
rect 84805 -16500 84812 -16489
rect 84816 -16500 84821 -16451
rect 85010 -16494 85051 -16460
rect 85055 -16494 85062 -16449
rect 85155 -16460 85162 -16449
rect 85364 -16453 85405 -16419
rect 85409 -16453 85416 -16408
rect 85509 -16419 85516 -16408
rect 85690 -16413 85731 -16379
rect 85754 -16413 85806 -16379
rect 85834 -16413 85875 -16379
rect 85520 -16453 85561 -16419
rect 85166 -16494 85207 -16460
rect 84816 -16534 84857 -16500
rect 84816 -16568 84821 -16534
rect 83466 -16740 83471 -16706
rect 83762 -16723 83803 -16689
rect 83807 -16723 83814 -16681
rect 83949 -16741 83961 -16673
rect 83990 -16707 83995 -16639
rect 84035 -16671 84040 -16603
rect 84069 -16637 84074 -16571
rect 85010 -16577 85051 -16543
rect 85055 -16577 85062 -16532
rect 85155 -16543 85162 -16532
rect 85364 -16537 85405 -16503
rect 85409 -16537 85416 -16492
rect 85509 -16503 85516 -16492
rect 85754 -16496 85795 -16462
rect 85799 -16496 85806 -16451
rect 85520 -16537 85561 -16503
rect 85166 -16577 85207 -16543
rect 84079 -16621 84120 -16587
rect 84280 -16666 84321 -16632
rect 84049 -16689 84056 -16681
rect 84060 -16723 84101 -16689
rect 84280 -16734 84321 -16700
rect 81213 -16906 81254 -16872
rect 81285 -16906 81326 -16872
rect 81357 -16906 81398 -16872
rect 81670 -16913 81711 -16879
rect 81715 -16913 81722 -16868
rect 81815 -16879 81822 -16868
rect 81826 -16913 81867 -16879
rect 82410 -16895 82451 -16861
rect 82455 -16895 82462 -16853
rect 80304 -16959 80786 -16925
rect 81638 -16949 81679 -16915
rect 81710 -16949 81751 -16915
rect 82024 -16956 82065 -16922
rect 82069 -16956 82076 -16911
rect 82169 -16922 82176 -16911
rect 82597 -16913 82609 -16845
rect 82638 -16879 82643 -16811
rect 82683 -16843 82688 -16775
rect 82717 -16809 82722 -16743
rect 83949 -16753 83956 -16741
rect 84329 -16750 84334 -16616
rect 82727 -16793 82768 -16759
rect 82930 -16838 82971 -16804
rect 82697 -16861 82704 -16853
rect 82708 -16895 82749 -16861
rect 82930 -16906 82971 -16872
rect 82180 -16956 82221 -16922
rect 80304 -16985 80773 -16959
rect 80308 -16993 80515 -16985
rect 80324 -17003 80499 -16993
rect 80050 -17140 80231 -17114
rect 79557 -17174 79598 -17140
rect 79653 -17174 79694 -17140
rect 79749 -17174 79790 -17140
rect 79845 -17174 79886 -17140
rect 79941 -17174 79982 -17140
rect 80037 -17174 80231 -17140
rect 80050 -17200 80231 -17174
rect 80250 -17174 80357 -17050
rect 80509 -17062 80515 -17051
rect 80128 -17870 80169 -17200
rect 80250 -17228 80259 -17174
rect 79935 -17936 80086 -17924
rect 79603 -17970 80086 -17936
rect 79935 -17971 80086 -17970
rect 80116 -17971 80169 -17870
rect 80262 -17971 80303 -17174
rect 80308 -17971 80314 -17174
rect 80520 -17971 80561 -17062
rect 80654 -17971 80695 -16985
rect 80907 -17002 80948 -16968
rect 81003 -17002 81044 -16968
rect 81099 -17002 81140 -16968
rect 81195 -17002 81236 -16968
rect 81291 -17002 81332 -16968
rect 81387 -17002 81428 -16968
rect 81483 -17002 81524 -16968
rect 81992 -16992 82033 -16958
rect 82064 -16992 82105 -16958
rect 82410 -16995 82451 -16961
rect 82455 -16995 82462 -16950
rect 82597 -17001 82604 -16913
rect 82979 -16922 82984 -16788
rect 82697 -16961 82704 -16950
rect 83013 -16956 83018 -16762
rect 83053 -16778 83060 -16767
rect 83049 -16809 83060 -16778
rect 83375 -16796 83416 -16762
rect 82708 -16995 82749 -16961
rect 81645 -17045 81686 -17011
rect 81741 -17045 81782 -17011
rect 81837 -17045 81878 -17011
rect 82346 -17035 82387 -17001
rect 82418 -17035 82459 -17001
rect 82490 -17035 82531 -17001
rect 82562 -17029 82604 -17001
rect 82908 -17025 82949 -16991
rect 82953 -17025 82960 -16980
rect 83049 -16992 83054 -16809
rect 83083 -16995 83088 -16812
rect 82562 -17035 82603 -17029
rect 81999 -17088 82040 -17054
rect 82095 -17088 82136 -17054
rect 82191 -17088 82232 -17054
rect 83095 -17076 83102 -16809
rect 83724 -16819 84117 -16753
rect 84363 -16784 84368 -16590
rect 84403 -16606 84410 -16595
rect 84399 -16637 84410 -16606
rect 84725 -16624 84766 -16590
rect 83111 -16860 83152 -16826
rect 83460 -16830 83477 -16819
rect 83460 -16832 83466 -16830
rect 83111 -16928 83152 -16894
rect 83163 -16995 83168 -16860
rect 83394 -16874 83466 -16832
rect 83522 -16874 84117 -16819
rect 84258 -16853 84299 -16819
rect 84303 -16853 84310 -16808
rect 84399 -16820 84404 -16637
rect 84433 -16823 84438 -16640
rect 83394 -16877 84117 -16874
rect 83197 -16980 83202 -16892
rect 83314 -16942 83355 -16908
rect 83359 -16942 83366 -16900
rect 83195 -16991 83202 -16980
rect 83197 -17025 83202 -16991
rect 83206 -17025 83247 -16991
rect 83314 -17042 83355 -17008
rect 83359 -17042 83366 -16997
rect 83207 -17078 83248 -17044
rect 83279 -17078 83320 -17044
rect 83351 -17078 83392 -17044
rect 82353 -17131 82394 -17097
rect 82449 -17131 82490 -17097
rect 82545 -17131 82586 -17097
rect 82641 -17131 82682 -17097
rect 82737 -17131 82778 -17097
rect 83394 -17114 83545 -16877
rect 83724 -16899 84117 -16877
rect 83648 -16925 84117 -16899
rect 84445 -16904 84452 -16637
rect 84461 -16688 84502 -16654
rect 84461 -16756 84502 -16722
rect 84513 -16823 84518 -16688
rect 85075 -16691 85116 -16657
rect 85127 -16718 85132 -16641
rect 84547 -16808 84552 -16720
rect 84664 -16770 84705 -16736
rect 84709 -16770 84716 -16728
rect 84809 -16740 84816 -16729
rect 84820 -16774 84861 -16740
rect 85161 -16752 85166 -16607
rect 85364 -16620 85405 -16586
rect 85409 -16620 85416 -16575
rect 85509 -16586 85516 -16575
rect 85754 -16580 85795 -16546
rect 85799 -16580 85806 -16535
rect 85520 -16620 85561 -16586
rect 85429 -16734 85470 -16700
rect 85481 -16761 85486 -16684
rect 84545 -16819 84552 -16808
rect 85014 -16813 85055 -16779
rect 85059 -16813 85066 -16771
rect 85159 -16779 85166 -16771
rect 85170 -16813 85211 -16779
rect 85515 -16795 85520 -16650
rect 85754 -16663 85795 -16629
rect 85799 -16663 85806 -16618
rect 85876 -16679 85881 -16363
rect 85899 -16379 85906 -16371
rect 85910 -16379 85915 -16363
rect 85910 -16413 85951 -16379
rect 85955 -16413 85962 -16371
rect 85899 -16462 85906 -16451
rect 85910 -16462 85915 -16413
rect 85910 -16496 85951 -16462
rect 85955 -16496 85962 -16451
rect 85899 -16546 85906 -16535
rect 85910 -16546 85915 -16496
rect 85910 -16580 85951 -16546
rect 85955 -16580 85962 -16535
rect 85899 -16629 85906 -16618
rect 85910 -16629 85915 -16580
rect 85910 -16663 85951 -16629
rect 85955 -16663 85962 -16618
rect 85899 -16697 85906 -16671
rect 85910 -16713 85915 -16663
rect 85819 -16777 85860 -16743
rect 84547 -16853 84552 -16819
rect 84556 -16853 84597 -16819
rect 84664 -16870 84705 -16836
rect 84709 -16870 84716 -16825
rect 84809 -16832 84816 -16821
rect 84820 -16866 84861 -16832
rect 85368 -16856 85409 -16822
rect 85413 -16856 85420 -16814
rect 85513 -16822 85520 -16814
rect 85524 -16856 85565 -16822
rect 85941 -16845 85948 -16697
rect 85964 -16713 85967 -16363
rect 85998 -16679 86001 -16363
rect 86055 -16379 86062 -16371
rect 86004 -16413 86045 -16379
rect 86066 -16413 86117 -16379
rect 86776 -16422 86781 -16406
rect 86799 -16422 86806 -16414
rect 86810 -16422 86815 -16406
rect 87106 -16408 87147 -16374
rect 87151 -16408 87158 -16363
rect 86055 -16462 86062 -16451
rect 86236 -16456 86277 -16422
rect 86308 -16456 86349 -16422
rect 86380 -16456 86421 -16422
rect 86524 -16456 86565 -16422
rect 86596 -16456 86709 -16422
rect 86740 -16456 86781 -16422
rect 86066 -16496 86107 -16462
rect 86055 -16546 86062 -16535
rect 86633 -16539 86674 -16505
rect 86066 -16580 86107 -16546
rect 86055 -16629 86062 -16618
rect 86066 -16663 86107 -16629
rect 86298 -16689 86339 -16655
rect 86343 -16689 86350 -16644
rect 86420 -16706 86425 -16588
rect 86443 -16655 86450 -16644
rect 86454 -16655 86459 -16622
rect 86490 -16655 86495 -16622
rect 86454 -16689 86495 -16655
rect 86499 -16689 86506 -16644
rect 86454 -16740 86459 -16689
rect 86490 -16740 86495 -16689
rect 86524 -16706 86529 -16589
rect 86633 -16623 86674 -16589
rect 86633 -16706 86674 -16672
rect 86776 -16706 86781 -16456
rect 86810 -16456 86851 -16422
rect 86799 -16505 86806 -16494
rect 86810 -16505 86815 -16456
rect 87106 -16491 87147 -16457
rect 87151 -16491 87158 -16446
rect 86810 -16539 86851 -16505
rect 86799 -16589 86806 -16578
rect 86810 -16589 86815 -16539
rect 86959 -16565 87068 -16499
rect 87228 -16507 87233 -16191
rect 87251 -16207 87258 -16199
rect 87262 -16207 87267 -16191
rect 87262 -16241 87303 -16207
rect 87307 -16241 87314 -16199
rect 87251 -16290 87258 -16279
rect 87262 -16290 87267 -16241
rect 87262 -16324 87303 -16290
rect 87307 -16324 87314 -16279
rect 87251 -16374 87258 -16363
rect 87262 -16374 87267 -16324
rect 87262 -16408 87303 -16374
rect 87307 -16408 87314 -16363
rect 87251 -16457 87258 -16446
rect 87262 -16457 87267 -16408
rect 87262 -16491 87303 -16457
rect 87307 -16491 87314 -16446
rect 87251 -16525 87258 -16499
rect 87262 -16541 87267 -16491
rect 86810 -16623 86851 -16589
rect 87171 -16605 87212 -16571
rect 86799 -16672 86806 -16661
rect 86810 -16672 86815 -16623
rect 86810 -16706 86851 -16672
rect 87293 -16673 87300 -16525
rect 87316 -16541 87319 -16191
rect 87350 -16507 87353 -16191
rect 87407 -16207 87414 -16199
rect 87356 -16241 87397 -16207
rect 87418 -16241 87469 -16207
rect 88333 -16231 88374 -16197
rect 88429 -16231 88470 -16197
rect 88525 -16231 88566 -16197
rect 90495 -16207 90502 -16199
rect 88126 -16250 88131 -16234
rect 88149 -16250 88156 -16242
rect 88160 -16250 88165 -16234
rect 87407 -16290 87414 -16279
rect 87586 -16284 87627 -16250
rect 87658 -16284 87699 -16250
rect 87730 -16284 87771 -16250
rect 87874 -16284 87915 -16250
rect 87946 -16284 88059 -16250
rect 88090 -16284 88131 -16250
rect 87418 -16324 87459 -16290
rect 87407 -16374 87414 -16363
rect 87983 -16367 88024 -16333
rect 87418 -16408 87459 -16374
rect 87407 -16457 87414 -16446
rect 87418 -16491 87459 -16457
rect 87648 -16517 87689 -16483
rect 87693 -16517 87700 -16472
rect 87770 -16534 87775 -16416
rect 87793 -16483 87800 -16472
rect 87804 -16483 87809 -16450
rect 87840 -16483 87845 -16450
rect 87804 -16517 87845 -16483
rect 87849 -16517 87856 -16472
rect 87804 -16568 87809 -16517
rect 87840 -16568 87845 -16517
rect 87874 -16534 87879 -16417
rect 87983 -16451 88024 -16417
rect 87983 -16534 88024 -16500
rect 88126 -16534 88131 -16284
rect 88160 -16284 88201 -16250
rect 88687 -16274 88728 -16240
rect 88783 -16274 88824 -16240
rect 88879 -16274 88920 -16240
rect 90386 -16241 90427 -16207
rect 90450 -16241 90502 -16207
rect 90530 -16241 90571 -16207
rect 88149 -16333 88156 -16322
rect 88160 -16333 88165 -16284
rect 88399 -16293 88406 -16285
rect 88499 -16293 88506 -16285
rect 88326 -16327 88395 -16293
rect 88398 -16327 88439 -16293
rect 88510 -16327 88551 -16293
rect 89041 -16317 89082 -16283
rect 89137 -16317 89178 -16283
rect 89233 -16317 89274 -16283
rect 89329 -16317 89370 -16283
rect 89425 -16317 89466 -16283
rect 90450 -16324 90491 -16290
rect 90495 -16324 90502 -16279
rect 88160 -16367 88201 -16333
rect 88753 -16336 88760 -16328
rect 88853 -16336 88860 -16328
rect 88149 -16417 88156 -16406
rect 88160 -16417 88165 -16367
rect 88354 -16410 88395 -16376
rect 88399 -16410 88406 -16365
rect 88499 -16376 88506 -16365
rect 88680 -16370 88749 -16336
rect 88752 -16370 88793 -16336
rect 88864 -16370 88905 -16336
rect 89589 -16360 89630 -16326
rect 89685 -16360 89726 -16326
rect 89781 -16360 89822 -16326
rect 89877 -16360 89918 -16326
rect 89973 -16360 90014 -16326
rect 90069 -16360 90110 -16326
rect 90165 -16360 90206 -16326
rect 88510 -16410 88551 -16376
rect 89143 -16379 89150 -16371
rect 88160 -16451 88201 -16417
rect 88149 -16500 88156 -16489
rect 88160 -16500 88165 -16451
rect 88354 -16494 88395 -16460
rect 88399 -16494 88406 -16449
rect 88499 -16460 88506 -16449
rect 88708 -16453 88749 -16419
rect 88753 -16453 88760 -16408
rect 88853 -16419 88860 -16408
rect 89034 -16413 89075 -16379
rect 89098 -16413 89150 -16379
rect 89178 -16413 89219 -16379
rect 88864 -16453 88905 -16419
rect 88510 -16494 88551 -16460
rect 88160 -16534 88201 -16500
rect 88160 -16568 88165 -16534
rect 86810 -16740 86815 -16706
rect 87106 -16723 87147 -16689
rect 87151 -16723 87158 -16681
rect 87293 -16741 87305 -16673
rect 87334 -16707 87339 -16639
rect 87379 -16671 87384 -16603
rect 87413 -16637 87418 -16571
rect 88354 -16577 88395 -16543
rect 88399 -16577 88406 -16532
rect 88499 -16543 88506 -16532
rect 88708 -16537 88749 -16503
rect 88753 -16537 88760 -16492
rect 88853 -16503 88860 -16492
rect 89098 -16496 89139 -16462
rect 89143 -16496 89150 -16451
rect 88864 -16537 88905 -16503
rect 88510 -16577 88551 -16543
rect 87423 -16621 87464 -16587
rect 87624 -16666 87665 -16632
rect 87393 -16689 87400 -16681
rect 87404 -16723 87445 -16689
rect 87624 -16734 87665 -16700
rect 84557 -16906 84598 -16872
rect 84629 -16906 84670 -16872
rect 84701 -16906 84742 -16872
rect 85014 -16913 85055 -16879
rect 85059 -16913 85066 -16868
rect 85159 -16879 85166 -16868
rect 85170 -16913 85211 -16879
rect 85754 -16895 85795 -16861
rect 85799 -16895 85806 -16853
rect 83648 -16959 84130 -16925
rect 84982 -16949 85023 -16915
rect 85054 -16949 85095 -16915
rect 85368 -16956 85409 -16922
rect 85413 -16956 85420 -16911
rect 85513 -16922 85520 -16911
rect 85941 -16913 85953 -16845
rect 85982 -16879 85987 -16811
rect 86027 -16843 86032 -16775
rect 86061 -16809 86066 -16743
rect 87293 -16753 87300 -16741
rect 87673 -16750 87678 -16616
rect 86071 -16793 86112 -16759
rect 86274 -16838 86315 -16804
rect 86041 -16861 86048 -16853
rect 86052 -16895 86093 -16861
rect 86274 -16906 86315 -16872
rect 85524 -16956 85565 -16922
rect 83648 -16985 84117 -16959
rect 83652 -16993 83859 -16985
rect 83668 -17003 83843 -16993
rect 83394 -17140 83575 -17114
rect 82901 -17174 82942 -17140
rect 82997 -17174 83038 -17140
rect 83093 -17174 83134 -17140
rect 83189 -17174 83230 -17140
rect 83285 -17174 83326 -17140
rect 83381 -17174 83575 -17140
rect 83394 -17200 83575 -17174
rect 83594 -17174 83701 -17050
rect 83853 -17062 83859 -17051
rect 83472 -17870 83513 -17200
rect 83594 -17228 83603 -17174
rect 83279 -17936 83430 -17924
rect 82947 -17970 83430 -17936
rect 83279 -17971 83430 -17970
rect 83460 -17971 83513 -17870
rect 83606 -17971 83647 -17174
rect 83652 -17971 83658 -17174
rect 83864 -17971 83905 -17062
rect 83998 -17971 84039 -16985
rect 84251 -17002 84292 -16968
rect 84347 -17002 84388 -16968
rect 84443 -17002 84484 -16968
rect 84539 -17002 84580 -16968
rect 84635 -17002 84676 -16968
rect 84731 -17002 84772 -16968
rect 84827 -17002 84868 -16968
rect 85336 -16992 85377 -16958
rect 85408 -16992 85449 -16958
rect 85754 -16995 85795 -16961
rect 85799 -16995 85806 -16950
rect 85941 -17001 85948 -16913
rect 86323 -16922 86328 -16788
rect 86041 -16961 86048 -16950
rect 86357 -16956 86362 -16762
rect 86397 -16778 86404 -16767
rect 86393 -16809 86404 -16778
rect 86719 -16796 86760 -16762
rect 86052 -16995 86093 -16961
rect 84989 -17045 85030 -17011
rect 85085 -17045 85126 -17011
rect 85181 -17045 85222 -17011
rect 85690 -17035 85731 -17001
rect 85762 -17035 85803 -17001
rect 85834 -17035 85875 -17001
rect 85906 -17029 85948 -17001
rect 86252 -17025 86293 -16991
rect 86297 -17025 86304 -16980
rect 86393 -16992 86398 -16809
rect 86427 -16995 86432 -16812
rect 85906 -17035 85947 -17029
rect 85343 -17088 85384 -17054
rect 85439 -17088 85480 -17054
rect 85535 -17088 85576 -17054
rect 86439 -17076 86446 -16809
rect 87068 -16819 87461 -16753
rect 87707 -16784 87712 -16590
rect 87747 -16606 87754 -16595
rect 87743 -16637 87754 -16606
rect 88069 -16624 88110 -16590
rect 86455 -16860 86496 -16826
rect 86804 -16830 86821 -16819
rect 86804 -16832 86810 -16830
rect 86455 -16928 86496 -16894
rect 86507 -16995 86512 -16860
rect 86738 -16874 86810 -16832
rect 86866 -16874 87461 -16819
rect 87602 -16853 87643 -16819
rect 87647 -16853 87654 -16808
rect 87743 -16820 87748 -16637
rect 87777 -16823 87782 -16640
rect 86738 -16877 87461 -16874
rect 86541 -16980 86546 -16892
rect 86658 -16942 86699 -16908
rect 86703 -16942 86710 -16900
rect 86539 -16991 86546 -16980
rect 86541 -17025 86546 -16991
rect 86550 -17025 86591 -16991
rect 86658 -17042 86699 -17008
rect 86703 -17042 86710 -16997
rect 86551 -17078 86592 -17044
rect 86623 -17078 86664 -17044
rect 86695 -17078 86736 -17044
rect 85697 -17131 85738 -17097
rect 85793 -17131 85834 -17097
rect 85889 -17131 85930 -17097
rect 85985 -17131 86026 -17097
rect 86081 -17131 86122 -17097
rect 86738 -17114 86889 -16877
rect 87068 -16899 87461 -16877
rect 86992 -16925 87461 -16899
rect 87789 -16904 87796 -16637
rect 87805 -16688 87846 -16654
rect 87805 -16756 87846 -16722
rect 87857 -16823 87862 -16688
rect 88419 -16691 88460 -16657
rect 88471 -16718 88476 -16641
rect 87891 -16808 87896 -16720
rect 88008 -16770 88049 -16736
rect 88053 -16770 88060 -16728
rect 88153 -16740 88160 -16729
rect 88164 -16774 88205 -16740
rect 88505 -16752 88510 -16607
rect 88708 -16620 88749 -16586
rect 88753 -16620 88760 -16575
rect 88853 -16586 88860 -16575
rect 89098 -16580 89139 -16546
rect 89143 -16580 89150 -16535
rect 88864 -16620 88905 -16586
rect 88773 -16734 88814 -16700
rect 88825 -16761 88830 -16684
rect 87889 -16819 87896 -16808
rect 88358 -16813 88399 -16779
rect 88403 -16813 88410 -16771
rect 88503 -16779 88510 -16771
rect 88514 -16813 88555 -16779
rect 88859 -16795 88864 -16650
rect 89098 -16663 89139 -16629
rect 89143 -16663 89150 -16618
rect 89220 -16679 89225 -16363
rect 89243 -16379 89250 -16371
rect 89254 -16379 89259 -16363
rect 89254 -16413 89295 -16379
rect 89299 -16413 89306 -16371
rect 89243 -16462 89250 -16451
rect 89254 -16462 89259 -16413
rect 89254 -16496 89295 -16462
rect 89299 -16496 89306 -16451
rect 89243 -16546 89250 -16535
rect 89254 -16546 89259 -16496
rect 89254 -16580 89295 -16546
rect 89299 -16580 89306 -16535
rect 89243 -16629 89250 -16618
rect 89254 -16629 89259 -16580
rect 89254 -16663 89295 -16629
rect 89299 -16663 89306 -16618
rect 89243 -16697 89250 -16671
rect 89254 -16713 89259 -16663
rect 89163 -16777 89204 -16743
rect 87891 -16853 87896 -16819
rect 87900 -16853 87941 -16819
rect 88008 -16870 88049 -16836
rect 88053 -16870 88060 -16825
rect 88153 -16832 88160 -16821
rect 88164 -16866 88205 -16832
rect 88712 -16856 88753 -16822
rect 88757 -16856 88764 -16814
rect 88857 -16822 88864 -16814
rect 88868 -16856 88909 -16822
rect 89285 -16845 89292 -16697
rect 89308 -16713 89311 -16363
rect 89342 -16679 89345 -16363
rect 89399 -16379 89406 -16371
rect 89348 -16413 89389 -16379
rect 89410 -16413 89461 -16379
rect 90120 -16422 90125 -16406
rect 90143 -16422 90150 -16414
rect 90154 -16422 90159 -16406
rect 90450 -16408 90491 -16374
rect 90495 -16408 90502 -16363
rect 89399 -16462 89406 -16451
rect 89580 -16456 89621 -16422
rect 89652 -16456 89693 -16422
rect 89724 -16456 89765 -16422
rect 89868 -16456 89909 -16422
rect 89940 -16456 90053 -16422
rect 90084 -16456 90125 -16422
rect 89410 -16496 89451 -16462
rect 89399 -16546 89406 -16535
rect 89977 -16539 90018 -16505
rect 89410 -16580 89451 -16546
rect 89399 -16629 89406 -16618
rect 89410 -16663 89451 -16629
rect 89642 -16689 89683 -16655
rect 89687 -16689 89694 -16644
rect 89764 -16706 89769 -16588
rect 89787 -16655 89794 -16644
rect 89798 -16655 89803 -16622
rect 89834 -16655 89839 -16622
rect 89798 -16689 89839 -16655
rect 89843 -16689 89850 -16644
rect 89798 -16740 89803 -16689
rect 89834 -16740 89839 -16689
rect 89868 -16706 89873 -16589
rect 89977 -16623 90018 -16589
rect 89977 -16706 90018 -16672
rect 90120 -16706 90125 -16456
rect 90154 -16456 90195 -16422
rect 90143 -16505 90150 -16494
rect 90154 -16505 90159 -16456
rect 90450 -16491 90491 -16457
rect 90495 -16491 90502 -16446
rect 90154 -16539 90195 -16505
rect 90143 -16589 90150 -16578
rect 90154 -16589 90159 -16539
rect 90303 -16565 90412 -16499
rect 90572 -16507 90577 -16191
rect 90595 -16207 90602 -16199
rect 90606 -16207 90611 -16191
rect 90606 -16241 90647 -16207
rect 90651 -16241 90658 -16199
rect 90595 -16290 90602 -16279
rect 90606 -16290 90611 -16241
rect 90606 -16324 90647 -16290
rect 90651 -16324 90658 -16279
rect 90595 -16374 90602 -16363
rect 90606 -16374 90611 -16324
rect 90606 -16408 90647 -16374
rect 90651 -16408 90658 -16363
rect 90595 -16457 90602 -16446
rect 90606 -16457 90611 -16408
rect 90606 -16491 90647 -16457
rect 90651 -16491 90658 -16446
rect 90595 -16525 90602 -16499
rect 90606 -16541 90611 -16491
rect 90154 -16623 90195 -16589
rect 90515 -16605 90556 -16571
rect 90143 -16672 90150 -16661
rect 90154 -16672 90159 -16623
rect 90154 -16706 90195 -16672
rect 90637 -16673 90644 -16525
rect 90660 -16541 90663 -16191
rect 90694 -16507 90697 -16191
rect 90751 -16207 90758 -16199
rect 90700 -16241 90741 -16207
rect 90762 -16241 90813 -16207
rect 91677 -16231 91718 -16197
rect 91773 -16231 91814 -16197
rect 91869 -16231 91910 -16197
rect 93839 -16207 93846 -16199
rect 91470 -16250 91475 -16234
rect 91493 -16250 91500 -16242
rect 91504 -16250 91509 -16234
rect 90751 -16290 90758 -16279
rect 90930 -16284 90971 -16250
rect 91002 -16284 91043 -16250
rect 91074 -16284 91115 -16250
rect 91218 -16284 91259 -16250
rect 91290 -16284 91403 -16250
rect 91434 -16284 91475 -16250
rect 90762 -16324 90803 -16290
rect 90751 -16374 90758 -16363
rect 91327 -16367 91368 -16333
rect 90762 -16408 90803 -16374
rect 90751 -16457 90758 -16446
rect 90762 -16491 90803 -16457
rect 90992 -16517 91033 -16483
rect 91037 -16517 91044 -16472
rect 91114 -16534 91119 -16416
rect 91137 -16483 91144 -16472
rect 91148 -16483 91153 -16450
rect 91184 -16483 91189 -16450
rect 91148 -16517 91189 -16483
rect 91193 -16517 91200 -16472
rect 91148 -16568 91153 -16517
rect 91184 -16568 91189 -16517
rect 91218 -16534 91223 -16417
rect 91327 -16451 91368 -16417
rect 91327 -16534 91368 -16500
rect 91470 -16534 91475 -16284
rect 91504 -16284 91545 -16250
rect 92031 -16274 92072 -16240
rect 92127 -16274 92168 -16240
rect 92223 -16274 92264 -16240
rect 93730 -16241 93771 -16207
rect 93794 -16241 93846 -16207
rect 93874 -16241 93915 -16207
rect 91493 -16333 91500 -16322
rect 91504 -16333 91509 -16284
rect 91743 -16293 91750 -16285
rect 91843 -16293 91850 -16285
rect 91670 -16327 91739 -16293
rect 91742 -16327 91783 -16293
rect 91854 -16327 91895 -16293
rect 92385 -16317 92426 -16283
rect 92481 -16317 92522 -16283
rect 92577 -16317 92618 -16283
rect 92673 -16317 92714 -16283
rect 92769 -16317 92810 -16283
rect 93794 -16324 93835 -16290
rect 93839 -16324 93846 -16279
rect 91504 -16367 91545 -16333
rect 92097 -16336 92104 -16328
rect 92197 -16336 92204 -16328
rect 91493 -16417 91500 -16406
rect 91504 -16417 91509 -16367
rect 91698 -16410 91739 -16376
rect 91743 -16410 91750 -16365
rect 91843 -16376 91850 -16365
rect 92024 -16370 92093 -16336
rect 92096 -16370 92137 -16336
rect 92208 -16370 92249 -16336
rect 92933 -16360 92974 -16326
rect 93029 -16360 93070 -16326
rect 93125 -16360 93166 -16326
rect 93221 -16360 93262 -16326
rect 93317 -16360 93358 -16326
rect 93413 -16360 93454 -16326
rect 93509 -16360 93550 -16326
rect 91854 -16410 91895 -16376
rect 92487 -16379 92494 -16371
rect 91504 -16451 91545 -16417
rect 91493 -16500 91500 -16489
rect 91504 -16500 91509 -16451
rect 91698 -16494 91739 -16460
rect 91743 -16494 91750 -16449
rect 91843 -16460 91850 -16449
rect 92052 -16453 92093 -16419
rect 92097 -16453 92104 -16408
rect 92197 -16419 92204 -16408
rect 92378 -16413 92419 -16379
rect 92442 -16413 92494 -16379
rect 92522 -16413 92563 -16379
rect 92208 -16453 92249 -16419
rect 91854 -16494 91895 -16460
rect 91504 -16534 91545 -16500
rect 91504 -16568 91509 -16534
rect 90154 -16740 90159 -16706
rect 90450 -16723 90491 -16689
rect 90495 -16723 90502 -16681
rect 90637 -16741 90649 -16673
rect 90678 -16707 90683 -16639
rect 90723 -16671 90728 -16603
rect 90757 -16637 90762 -16571
rect 91698 -16577 91739 -16543
rect 91743 -16577 91750 -16532
rect 91843 -16543 91850 -16532
rect 92052 -16537 92093 -16503
rect 92097 -16537 92104 -16492
rect 92197 -16503 92204 -16492
rect 92442 -16496 92483 -16462
rect 92487 -16496 92494 -16451
rect 92208 -16537 92249 -16503
rect 91854 -16577 91895 -16543
rect 90767 -16621 90808 -16587
rect 90968 -16666 91009 -16632
rect 90737 -16689 90744 -16681
rect 90748 -16723 90789 -16689
rect 90968 -16734 91009 -16700
rect 87901 -16906 87942 -16872
rect 87973 -16906 88014 -16872
rect 88045 -16906 88086 -16872
rect 88358 -16913 88399 -16879
rect 88403 -16913 88410 -16868
rect 88503 -16879 88510 -16868
rect 88514 -16913 88555 -16879
rect 89098 -16895 89139 -16861
rect 89143 -16895 89150 -16853
rect 86992 -16959 87474 -16925
rect 88326 -16949 88367 -16915
rect 88398 -16949 88439 -16915
rect 88712 -16956 88753 -16922
rect 88757 -16956 88764 -16911
rect 88857 -16922 88864 -16911
rect 89285 -16913 89297 -16845
rect 89326 -16879 89331 -16811
rect 89371 -16843 89376 -16775
rect 89405 -16809 89410 -16743
rect 90637 -16753 90644 -16741
rect 91017 -16750 91022 -16616
rect 89415 -16793 89456 -16759
rect 89618 -16838 89659 -16804
rect 89385 -16861 89392 -16853
rect 89396 -16895 89437 -16861
rect 89618 -16906 89659 -16872
rect 88868 -16956 88909 -16922
rect 86992 -16985 87461 -16959
rect 86996 -16993 87203 -16985
rect 87012 -17003 87187 -16993
rect 86738 -17140 86919 -17114
rect 86245 -17174 86286 -17140
rect 86341 -17174 86382 -17140
rect 86437 -17174 86478 -17140
rect 86533 -17174 86574 -17140
rect 86629 -17174 86670 -17140
rect 86725 -17174 86919 -17140
rect 86738 -17200 86919 -17174
rect 86938 -17174 87045 -17050
rect 87197 -17062 87203 -17051
rect 86816 -17870 86857 -17200
rect 86938 -17228 86947 -17174
rect 86623 -17936 86774 -17924
rect 86291 -17970 86774 -17936
rect 86623 -17971 86774 -17970
rect 86804 -17971 86857 -17870
rect 86950 -17971 86991 -17174
rect 86996 -17971 87002 -17174
rect 87208 -17971 87249 -17062
rect 87342 -17971 87383 -16985
rect 87595 -17002 87636 -16968
rect 87691 -17002 87732 -16968
rect 87787 -17002 87828 -16968
rect 87883 -17002 87924 -16968
rect 87979 -17002 88020 -16968
rect 88075 -17002 88116 -16968
rect 88171 -17002 88212 -16968
rect 88680 -16992 88721 -16958
rect 88752 -16992 88793 -16958
rect 89098 -16995 89139 -16961
rect 89143 -16995 89150 -16950
rect 89285 -17001 89292 -16913
rect 89667 -16922 89672 -16788
rect 89385 -16961 89392 -16950
rect 89701 -16956 89706 -16762
rect 89741 -16778 89748 -16767
rect 89737 -16809 89748 -16778
rect 90063 -16796 90104 -16762
rect 89396 -16995 89437 -16961
rect 88333 -17045 88374 -17011
rect 88429 -17045 88470 -17011
rect 88525 -17045 88566 -17011
rect 89034 -17035 89075 -17001
rect 89106 -17035 89147 -17001
rect 89178 -17035 89219 -17001
rect 89250 -17029 89292 -17001
rect 89596 -17025 89637 -16991
rect 89641 -17025 89648 -16980
rect 89737 -16992 89742 -16809
rect 89771 -16995 89776 -16812
rect 89250 -17035 89291 -17029
rect 88687 -17088 88728 -17054
rect 88783 -17088 88824 -17054
rect 88879 -17088 88920 -17054
rect 89783 -17076 89790 -16809
rect 90412 -16819 90805 -16753
rect 91051 -16784 91056 -16590
rect 91091 -16606 91098 -16595
rect 91087 -16637 91098 -16606
rect 91413 -16624 91454 -16590
rect 89799 -16860 89840 -16826
rect 90148 -16830 90165 -16819
rect 90148 -16832 90154 -16830
rect 89799 -16928 89840 -16894
rect 89851 -16995 89856 -16860
rect 90082 -16874 90154 -16832
rect 90210 -16874 90805 -16819
rect 90946 -16853 90987 -16819
rect 90991 -16853 90998 -16808
rect 91087 -16820 91092 -16637
rect 91121 -16823 91126 -16640
rect 90082 -16877 90805 -16874
rect 89885 -16980 89890 -16892
rect 90002 -16942 90043 -16908
rect 90047 -16942 90054 -16900
rect 89883 -16991 89890 -16980
rect 89885 -17025 89890 -16991
rect 89894 -17025 89935 -16991
rect 90002 -17042 90043 -17008
rect 90047 -17042 90054 -16997
rect 89895 -17078 89936 -17044
rect 89967 -17078 90008 -17044
rect 90039 -17078 90080 -17044
rect 89041 -17131 89082 -17097
rect 89137 -17131 89178 -17097
rect 89233 -17131 89274 -17097
rect 89329 -17131 89370 -17097
rect 89425 -17131 89466 -17097
rect 90082 -17114 90233 -16877
rect 90412 -16899 90805 -16877
rect 90336 -16925 90805 -16899
rect 91133 -16904 91140 -16637
rect 91149 -16688 91190 -16654
rect 91149 -16756 91190 -16722
rect 91201 -16823 91206 -16688
rect 91763 -16691 91804 -16657
rect 91815 -16718 91820 -16641
rect 91235 -16808 91240 -16720
rect 91352 -16770 91393 -16736
rect 91397 -16770 91404 -16728
rect 91497 -16740 91504 -16729
rect 91508 -16774 91549 -16740
rect 91849 -16752 91854 -16607
rect 92052 -16620 92093 -16586
rect 92097 -16620 92104 -16575
rect 92197 -16586 92204 -16575
rect 92442 -16580 92483 -16546
rect 92487 -16580 92494 -16535
rect 92208 -16620 92249 -16586
rect 92117 -16734 92158 -16700
rect 92169 -16761 92174 -16684
rect 91233 -16819 91240 -16808
rect 91702 -16813 91743 -16779
rect 91747 -16813 91754 -16771
rect 91847 -16779 91854 -16771
rect 91858 -16813 91899 -16779
rect 92203 -16795 92208 -16650
rect 92442 -16663 92483 -16629
rect 92487 -16663 92494 -16618
rect 92564 -16679 92569 -16363
rect 92587 -16379 92594 -16371
rect 92598 -16379 92603 -16363
rect 92598 -16413 92639 -16379
rect 92643 -16413 92650 -16371
rect 92587 -16462 92594 -16451
rect 92598 -16462 92603 -16413
rect 92598 -16496 92639 -16462
rect 92643 -16496 92650 -16451
rect 92587 -16546 92594 -16535
rect 92598 -16546 92603 -16496
rect 92598 -16580 92639 -16546
rect 92643 -16580 92650 -16535
rect 92587 -16629 92594 -16618
rect 92598 -16629 92603 -16580
rect 92598 -16663 92639 -16629
rect 92643 -16663 92650 -16618
rect 92587 -16697 92594 -16671
rect 92598 -16713 92603 -16663
rect 92507 -16777 92548 -16743
rect 91235 -16853 91240 -16819
rect 91244 -16853 91285 -16819
rect 91352 -16870 91393 -16836
rect 91397 -16870 91404 -16825
rect 91497 -16832 91504 -16821
rect 91508 -16866 91549 -16832
rect 92056 -16856 92097 -16822
rect 92101 -16856 92108 -16814
rect 92201 -16822 92208 -16814
rect 92212 -16856 92253 -16822
rect 92629 -16845 92636 -16697
rect 92652 -16713 92655 -16363
rect 92686 -16679 92689 -16363
rect 92743 -16379 92750 -16371
rect 92692 -16413 92733 -16379
rect 92754 -16413 92805 -16379
rect 93464 -16422 93469 -16406
rect 93487 -16422 93494 -16414
rect 93498 -16422 93503 -16406
rect 93794 -16408 93835 -16374
rect 93839 -16408 93846 -16363
rect 92743 -16462 92750 -16451
rect 92924 -16456 92965 -16422
rect 92996 -16456 93037 -16422
rect 93068 -16456 93109 -16422
rect 93212 -16456 93253 -16422
rect 93284 -16456 93397 -16422
rect 93428 -16456 93469 -16422
rect 92754 -16496 92795 -16462
rect 92743 -16546 92750 -16535
rect 93321 -16539 93362 -16505
rect 92754 -16580 92795 -16546
rect 92743 -16629 92750 -16618
rect 92754 -16663 92795 -16629
rect 92986 -16689 93027 -16655
rect 93031 -16689 93038 -16644
rect 93108 -16706 93113 -16588
rect 93131 -16655 93138 -16644
rect 93142 -16655 93147 -16622
rect 93178 -16655 93183 -16622
rect 93142 -16689 93183 -16655
rect 93187 -16689 93194 -16644
rect 93142 -16740 93147 -16689
rect 93178 -16740 93183 -16689
rect 93212 -16706 93217 -16589
rect 93321 -16623 93362 -16589
rect 93321 -16706 93362 -16672
rect 93464 -16706 93469 -16456
rect 93498 -16456 93539 -16422
rect 93487 -16505 93494 -16494
rect 93498 -16505 93503 -16456
rect 93794 -16491 93835 -16457
rect 93839 -16491 93846 -16446
rect 93498 -16539 93539 -16505
rect 93487 -16589 93494 -16578
rect 93498 -16589 93503 -16539
rect 93647 -16565 93756 -16499
rect 93916 -16507 93921 -16191
rect 93939 -16207 93946 -16199
rect 93950 -16207 93955 -16191
rect 93950 -16241 93991 -16207
rect 93995 -16241 94002 -16199
rect 93939 -16290 93946 -16279
rect 93950 -16290 93955 -16241
rect 93950 -16324 93991 -16290
rect 93995 -16324 94002 -16279
rect 93939 -16374 93946 -16363
rect 93950 -16374 93955 -16324
rect 93950 -16408 93991 -16374
rect 93995 -16408 94002 -16363
rect 93939 -16457 93946 -16446
rect 93950 -16457 93955 -16408
rect 93950 -16491 93991 -16457
rect 93995 -16491 94002 -16446
rect 93939 -16525 93946 -16499
rect 93950 -16541 93955 -16491
rect 93498 -16623 93539 -16589
rect 93859 -16605 93900 -16571
rect 93487 -16672 93494 -16661
rect 93498 -16672 93503 -16623
rect 93498 -16706 93539 -16672
rect 93981 -16673 93988 -16525
rect 94004 -16541 94007 -16191
rect 94038 -16507 94041 -16191
rect 94095 -16207 94102 -16199
rect 94044 -16241 94085 -16207
rect 94106 -16241 94157 -16207
rect 95021 -16231 95062 -16197
rect 95117 -16231 95158 -16197
rect 95213 -16231 95254 -16197
rect 97183 -16207 97190 -16199
rect 94814 -16250 94819 -16234
rect 94837 -16250 94844 -16242
rect 94848 -16250 94853 -16234
rect 94095 -16290 94102 -16279
rect 94274 -16284 94315 -16250
rect 94346 -16284 94387 -16250
rect 94418 -16284 94459 -16250
rect 94562 -16284 94603 -16250
rect 94634 -16284 94747 -16250
rect 94778 -16284 94819 -16250
rect 94106 -16324 94147 -16290
rect 94095 -16374 94102 -16363
rect 94671 -16367 94712 -16333
rect 94106 -16408 94147 -16374
rect 94095 -16457 94102 -16446
rect 94106 -16491 94147 -16457
rect 94336 -16517 94377 -16483
rect 94381 -16517 94388 -16472
rect 94458 -16534 94463 -16416
rect 94481 -16483 94488 -16472
rect 94492 -16483 94497 -16450
rect 94528 -16483 94533 -16450
rect 94492 -16517 94533 -16483
rect 94537 -16517 94544 -16472
rect 94492 -16568 94497 -16517
rect 94528 -16568 94533 -16517
rect 94562 -16534 94567 -16417
rect 94671 -16451 94712 -16417
rect 94671 -16534 94712 -16500
rect 94814 -16534 94819 -16284
rect 94848 -16284 94889 -16250
rect 95375 -16274 95416 -16240
rect 95471 -16274 95512 -16240
rect 95567 -16274 95608 -16240
rect 97074 -16241 97115 -16207
rect 97138 -16241 97190 -16207
rect 97218 -16241 97259 -16207
rect 94837 -16333 94844 -16322
rect 94848 -16333 94853 -16284
rect 95087 -16293 95094 -16285
rect 95187 -16293 95194 -16285
rect 95014 -16327 95083 -16293
rect 95086 -16327 95127 -16293
rect 95198 -16327 95239 -16293
rect 95729 -16317 95770 -16283
rect 95825 -16317 95866 -16283
rect 95921 -16317 95962 -16283
rect 96017 -16317 96058 -16283
rect 96113 -16317 96154 -16283
rect 97138 -16324 97179 -16290
rect 97183 -16324 97190 -16279
rect 94848 -16367 94889 -16333
rect 95441 -16336 95448 -16328
rect 95541 -16336 95548 -16328
rect 94837 -16417 94844 -16406
rect 94848 -16417 94853 -16367
rect 95042 -16410 95083 -16376
rect 95087 -16410 95094 -16365
rect 95187 -16376 95194 -16365
rect 95368 -16370 95437 -16336
rect 95440 -16370 95481 -16336
rect 95552 -16370 95593 -16336
rect 96277 -16360 96318 -16326
rect 96373 -16360 96414 -16326
rect 96469 -16360 96510 -16326
rect 96565 -16360 96606 -16326
rect 96661 -16360 96702 -16326
rect 96757 -16360 96798 -16326
rect 96853 -16360 96894 -16326
rect 95198 -16410 95239 -16376
rect 95831 -16379 95838 -16371
rect 94848 -16451 94889 -16417
rect 94837 -16500 94844 -16489
rect 94848 -16500 94853 -16451
rect 95042 -16494 95083 -16460
rect 95087 -16494 95094 -16449
rect 95187 -16460 95194 -16449
rect 95396 -16453 95437 -16419
rect 95441 -16453 95448 -16408
rect 95541 -16419 95548 -16408
rect 95722 -16413 95763 -16379
rect 95786 -16413 95838 -16379
rect 95866 -16413 95907 -16379
rect 95552 -16453 95593 -16419
rect 95198 -16494 95239 -16460
rect 94848 -16534 94889 -16500
rect 94848 -16568 94853 -16534
rect 93498 -16740 93503 -16706
rect 93794 -16723 93835 -16689
rect 93839 -16723 93846 -16681
rect 93981 -16741 93993 -16673
rect 94022 -16707 94027 -16639
rect 94067 -16671 94072 -16603
rect 94101 -16637 94106 -16571
rect 95042 -16577 95083 -16543
rect 95087 -16577 95094 -16532
rect 95187 -16543 95194 -16532
rect 95396 -16537 95437 -16503
rect 95441 -16537 95448 -16492
rect 95541 -16503 95548 -16492
rect 95786 -16496 95827 -16462
rect 95831 -16496 95838 -16451
rect 95552 -16537 95593 -16503
rect 95198 -16577 95239 -16543
rect 94111 -16621 94152 -16587
rect 94312 -16666 94353 -16632
rect 94081 -16689 94088 -16681
rect 94092 -16723 94133 -16689
rect 94312 -16734 94353 -16700
rect 91245 -16906 91286 -16872
rect 91317 -16906 91358 -16872
rect 91389 -16906 91430 -16872
rect 91702 -16913 91743 -16879
rect 91747 -16913 91754 -16868
rect 91847 -16879 91854 -16868
rect 91858 -16913 91899 -16879
rect 92442 -16895 92483 -16861
rect 92487 -16895 92494 -16853
rect 90336 -16959 90818 -16925
rect 91670 -16949 91711 -16915
rect 91742 -16949 91783 -16915
rect 92056 -16956 92097 -16922
rect 92101 -16956 92108 -16911
rect 92201 -16922 92208 -16911
rect 92629 -16913 92641 -16845
rect 92670 -16879 92675 -16811
rect 92715 -16843 92720 -16775
rect 92749 -16809 92754 -16743
rect 93981 -16753 93988 -16741
rect 94361 -16750 94366 -16616
rect 92759 -16793 92800 -16759
rect 92962 -16838 93003 -16804
rect 92729 -16861 92736 -16853
rect 92740 -16895 92781 -16861
rect 92962 -16906 93003 -16872
rect 92212 -16956 92253 -16922
rect 90336 -16985 90805 -16959
rect 90340 -16993 90547 -16985
rect 90356 -17003 90531 -16993
rect 90082 -17140 90263 -17114
rect 89589 -17174 89630 -17140
rect 89685 -17174 89726 -17140
rect 89781 -17174 89822 -17140
rect 89877 -17174 89918 -17140
rect 89973 -17174 90014 -17140
rect 90069 -17174 90263 -17140
rect 90082 -17200 90263 -17174
rect 90282 -17174 90389 -17050
rect 90541 -17062 90547 -17051
rect 90160 -17870 90201 -17200
rect 90282 -17228 90291 -17174
rect 89967 -17936 90118 -17924
rect 89635 -17970 90118 -17936
rect 89967 -17971 90118 -17970
rect 90148 -17971 90201 -17870
rect 90294 -17971 90335 -17174
rect 90340 -17971 90346 -17174
rect 90552 -17971 90593 -17062
rect 90686 -17971 90727 -16985
rect 90939 -17002 90980 -16968
rect 91035 -17002 91076 -16968
rect 91131 -17002 91172 -16968
rect 91227 -17002 91268 -16968
rect 91323 -17002 91364 -16968
rect 91419 -17002 91460 -16968
rect 91515 -17002 91556 -16968
rect 92024 -16992 92065 -16958
rect 92096 -16992 92137 -16958
rect 92442 -16995 92483 -16961
rect 92487 -16995 92494 -16950
rect 92629 -17001 92636 -16913
rect 93011 -16922 93016 -16788
rect 92729 -16961 92736 -16950
rect 93045 -16956 93050 -16762
rect 93085 -16778 93092 -16767
rect 93081 -16809 93092 -16778
rect 93407 -16796 93448 -16762
rect 92740 -16995 92781 -16961
rect 91677 -17045 91718 -17011
rect 91773 -17045 91814 -17011
rect 91869 -17045 91910 -17011
rect 92378 -17035 92419 -17001
rect 92450 -17035 92491 -17001
rect 92522 -17035 92563 -17001
rect 92594 -17029 92636 -17001
rect 92940 -17025 92981 -16991
rect 92985 -17025 92992 -16980
rect 93081 -16992 93086 -16809
rect 93115 -16995 93120 -16812
rect 92594 -17035 92635 -17029
rect 92031 -17088 92072 -17054
rect 92127 -17088 92168 -17054
rect 92223 -17088 92264 -17054
rect 93127 -17076 93134 -16809
rect 93756 -16819 94149 -16753
rect 94395 -16784 94400 -16590
rect 94435 -16606 94442 -16595
rect 94431 -16637 94442 -16606
rect 94757 -16624 94798 -16590
rect 93143 -16860 93184 -16826
rect 93492 -16830 93509 -16819
rect 93492 -16832 93498 -16830
rect 93143 -16928 93184 -16894
rect 93195 -16995 93200 -16860
rect 93426 -16874 93498 -16832
rect 93554 -16874 94149 -16819
rect 94290 -16853 94331 -16819
rect 94335 -16853 94342 -16808
rect 94431 -16820 94436 -16637
rect 94465 -16823 94470 -16640
rect 93426 -16877 94149 -16874
rect 93229 -16980 93234 -16892
rect 93346 -16942 93387 -16908
rect 93391 -16942 93398 -16900
rect 93227 -16991 93234 -16980
rect 93229 -17025 93234 -16991
rect 93238 -17025 93279 -16991
rect 93346 -17042 93387 -17008
rect 93391 -17042 93398 -16997
rect 93239 -17078 93280 -17044
rect 93311 -17078 93352 -17044
rect 93383 -17078 93424 -17044
rect 92385 -17131 92426 -17097
rect 92481 -17131 92522 -17097
rect 92577 -17131 92618 -17097
rect 92673 -17131 92714 -17097
rect 92769 -17131 92810 -17097
rect 93426 -17114 93577 -16877
rect 93756 -16899 94149 -16877
rect 93680 -16925 94149 -16899
rect 94477 -16904 94484 -16637
rect 94493 -16688 94534 -16654
rect 94493 -16756 94534 -16722
rect 94545 -16823 94550 -16688
rect 95107 -16691 95148 -16657
rect 95159 -16718 95164 -16641
rect 94579 -16808 94584 -16720
rect 94696 -16770 94737 -16736
rect 94741 -16770 94748 -16728
rect 94841 -16740 94848 -16729
rect 94852 -16774 94893 -16740
rect 95193 -16752 95198 -16607
rect 95396 -16620 95437 -16586
rect 95441 -16620 95448 -16575
rect 95541 -16586 95548 -16575
rect 95786 -16580 95827 -16546
rect 95831 -16580 95838 -16535
rect 95552 -16620 95593 -16586
rect 95461 -16734 95502 -16700
rect 95513 -16761 95518 -16684
rect 94577 -16819 94584 -16808
rect 95046 -16813 95087 -16779
rect 95091 -16813 95098 -16771
rect 95191 -16779 95198 -16771
rect 95202 -16813 95243 -16779
rect 95547 -16795 95552 -16650
rect 95786 -16663 95827 -16629
rect 95831 -16663 95838 -16618
rect 95908 -16679 95913 -16363
rect 95931 -16379 95938 -16371
rect 95942 -16379 95947 -16363
rect 95942 -16413 95983 -16379
rect 95987 -16413 95994 -16371
rect 95931 -16462 95938 -16451
rect 95942 -16462 95947 -16413
rect 95942 -16496 95983 -16462
rect 95987 -16496 95994 -16451
rect 95931 -16546 95938 -16535
rect 95942 -16546 95947 -16496
rect 95942 -16580 95983 -16546
rect 95987 -16580 95994 -16535
rect 95931 -16629 95938 -16618
rect 95942 -16629 95947 -16580
rect 95942 -16663 95983 -16629
rect 95987 -16663 95994 -16618
rect 95931 -16697 95938 -16671
rect 95942 -16713 95947 -16663
rect 95851 -16777 95892 -16743
rect 94579 -16853 94584 -16819
rect 94588 -16853 94629 -16819
rect 94696 -16870 94737 -16836
rect 94741 -16870 94748 -16825
rect 94841 -16832 94848 -16821
rect 94852 -16866 94893 -16832
rect 95400 -16856 95441 -16822
rect 95445 -16856 95452 -16814
rect 95545 -16822 95552 -16814
rect 95556 -16856 95597 -16822
rect 95973 -16845 95980 -16697
rect 95996 -16713 95999 -16363
rect 96030 -16679 96033 -16363
rect 96087 -16379 96094 -16371
rect 96036 -16413 96077 -16379
rect 96098 -16413 96149 -16379
rect 96808 -16422 96813 -16406
rect 96831 -16422 96838 -16414
rect 96842 -16422 96847 -16406
rect 97138 -16408 97179 -16374
rect 97183 -16408 97190 -16363
rect 96087 -16462 96094 -16451
rect 96268 -16456 96309 -16422
rect 96340 -16456 96381 -16422
rect 96412 -16456 96453 -16422
rect 96556 -16456 96597 -16422
rect 96628 -16456 96741 -16422
rect 96772 -16456 96813 -16422
rect 96098 -16496 96139 -16462
rect 96087 -16546 96094 -16535
rect 96665 -16539 96706 -16505
rect 96098 -16580 96139 -16546
rect 96087 -16629 96094 -16618
rect 96098 -16663 96139 -16629
rect 96330 -16689 96371 -16655
rect 96375 -16689 96382 -16644
rect 96452 -16706 96457 -16588
rect 96475 -16655 96482 -16644
rect 96486 -16655 96491 -16622
rect 96522 -16655 96527 -16622
rect 96486 -16689 96527 -16655
rect 96531 -16689 96538 -16644
rect 96486 -16740 96491 -16689
rect 96522 -16740 96527 -16689
rect 96556 -16706 96561 -16589
rect 96665 -16623 96706 -16589
rect 96665 -16706 96706 -16672
rect 96808 -16706 96813 -16456
rect 96842 -16456 96883 -16422
rect 96831 -16505 96838 -16494
rect 96842 -16505 96847 -16456
rect 97138 -16491 97179 -16457
rect 97183 -16491 97190 -16446
rect 96842 -16539 96883 -16505
rect 96831 -16589 96838 -16578
rect 96842 -16589 96847 -16539
rect 96991 -16565 97100 -16499
rect 97260 -16507 97265 -16191
rect 97283 -16207 97290 -16199
rect 97294 -16207 97299 -16191
rect 97294 -16241 97335 -16207
rect 97339 -16241 97346 -16199
rect 97283 -16290 97290 -16279
rect 97294 -16290 97299 -16241
rect 97294 -16324 97335 -16290
rect 97339 -16324 97346 -16279
rect 97283 -16374 97290 -16363
rect 97294 -16374 97299 -16324
rect 97294 -16408 97335 -16374
rect 97339 -16408 97346 -16363
rect 97283 -16457 97290 -16446
rect 97294 -16457 97299 -16408
rect 97294 -16491 97335 -16457
rect 97339 -16491 97346 -16446
rect 97283 -16525 97290 -16499
rect 97294 -16541 97299 -16491
rect 96842 -16623 96883 -16589
rect 97203 -16605 97244 -16571
rect 96831 -16672 96838 -16661
rect 96842 -16672 96847 -16623
rect 96842 -16706 96883 -16672
rect 97325 -16673 97332 -16525
rect 97348 -16541 97351 -16191
rect 97382 -16507 97385 -16191
rect 97439 -16207 97446 -16199
rect 97388 -16241 97429 -16207
rect 97450 -16241 97501 -16207
rect 98365 -16231 98406 -16197
rect 98461 -16231 98502 -16197
rect 98557 -16231 98598 -16197
rect 100527 -16207 100534 -16199
rect 98158 -16250 98163 -16234
rect 98181 -16250 98188 -16242
rect 98192 -16250 98197 -16234
rect 97439 -16290 97446 -16279
rect 97618 -16284 97659 -16250
rect 97690 -16284 97731 -16250
rect 97762 -16284 97803 -16250
rect 97906 -16284 97947 -16250
rect 97978 -16284 98091 -16250
rect 98122 -16284 98163 -16250
rect 97450 -16324 97491 -16290
rect 97439 -16374 97446 -16363
rect 98015 -16367 98056 -16333
rect 97450 -16408 97491 -16374
rect 97439 -16457 97446 -16446
rect 97450 -16491 97491 -16457
rect 97680 -16517 97721 -16483
rect 97725 -16517 97732 -16472
rect 97802 -16534 97807 -16416
rect 97825 -16483 97832 -16472
rect 97836 -16483 97841 -16450
rect 97872 -16483 97877 -16450
rect 97836 -16517 97877 -16483
rect 97881 -16517 97888 -16472
rect 97836 -16568 97841 -16517
rect 97872 -16568 97877 -16517
rect 97906 -16534 97911 -16417
rect 98015 -16451 98056 -16417
rect 98015 -16534 98056 -16500
rect 98158 -16534 98163 -16284
rect 98192 -16284 98233 -16250
rect 98719 -16274 98760 -16240
rect 98815 -16274 98856 -16240
rect 98911 -16274 98952 -16240
rect 100418 -16241 100459 -16207
rect 100482 -16241 100534 -16207
rect 100562 -16241 100603 -16207
rect 98181 -16333 98188 -16322
rect 98192 -16333 98197 -16284
rect 98431 -16293 98438 -16285
rect 98531 -16293 98538 -16285
rect 98358 -16327 98427 -16293
rect 98430 -16327 98471 -16293
rect 98542 -16327 98583 -16293
rect 99073 -16317 99114 -16283
rect 99169 -16317 99210 -16283
rect 99265 -16317 99306 -16283
rect 99361 -16317 99402 -16283
rect 99457 -16317 99498 -16283
rect 100482 -16324 100523 -16290
rect 100527 -16324 100534 -16279
rect 98192 -16367 98233 -16333
rect 98785 -16336 98792 -16328
rect 98885 -16336 98892 -16328
rect 98181 -16417 98188 -16406
rect 98192 -16417 98197 -16367
rect 98386 -16410 98427 -16376
rect 98431 -16410 98438 -16365
rect 98531 -16376 98538 -16365
rect 98712 -16370 98781 -16336
rect 98784 -16370 98825 -16336
rect 98896 -16370 98937 -16336
rect 99621 -16360 99662 -16326
rect 99717 -16360 99758 -16326
rect 99813 -16360 99854 -16326
rect 99909 -16360 99950 -16326
rect 100005 -16360 100046 -16326
rect 100101 -16360 100142 -16326
rect 100197 -16360 100238 -16326
rect 98542 -16410 98583 -16376
rect 99175 -16379 99182 -16371
rect 98192 -16451 98233 -16417
rect 98181 -16500 98188 -16489
rect 98192 -16500 98197 -16451
rect 98386 -16494 98427 -16460
rect 98431 -16494 98438 -16449
rect 98531 -16460 98538 -16449
rect 98740 -16453 98781 -16419
rect 98785 -16453 98792 -16408
rect 98885 -16419 98892 -16408
rect 99066 -16413 99107 -16379
rect 99130 -16413 99182 -16379
rect 99210 -16413 99251 -16379
rect 98896 -16453 98937 -16419
rect 98542 -16494 98583 -16460
rect 98192 -16534 98233 -16500
rect 98192 -16568 98197 -16534
rect 96842 -16740 96847 -16706
rect 97138 -16723 97179 -16689
rect 97183 -16723 97190 -16681
rect 97325 -16741 97337 -16673
rect 97366 -16707 97371 -16639
rect 97411 -16671 97416 -16603
rect 97445 -16637 97450 -16571
rect 98386 -16577 98427 -16543
rect 98431 -16577 98438 -16532
rect 98531 -16543 98538 -16532
rect 98740 -16537 98781 -16503
rect 98785 -16537 98792 -16492
rect 98885 -16503 98892 -16492
rect 99130 -16496 99171 -16462
rect 99175 -16496 99182 -16451
rect 98896 -16537 98937 -16503
rect 98542 -16577 98583 -16543
rect 97455 -16621 97496 -16587
rect 97656 -16666 97697 -16632
rect 97425 -16689 97432 -16681
rect 97436 -16723 97477 -16689
rect 97656 -16734 97697 -16700
rect 94589 -16906 94630 -16872
rect 94661 -16906 94702 -16872
rect 94733 -16906 94774 -16872
rect 95046 -16913 95087 -16879
rect 95091 -16913 95098 -16868
rect 95191 -16879 95198 -16868
rect 95202 -16913 95243 -16879
rect 95786 -16895 95827 -16861
rect 95831 -16895 95838 -16853
rect 93680 -16959 94162 -16925
rect 95014 -16949 95055 -16915
rect 95086 -16949 95127 -16915
rect 95400 -16956 95441 -16922
rect 95445 -16956 95452 -16911
rect 95545 -16922 95552 -16911
rect 95973 -16913 95985 -16845
rect 96014 -16879 96019 -16811
rect 96059 -16843 96064 -16775
rect 96093 -16809 96098 -16743
rect 97325 -16753 97332 -16741
rect 97705 -16750 97710 -16616
rect 96103 -16793 96144 -16759
rect 96306 -16838 96347 -16804
rect 96073 -16861 96080 -16853
rect 96084 -16895 96125 -16861
rect 96306 -16906 96347 -16872
rect 95556 -16956 95597 -16922
rect 93680 -16985 94149 -16959
rect 93684 -16993 93891 -16985
rect 93700 -17003 93875 -16993
rect 93426 -17140 93607 -17114
rect 92933 -17174 92974 -17140
rect 93029 -17174 93070 -17140
rect 93125 -17174 93166 -17140
rect 93221 -17174 93262 -17140
rect 93317 -17174 93358 -17140
rect 93413 -17174 93607 -17140
rect 93426 -17200 93607 -17174
rect 93626 -17174 93733 -17050
rect 93885 -17062 93891 -17051
rect 93504 -17870 93545 -17200
rect 93626 -17228 93635 -17174
rect 93311 -17936 93462 -17924
rect 92979 -17970 93462 -17936
rect 93311 -17971 93462 -17970
rect 93492 -17971 93545 -17870
rect 93638 -17971 93679 -17174
rect 93684 -17971 93690 -17174
rect 93896 -17971 93937 -17062
rect 94030 -17971 94071 -16985
rect 94283 -17002 94324 -16968
rect 94379 -17002 94420 -16968
rect 94475 -17002 94516 -16968
rect 94571 -17002 94612 -16968
rect 94667 -17002 94708 -16968
rect 94763 -17002 94804 -16968
rect 94859 -17002 94900 -16968
rect 95368 -16992 95409 -16958
rect 95440 -16992 95481 -16958
rect 95786 -16995 95827 -16961
rect 95831 -16995 95838 -16950
rect 95973 -17001 95980 -16913
rect 96355 -16922 96360 -16788
rect 96073 -16961 96080 -16950
rect 96389 -16956 96394 -16762
rect 96429 -16778 96436 -16767
rect 96425 -16809 96436 -16778
rect 96751 -16796 96792 -16762
rect 96084 -16995 96125 -16961
rect 95021 -17045 95062 -17011
rect 95117 -17045 95158 -17011
rect 95213 -17045 95254 -17011
rect 95722 -17035 95763 -17001
rect 95794 -17035 95835 -17001
rect 95866 -17035 95907 -17001
rect 95938 -17029 95980 -17001
rect 96284 -17025 96325 -16991
rect 96329 -17025 96336 -16980
rect 96425 -16992 96430 -16809
rect 96459 -16995 96464 -16812
rect 95938 -17035 95979 -17029
rect 95375 -17088 95416 -17054
rect 95471 -17088 95512 -17054
rect 95567 -17088 95608 -17054
rect 96471 -17076 96478 -16809
rect 97100 -16819 97493 -16753
rect 97739 -16784 97744 -16590
rect 97779 -16606 97786 -16595
rect 97775 -16637 97786 -16606
rect 98101 -16624 98142 -16590
rect 96487 -16860 96528 -16826
rect 96836 -16830 96853 -16819
rect 96836 -16832 96842 -16830
rect 96487 -16928 96528 -16894
rect 96539 -16995 96544 -16860
rect 96770 -16874 96842 -16832
rect 96898 -16874 97493 -16819
rect 97634 -16853 97675 -16819
rect 97679 -16853 97686 -16808
rect 97775 -16820 97780 -16637
rect 97809 -16823 97814 -16640
rect 96770 -16877 97493 -16874
rect 96573 -16980 96578 -16892
rect 96690 -16942 96731 -16908
rect 96735 -16942 96742 -16900
rect 96571 -16991 96578 -16980
rect 96573 -17025 96578 -16991
rect 96582 -17025 96623 -16991
rect 96690 -17042 96731 -17008
rect 96735 -17042 96742 -16997
rect 96583 -17078 96624 -17044
rect 96655 -17078 96696 -17044
rect 96727 -17078 96768 -17044
rect 95729 -17131 95770 -17097
rect 95825 -17131 95866 -17097
rect 95921 -17131 95962 -17097
rect 96017 -17131 96058 -17097
rect 96113 -17131 96154 -17097
rect 96770 -17114 96921 -16877
rect 97100 -16899 97493 -16877
rect 97024 -16925 97493 -16899
rect 97821 -16904 97828 -16637
rect 97837 -16688 97878 -16654
rect 97837 -16756 97878 -16722
rect 97889 -16823 97894 -16688
rect 98451 -16691 98492 -16657
rect 98503 -16718 98508 -16641
rect 97923 -16808 97928 -16720
rect 98040 -16770 98081 -16736
rect 98085 -16770 98092 -16728
rect 98185 -16740 98192 -16729
rect 98196 -16774 98237 -16740
rect 98537 -16752 98542 -16607
rect 98740 -16620 98781 -16586
rect 98785 -16620 98792 -16575
rect 98885 -16586 98892 -16575
rect 99130 -16580 99171 -16546
rect 99175 -16580 99182 -16535
rect 98896 -16620 98937 -16586
rect 98805 -16734 98846 -16700
rect 98857 -16761 98862 -16684
rect 97921 -16819 97928 -16808
rect 98390 -16813 98431 -16779
rect 98435 -16813 98442 -16771
rect 98535 -16779 98542 -16771
rect 98546 -16813 98587 -16779
rect 98891 -16795 98896 -16650
rect 99130 -16663 99171 -16629
rect 99175 -16663 99182 -16618
rect 99252 -16679 99257 -16363
rect 99275 -16379 99282 -16371
rect 99286 -16379 99291 -16363
rect 99286 -16413 99327 -16379
rect 99331 -16413 99338 -16371
rect 99275 -16462 99282 -16451
rect 99286 -16462 99291 -16413
rect 99286 -16496 99327 -16462
rect 99331 -16496 99338 -16451
rect 99275 -16546 99282 -16535
rect 99286 -16546 99291 -16496
rect 99286 -16580 99327 -16546
rect 99331 -16580 99338 -16535
rect 99275 -16629 99282 -16618
rect 99286 -16629 99291 -16580
rect 99286 -16663 99327 -16629
rect 99331 -16663 99338 -16618
rect 99275 -16697 99282 -16671
rect 99286 -16713 99291 -16663
rect 99195 -16777 99236 -16743
rect 97923 -16853 97928 -16819
rect 97932 -16853 97973 -16819
rect 98040 -16870 98081 -16836
rect 98085 -16870 98092 -16825
rect 98185 -16832 98192 -16821
rect 98196 -16866 98237 -16832
rect 98744 -16856 98785 -16822
rect 98789 -16856 98796 -16814
rect 98889 -16822 98896 -16814
rect 98900 -16856 98941 -16822
rect 99317 -16845 99324 -16697
rect 99340 -16713 99343 -16363
rect 99374 -16679 99377 -16363
rect 99431 -16379 99438 -16371
rect 99380 -16413 99421 -16379
rect 99442 -16413 99493 -16379
rect 100152 -16422 100157 -16406
rect 100175 -16422 100182 -16414
rect 100186 -16422 100191 -16406
rect 100482 -16408 100523 -16374
rect 100527 -16408 100534 -16363
rect 99431 -16462 99438 -16451
rect 99612 -16456 99653 -16422
rect 99684 -16456 99725 -16422
rect 99756 -16456 99797 -16422
rect 99900 -16456 99941 -16422
rect 99972 -16456 100085 -16422
rect 100116 -16456 100157 -16422
rect 99442 -16496 99483 -16462
rect 99431 -16546 99438 -16535
rect 100009 -16539 100050 -16505
rect 99442 -16580 99483 -16546
rect 99431 -16629 99438 -16618
rect 99442 -16663 99483 -16629
rect 99674 -16689 99715 -16655
rect 99719 -16689 99726 -16644
rect 99796 -16706 99801 -16588
rect 99819 -16655 99826 -16644
rect 99830 -16655 99835 -16622
rect 99866 -16655 99871 -16622
rect 99830 -16689 99871 -16655
rect 99875 -16689 99882 -16644
rect 99830 -16740 99835 -16689
rect 99866 -16740 99871 -16689
rect 99900 -16706 99905 -16589
rect 100009 -16623 100050 -16589
rect 100009 -16706 100050 -16672
rect 100152 -16706 100157 -16456
rect 100186 -16456 100227 -16422
rect 100175 -16505 100182 -16494
rect 100186 -16505 100191 -16456
rect 100482 -16491 100523 -16457
rect 100527 -16491 100534 -16446
rect 100186 -16539 100227 -16505
rect 100175 -16589 100182 -16578
rect 100186 -16589 100191 -16539
rect 100335 -16565 100444 -16499
rect 100604 -16507 100609 -16191
rect 100627 -16207 100634 -16199
rect 100638 -16207 100643 -16191
rect 100638 -16241 100679 -16207
rect 100683 -16241 100690 -16199
rect 100627 -16290 100634 -16279
rect 100638 -16290 100643 -16241
rect 100638 -16324 100679 -16290
rect 100683 -16324 100690 -16279
rect 100627 -16374 100634 -16363
rect 100638 -16374 100643 -16324
rect 100638 -16408 100679 -16374
rect 100683 -16408 100690 -16363
rect 100627 -16457 100634 -16446
rect 100638 -16457 100643 -16408
rect 100638 -16491 100679 -16457
rect 100683 -16491 100690 -16446
rect 100627 -16525 100634 -16499
rect 100638 -16541 100643 -16491
rect 100186 -16623 100227 -16589
rect 100547 -16605 100588 -16571
rect 100175 -16672 100182 -16661
rect 100186 -16672 100191 -16623
rect 100186 -16706 100227 -16672
rect 100669 -16673 100676 -16525
rect 100692 -16541 100695 -16191
rect 100726 -16507 100729 -16191
rect 100783 -16207 100790 -16199
rect 100732 -16241 100773 -16207
rect 100794 -16241 100845 -16207
rect 101709 -16231 101750 -16197
rect 101805 -16231 101846 -16197
rect 101901 -16231 101942 -16197
rect 103871 -16207 103878 -16199
rect 101502 -16250 101507 -16234
rect 101525 -16250 101532 -16242
rect 101536 -16250 101541 -16234
rect 100783 -16290 100790 -16279
rect 100962 -16284 101003 -16250
rect 101034 -16284 101075 -16250
rect 101106 -16284 101147 -16250
rect 101250 -16284 101291 -16250
rect 101322 -16284 101435 -16250
rect 101466 -16284 101507 -16250
rect 100794 -16324 100835 -16290
rect 100783 -16374 100790 -16363
rect 101359 -16367 101400 -16333
rect 100794 -16408 100835 -16374
rect 100783 -16457 100790 -16446
rect 100794 -16491 100835 -16457
rect 101024 -16517 101065 -16483
rect 101069 -16517 101076 -16472
rect 101146 -16534 101151 -16416
rect 101169 -16483 101176 -16472
rect 101180 -16483 101185 -16450
rect 101216 -16483 101221 -16450
rect 101180 -16517 101221 -16483
rect 101225 -16517 101232 -16472
rect 101180 -16568 101185 -16517
rect 101216 -16568 101221 -16517
rect 101250 -16534 101255 -16417
rect 101359 -16451 101400 -16417
rect 101359 -16534 101400 -16500
rect 101502 -16534 101507 -16284
rect 101536 -16284 101577 -16250
rect 102063 -16274 102104 -16240
rect 102159 -16274 102200 -16240
rect 102255 -16274 102296 -16240
rect 103762 -16241 103803 -16207
rect 103826 -16241 103878 -16207
rect 103906 -16241 103947 -16207
rect 101525 -16333 101532 -16322
rect 101536 -16333 101541 -16284
rect 101775 -16293 101782 -16285
rect 101875 -16293 101882 -16285
rect 101702 -16327 101771 -16293
rect 101774 -16327 101815 -16293
rect 101886 -16327 101927 -16293
rect 102417 -16317 102458 -16283
rect 102513 -16317 102554 -16283
rect 102609 -16317 102650 -16283
rect 102705 -16317 102746 -16283
rect 102801 -16317 102842 -16283
rect 103826 -16324 103867 -16290
rect 103871 -16324 103878 -16279
rect 101536 -16367 101577 -16333
rect 102129 -16336 102136 -16328
rect 102229 -16336 102236 -16328
rect 101525 -16417 101532 -16406
rect 101536 -16417 101541 -16367
rect 101730 -16410 101771 -16376
rect 101775 -16410 101782 -16365
rect 101875 -16376 101882 -16365
rect 102056 -16370 102125 -16336
rect 102128 -16370 102169 -16336
rect 102240 -16370 102281 -16336
rect 102965 -16360 103006 -16326
rect 103061 -16360 103102 -16326
rect 103157 -16360 103198 -16326
rect 103253 -16360 103294 -16326
rect 103349 -16360 103390 -16326
rect 103445 -16360 103486 -16326
rect 103541 -16360 103582 -16326
rect 101886 -16410 101927 -16376
rect 102519 -16379 102526 -16371
rect 101536 -16451 101577 -16417
rect 101525 -16500 101532 -16489
rect 101536 -16500 101541 -16451
rect 101730 -16494 101771 -16460
rect 101775 -16494 101782 -16449
rect 101875 -16460 101882 -16449
rect 102084 -16453 102125 -16419
rect 102129 -16453 102136 -16408
rect 102229 -16419 102236 -16408
rect 102410 -16413 102451 -16379
rect 102474 -16413 102526 -16379
rect 102554 -16413 102595 -16379
rect 102240 -16453 102281 -16419
rect 101886 -16494 101927 -16460
rect 101536 -16534 101577 -16500
rect 101536 -16568 101541 -16534
rect 100186 -16740 100191 -16706
rect 100482 -16723 100523 -16689
rect 100527 -16723 100534 -16681
rect 100669 -16741 100681 -16673
rect 100710 -16707 100715 -16639
rect 100755 -16671 100760 -16603
rect 100789 -16637 100794 -16571
rect 101730 -16577 101771 -16543
rect 101775 -16577 101782 -16532
rect 101875 -16543 101882 -16532
rect 102084 -16537 102125 -16503
rect 102129 -16537 102136 -16492
rect 102229 -16503 102236 -16492
rect 102474 -16496 102515 -16462
rect 102519 -16496 102526 -16451
rect 102240 -16537 102281 -16503
rect 101886 -16577 101927 -16543
rect 100800 -16621 100840 -16587
rect 101000 -16666 101041 -16632
rect 100769 -16689 100776 -16681
rect 100780 -16723 100821 -16689
rect 101000 -16734 101041 -16700
rect 97933 -16906 97974 -16872
rect 98005 -16906 98046 -16872
rect 98077 -16906 98118 -16872
rect 98390 -16913 98431 -16879
rect 98435 -16913 98442 -16868
rect 98535 -16879 98542 -16868
rect 98546 -16913 98587 -16879
rect 99130 -16895 99171 -16861
rect 99175 -16895 99182 -16853
rect 97024 -16959 97506 -16925
rect 98358 -16949 98399 -16915
rect 98430 -16949 98471 -16915
rect 98744 -16956 98785 -16922
rect 98789 -16956 98796 -16911
rect 98889 -16922 98896 -16911
rect 99317 -16913 99329 -16845
rect 99358 -16879 99363 -16811
rect 99403 -16843 99408 -16775
rect 99437 -16809 99442 -16743
rect 100669 -16753 100676 -16741
rect 101049 -16750 101054 -16616
rect 99447 -16793 99488 -16759
rect 99650 -16838 99691 -16804
rect 99417 -16861 99424 -16853
rect 99428 -16895 99469 -16861
rect 99650 -16906 99691 -16872
rect 98900 -16956 98941 -16922
rect 97024 -16985 97493 -16959
rect 97028 -16993 97235 -16985
rect 97044 -17003 97219 -16993
rect 96770 -17140 96951 -17114
rect 96277 -17174 96318 -17140
rect 96373 -17174 96414 -17140
rect 96469 -17174 96510 -17140
rect 96565 -17174 96606 -17140
rect 96661 -17174 96702 -17140
rect 96757 -17174 96951 -17140
rect 96770 -17200 96951 -17174
rect 96970 -17174 97077 -17050
rect 97229 -17062 97235 -17051
rect 96848 -17870 96889 -17200
rect 96970 -17228 96979 -17174
rect 96655 -17936 96806 -17924
rect 96323 -17970 96806 -17936
rect 96655 -17971 96806 -17970
rect 96836 -17971 96889 -17870
rect 96982 -17971 97023 -17174
rect 97028 -17971 97034 -17174
rect 97240 -17971 97281 -17062
rect 97374 -17971 97415 -16985
rect 97627 -17002 97668 -16968
rect 97723 -17002 97764 -16968
rect 97819 -17002 97860 -16968
rect 97915 -17002 97956 -16968
rect 98011 -17002 98052 -16968
rect 98107 -17002 98148 -16968
rect 98203 -17002 98244 -16968
rect 98712 -16992 98753 -16958
rect 98784 -16992 98825 -16958
rect 99130 -16995 99171 -16961
rect 99175 -16995 99182 -16950
rect 99317 -17001 99324 -16913
rect 99699 -16922 99704 -16788
rect 99417 -16961 99424 -16950
rect 99733 -16956 99738 -16762
rect 99773 -16778 99780 -16767
rect 99769 -16809 99780 -16778
rect 100095 -16796 100136 -16762
rect 99428 -16995 99469 -16961
rect 98365 -17045 98406 -17011
rect 98461 -17045 98502 -17011
rect 98557 -17045 98598 -17011
rect 99066 -17035 99107 -17001
rect 99138 -17035 99179 -17001
rect 99210 -17035 99251 -17001
rect 99282 -17029 99324 -17001
rect 99628 -17025 99669 -16991
rect 99673 -17025 99680 -16980
rect 99769 -16992 99774 -16809
rect 99803 -16995 99808 -16812
rect 99282 -17035 99323 -17029
rect 98719 -17088 98760 -17054
rect 98815 -17088 98856 -17054
rect 98911 -17088 98952 -17054
rect 99815 -17076 99822 -16809
rect 100444 -16819 100837 -16753
rect 101083 -16784 101088 -16590
rect 101123 -16606 101130 -16595
rect 101119 -16637 101130 -16606
rect 101445 -16624 101486 -16590
rect 99831 -16860 99872 -16826
rect 100180 -16830 100197 -16819
rect 100180 -16832 100186 -16830
rect 99831 -16928 99872 -16894
rect 99883 -16995 99888 -16860
rect 100114 -16874 100186 -16832
rect 100242 -16874 100837 -16819
rect 100978 -16853 101019 -16819
rect 101023 -16853 101030 -16808
rect 101119 -16820 101124 -16637
rect 101153 -16823 101158 -16640
rect 100114 -16877 100837 -16874
rect 99917 -16980 99922 -16892
rect 100034 -16942 100075 -16908
rect 100079 -16942 100086 -16900
rect 99915 -16991 99922 -16980
rect 99917 -17025 99922 -16991
rect 99926 -17025 99967 -16991
rect 100034 -17042 100075 -17008
rect 100079 -17042 100086 -16997
rect 99927 -17078 99968 -17044
rect 99999 -17078 100040 -17044
rect 100071 -17078 100112 -17044
rect 99073 -17131 99114 -17097
rect 99169 -17131 99210 -17097
rect 99265 -17131 99306 -17097
rect 99361 -17131 99402 -17097
rect 99457 -17131 99498 -17097
rect 100114 -17114 100265 -16877
rect 100444 -16899 100837 -16877
rect 100368 -16925 100837 -16899
rect 101165 -16904 101172 -16637
rect 101181 -16688 101222 -16654
rect 101181 -16756 101222 -16722
rect 101233 -16823 101238 -16688
rect 101795 -16691 101836 -16657
rect 101847 -16718 101852 -16641
rect 101267 -16808 101272 -16720
rect 101384 -16770 101425 -16736
rect 101429 -16770 101436 -16728
rect 101529 -16740 101536 -16729
rect 101540 -16774 101581 -16740
rect 101881 -16752 101886 -16607
rect 102084 -16620 102125 -16586
rect 102129 -16620 102136 -16575
rect 102229 -16586 102236 -16575
rect 102474 -16580 102515 -16546
rect 102519 -16580 102526 -16535
rect 102240 -16620 102281 -16586
rect 102149 -16734 102190 -16700
rect 102201 -16761 102206 -16684
rect 101265 -16819 101272 -16808
rect 101734 -16813 101775 -16779
rect 101779 -16813 101786 -16771
rect 101879 -16779 101886 -16771
rect 101890 -16813 101931 -16779
rect 102235 -16795 102240 -16650
rect 102474 -16663 102515 -16629
rect 102519 -16663 102526 -16618
rect 102596 -16679 102601 -16363
rect 102619 -16379 102626 -16371
rect 102630 -16379 102635 -16363
rect 102630 -16413 102671 -16379
rect 102675 -16413 102682 -16371
rect 102619 -16462 102626 -16451
rect 102630 -16462 102635 -16413
rect 102630 -16496 102671 -16462
rect 102675 -16496 102682 -16451
rect 102619 -16546 102626 -16535
rect 102630 -16546 102635 -16496
rect 102630 -16580 102671 -16546
rect 102675 -16580 102682 -16535
rect 102619 -16629 102626 -16618
rect 102630 -16629 102635 -16580
rect 102630 -16663 102671 -16629
rect 102675 -16663 102682 -16618
rect 102619 -16697 102626 -16671
rect 102630 -16713 102635 -16663
rect 102539 -16777 102580 -16743
rect 101267 -16853 101272 -16819
rect 101276 -16853 101317 -16819
rect 101384 -16870 101425 -16836
rect 101429 -16870 101436 -16825
rect 101529 -16832 101536 -16821
rect 101540 -16866 101581 -16832
rect 102088 -16856 102129 -16822
rect 102133 -16856 102140 -16814
rect 102233 -16822 102240 -16814
rect 102244 -16856 102285 -16822
rect 102661 -16845 102668 -16697
rect 102684 -16713 102687 -16363
rect 102718 -16679 102721 -16363
rect 102775 -16379 102782 -16371
rect 102724 -16413 102765 -16379
rect 102786 -16413 102837 -16379
rect 103496 -16422 103501 -16406
rect 103519 -16422 103526 -16414
rect 103530 -16422 103535 -16406
rect 103826 -16408 103867 -16374
rect 103871 -16408 103878 -16363
rect 102775 -16462 102782 -16451
rect 102956 -16456 102997 -16422
rect 103028 -16456 103069 -16422
rect 103100 -16456 103141 -16422
rect 103244 -16456 103285 -16422
rect 103316 -16456 103429 -16422
rect 103460 -16456 103501 -16422
rect 102786 -16496 102827 -16462
rect 102775 -16546 102782 -16535
rect 103353 -16539 103394 -16505
rect 102786 -16580 102827 -16546
rect 102775 -16629 102782 -16618
rect 102786 -16663 102827 -16629
rect 103018 -16689 103059 -16655
rect 103063 -16689 103070 -16644
rect 103140 -16706 103145 -16588
rect 103163 -16655 103170 -16644
rect 103174 -16655 103179 -16622
rect 103210 -16655 103215 -16622
rect 103174 -16689 103215 -16655
rect 103219 -16689 103226 -16644
rect 103174 -16740 103179 -16689
rect 103210 -16740 103215 -16689
rect 103244 -16706 103249 -16589
rect 103353 -16623 103394 -16589
rect 103353 -16706 103394 -16672
rect 103496 -16706 103501 -16456
rect 103530 -16456 103571 -16422
rect 103519 -16505 103526 -16494
rect 103530 -16505 103535 -16456
rect 103826 -16491 103867 -16457
rect 103871 -16491 103878 -16446
rect 103530 -16539 103571 -16505
rect 103519 -16589 103526 -16578
rect 103530 -16589 103535 -16539
rect 103679 -16565 103788 -16499
rect 103948 -16507 103953 -16191
rect 103971 -16207 103978 -16199
rect 103982 -16207 103987 -16191
rect 103982 -16241 104023 -16207
rect 104027 -16241 104034 -16199
rect 103971 -16290 103978 -16279
rect 103982 -16290 103987 -16241
rect 103982 -16324 104023 -16290
rect 104027 -16324 104034 -16279
rect 103971 -16374 103978 -16363
rect 103982 -16374 103987 -16324
rect 103982 -16408 104023 -16374
rect 104027 -16408 104034 -16363
rect 103971 -16457 103978 -16446
rect 103982 -16457 103987 -16408
rect 103982 -16491 104023 -16457
rect 104027 -16491 104034 -16446
rect 103971 -16525 103978 -16499
rect 103982 -16541 103987 -16491
rect 103530 -16623 103571 -16589
rect 103891 -16605 103932 -16571
rect 103519 -16672 103526 -16661
rect 103530 -16672 103535 -16623
rect 103530 -16706 103571 -16672
rect 104013 -16673 104020 -16525
rect 104036 -16541 104039 -16191
rect 104070 -16507 104073 -16191
rect 104127 -16207 104134 -16199
rect 104076 -16241 104117 -16207
rect 104138 -16241 104189 -16207
rect 105053 -16231 105094 -16197
rect 105149 -16231 105190 -16197
rect 105245 -16231 105286 -16197
rect 104846 -16250 104851 -16234
rect 104869 -16250 104876 -16242
rect 104880 -16250 104885 -16234
rect 104127 -16290 104134 -16279
rect 104306 -16284 104347 -16250
rect 104378 -16284 104419 -16250
rect 104450 -16284 104491 -16250
rect 104594 -16284 104635 -16250
rect 104666 -16284 104779 -16250
rect 104810 -16284 104851 -16250
rect 104138 -16324 104179 -16290
rect 104127 -16374 104134 -16363
rect 104703 -16367 104744 -16333
rect 104138 -16408 104179 -16374
rect 104127 -16457 104134 -16446
rect 104138 -16491 104179 -16457
rect 104368 -16517 104409 -16483
rect 104413 -16517 104420 -16472
rect 104490 -16534 104495 -16416
rect 104513 -16483 104520 -16472
rect 104524 -16483 104529 -16450
rect 104560 -16483 104565 -16450
rect 104524 -16517 104565 -16483
rect 104569 -16517 104576 -16472
rect 104524 -16568 104529 -16517
rect 104560 -16568 104565 -16517
rect 104594 -16534 104599 -16417
rect 104703 -16451 104744 -16417
rect 104703 -16534 104744 -16500
rect 104846 -16534 104851 -16284
rect 104880 -16284 104921 -16250
rect 105407 -16274 105448 -16240
rect 105503 -16274 105544 -16240
rect 105599 -16274 105640 -16240
rect 107112 -16241 107147 -16207
rect 107176 -16241 107219 -16207
rect 107221 -16241 107222 -16199
rect 107321 -16207 107322 -16199
rect 107256 -16241 107291 -16207
rect 107332 -16241 107367 -16207
rect 107377 -16241 107378 -16199
rect 107477 -16207 107478 -16199
rect 107426 -16241 107461 -16207
rect 107488 -16241 107533 -16207
rect 108403 -16231 108438 -16197
rect 108499 -16231 108534 -16197
rect 108595 -16231 108630 -16197
rect 108219 -16250 108220 -16242
rect 104869 -16333 104876 -16322
rect 104880 -16333 104885 -16284
rect 105119 -16293 105126 -16285
rect 105219 -16293 105226 -16285
rect 105046 -16327 105115 -16293
rect 105118 -16327 105159 -16293
rect 105230 -16327 105271 -16293
rect 105761 -16317 105802 -16283
rect 105857 -16317 105898 -16283
rect 105953 -16317 105994 -16283
rect 106049 -16317 106090 -16283
rect 106145 -16317 106186 -16283
rect 107176 -16324 107211 -16290
rect 107221 -16324 107222 -16279
rect 107321 -16290 107322 -16279
rect 107332 -16324 107367 -16290
rect 107377 -16324 107378 -16279
rect 107477 -16290 107478 -16279
rect 107656 -16284 107691 -16250
rect 107728 -16284 107763 -16250
rect 107800 -16284 107835 -16250
rect 107944 -16284 107979 -16250
rect 108016 -16284 108051 -16250
rect 108053 -16284 108123 -16250
rect 108160 -16284 108195 -16250
rect 108230 -16284 108265 -16250
rect 108757 -16274 108792 -16240
rect 108853 -16274 108888 -16240
rect 108949 -16274 108984 -16240
rect 110456 -16241 110491 -16207
rect 110520 -16241 110563 -16207
rect 110565 -16241 110566 -16199
rect 110665 -16207 110666 -16199
rect 110600 -16241 110635 -16207
rect 110676 -16241 110711 -16207
rect 110721 -16241 110722 -16199
rect 110821 -16207 110822 -16199
rect 110770 -16241 110805 -16207
rect 110832 -16241 110877 -16207
rect 111747 -16231 111782 -16197
rect 111843 -16231 111878 -16197
rect 111939 -16231 111974 -16197
rect 111563 -16250 111564 -16242
rect 107488 -16324 107523 -16290
rect 108469 -16293 108470 -16285
rect 108569 -16293 108570 -16285
rect 104880 -16367 104921 -16333
rect 105473 -16336 105480 -16328
rect 105573 -16336 105580 -16328
rect 104869 -16417 104876 -16406
rect 104880 -16417 104885 -16367
rect 105074 -16410 105115 -16376
rect 105119 -16410 105126 -16365
rect 105219 -16376 105226 -16365
rect 105400 -16370 105469 -16336
rect 105472 -16370 105513 -16336
rect 105584 -16370 105625 -16336
rect 106309 -16360 106350 -16326
rect 106405 -16360 106446 -16326
rect 106501 -16360 106542 -16326
rect 106597 -16360 106638 -16326
rect 106693 -16360 106734 -16326
rect 106789 -16360 106830 -16326
rect 106885 -16360 106926 -16326
rect 108219 -16333 108220 -16322
rect 108396 -16327 108459 -16293
rect 108468 -16327 108503 -16293
rect 108580 -16327 108615 -16293
rect 109111 -16317 109146 -16283
rect 109207 -16317 109242 -16283
rect 109303 -16317 109338 -16283
rect 109399 -16317 109434 -16283
rect 109495 -16317 109530 -16283
rect 110520 -16324 110555 -16290
rect 110565 -16324 110566 -16279
rect 110665 -16290 110666 -16279
rect 110676 -16324 110711 -16290
rect 110721 -16324 110722 -16279
rect 110821 -16290 110822 -16279
rect 111000 -16284 111035 -16250
rect 111072 -16284 111107 -16250
rect 111144 -16284 111179 -16250
rect 111288 -16284 111323 -16250
rect 111360 -16284 111395 -16250
rect 111397 -16284 111467 -16250
rect 111504 -16284 111539 -16250
rect 111574 -16284 111609 -16250
rect 112101 -16274 112136 -16240
rect 112197 -16274 112232 -16240
rect 112293 -16274 112328 -16240
rect 113800 -16241 113835 -16207
rect 113864 -16241 113907 -16207
rect 113909 -16241 113910 -16199
rect 114009 -16207 114010 -16199
rect 113944 -16241 113979 -16207
rect 114020 -16241 114055 -16207
rect 114065 -16241 114066 -16199
rect 114165 -16207 114166 -16199
rect 114114 -16241 114149 -16207
rect 114176 -16241 114221 -16207
rect 115091 -16231 115126 -16197
rect 115187 -16231 115222 -16197
rect 115283 -16231 115318 -16197
rect 114907 -16250 114908 -16242
rect 110832 -16324 110867 -16290
rect 111813 -16293 111814 -16285
rect 111913 -16293 111914 -16285
rect 105230 -16410 105271 -16376
rect 105863 -16379 105870 -16371
rect 104880 -16451 104921 -16417
rect 104869 -16500 104876 -16489
rect 104880 -16500 104885 -16451
rect 105074 -16494 105115 -16460
rect 105119 -16494 105126 -16449
rect 105219 -16460 105226 -16449
rect 105428 -16453 105469 -16419
rect 105473 -16453 105480 -16408
rect 105573 -16419 105580 -16408
rect 105754 -16413 105795 -16379
rect 105818 -16413 105870 -16379
rect 105898 -16413 105939 -16379
rect 105584 -16453 105625 -16419
rect 105230 -16494 105271 -16460
rect 104880 -16534 104921 -16500
rect 104880 -16568 104885 -16534
rect 103530 -16740 103535 -16706
rect 103826 -16723 103867 -16689
rect 103871 -16723 103878 -16681
rect 104013 -16741 104025 -16673
rect 104054 -16707 104059 -16639
rect 104099 -16671 104104 -16603
rect 104133 -16637 104138 -16571
rect 105074 -16577 105115 -16543
rect 105119 -16577 105126 -16532
rect 105219 -16543 105226 -16532
rect 105428 -16537 105469 -16503
rect 105473 -16537 105480 -16492
rect 105573 -16503 105580 -16492
rect 105818 -16496 105859 -16462
rect 105863 -16496 105870 -16451
rect 105584 -16537 105625 -16503
rect 105230 -16577 105271 -16543
rect 104143 -16621 104184 -16587
rect 104344 -16666 104385 -16632
rect 104113 -16689 104120 -16681
rect 104124 -16723 104165 -16689
rect 104344 -16734 104385 -16700
rect 101277 -16906 101318 -16872
rect 101349 -16906 101390 -16872
rect 101421 -16906 101462 -16872
rect 101734 -16913 101775 -16879
rect 101779 -16913 101786 -16868
rect 101879 -16879 101886 -16868
rect 101890 -16913 101931 -16879
rect 102474 -16895 102515 -16861
rect 102519 -16895 102526 -16853
rect 100368 -16959 100850 -16925
rect 101702 -16949 101743 -16915
rect 101774 -16949 101815 -16915
rect 102088 -16956 102129 -16922
rect 102133 -16956 102140 -16911
rect 102233 -16922 102240 -16911
rect 102661 -16913 102673 -16845
rect 102702 -16879 102707 -16811
rect 102747 -16843 102752 -16775
rect 102781 -16809 102786 -16743
rect 104013 -16753 104020 -16741
rect 104393 -16750 104398 -16616
rect 102791 -16793 102832 -16759
rect 102994 -16838 103035 -16804
rect 102761 -16861 102768 -16853
rect 102772 -16895 102813 -16861
rect 102994 -16906 103035 -16872
rect 102244 -16956 102285 -16922
rect 100368 -16985 100837 -16959
rect 100372 -16993 100579 -16985
rect 100388 -17003 100563 -16993
rect 100114 -17140 100295 -17114
rect 99621 -17174 99662 -17140
rect 99717 -17174 99758 -17140
rect 99813 -17174 99854 -17140
rect 99909 -17174 99950 -17140
rect 100005 -17174 100046 -17140
rect 100101 -17174 100295 -17140
rect 100114 -17200 100295 -17174
rect 100314 -17174 100421 -17050
rect 100573 -17062 100579 -17051
rect 100192 -17870 100233 -17200
rect 100314 -17228 100323 -17174
rect 99999 -17936 100150 -17924
rect 99667 -17970 100150 -17936
rect 99999 -17971 100150 -17970
rect 100180 -17971 100233 -17870
rect 100326 -17971 100367 -17174
rect 100372 -17971 100378 -17174
rect 100584 -17971 100625 -17062
rect 100718 -17971 100759 -16985
rect 100971 -17002 101012 -16968
rect 101067 -17002 101108 -16968
rect 101163 -17002 101204 -16968
rect 101259 -17002 101300 -16968
rect 101355 -17002 101396 -16968
rect 101451 -17002 101492 -16968
rect 101547 -17002 101588 -16968
rect 102056 -16992 102097 -16958
rect 102128 -16992 102169 -16958
rect 102474 -16995 102515 -16961
rect 102519 -16995 102526 -16950
rect 102661 -17001 102668 -16913
rect 103043 -16922 103048 -16788
rect 102761 -16961 102768 -16950
rect 103077 -16956 103082 -16762
rect 103117 -16778 103124 -16767
rect 103113 -16809 103124 -16778
rect 103439 -16796 103480 -16762
rect 102772 -16995 102813 -16961
rect 101709 -17045 101750 -17011
rect 101805 -17045 101846 -17011
rect 101901 -17045 101942 -17011
rect 102410 -17035 102451 -17001
rect 102482 -17035 102523 -17001
rect 102554 -17035 102595 -17001
rect 102626 -17029 102668 -17001
rect 102972 -17025 103013 -16991
rect 103017 -17025 103024 -16980
rect 103113 -16992 103118 -16809
rect 103147 -16995 103152 -16812
rect 102626 -17035 102667 -17029
rect 102063 -17088 102104 -17054
rect 102159 -17088 102200 -17054
rect 102255 -17088 102296 -17054
rect 103159 -17076 103166 -16809
rect 103788 -16819 104181 -16753
rect 104427 -16784 104432 -16590
rect 104467 -16606 104474 -16595
rect 104463 -16637 104474 -16606
rect 104789 -16624 104830 -16590
rect 103175 -16860 103216 -16826
rect 103524 -16830 103541 -16819
rect 103524 -16832 103530 -16830
rect 103175 -16928 103216 -16894
rect 103227 -16995 103232 -16860
rect 103458 -16874 103530 -16832
rect 103586 -16874 104181 -16819
rect 104322 -16853 104363 -16819
rect 104367 -16853 104374 -16808
rect 104463 -16820 104468 -16637
rect 104497 -16823 104502 -16640
rect 103458 -16877 104181 -16874
rect 103261 -16980 103266 -16892
rect 103378 -16942 103419 -16908
rect 103423 -16942 103430 -16900
rect 103259 -16991 103266 -16980
rect 103261 -17025 103266 -16991
rect 103270 -17025 103311 -16991
rect 103378 -17042 103419 -17008
rect 103423 -17042 103430 -16997
rect 103271 -17078 103312 -17044
rect 103343 -17078 103384 -17044
rect 103415 -17078 103456 -17044
rect 102417 -17131 102458 -17097
rect 102513 -17131 102554 -17097
rect 102609 -17131 102650 -17097
rect 102705 -17131 102746 -17097
rect 102801 -17131 102842 -17097
rect 103458 -17114 103609 -16877
rect 103788 -16899 104181 -16877
rect 103712 -16925 104181 -16899
rect 104509 -16904 104516 -16637
rect 104525 -16688 104566 -16654
rect 104525 -16756 104566 -16722
rect 104577 -16823 104582 -16688
rect 105139 -16691 105180 -16657
rect 105191 -16718 105196 -16641
rect 104611 -16808 104616 -16720
rect 104728 -16770 104769 -16736
rect 104773 -16770 104780 -16728
rect 104873 -16740 104880 -16729
rect 104884 -16774 104925 -16740
rect 105225 -16752 105230 -16607
rect 105428 -16620 105469 -16586
rect 105473 -16620 105480 -16575
rect 105573 -16586 105580 -16575
rect 105818 -16580 105859 -16546
rect 105863 -16580 105870 -16535
rect 105584 -16620 105625 -16586
rect 105493 -16734 105534 -16700
rect 105545 -16761 105550 -16684
rect 104609 -16819 104616 -16808
rect 105078 -16813 105119 -16779
rect 105123 -16813 105130 -16771
rect 105223 -16779 105230 -16771
rect 105234 -16813 105275 -16779
rect 105579 -16795 105584 -16650
rect 105818 -16663 105859 -16629
rect 105863 -16663 105870 -16618
rect 105940 -16679 105945 -16363
rect 105963 -16379 105970 -16371
rect 105974 -16379 105979 -16363
rect 105974 -16413 106015 -16379
rect 106019 -16413 106026 -16371
rect 105963 -16462 105970 -16451
rect 105974 -16462 105979 -16413
rect 105974 -16496 106015 -16462
rect 106019 -16496 106026 -16451
rect 105963 -16546 105970 -16535
rect 105974 -16546 105979 -16496
rect 105974 -16580 106015 -16546
rect 106019 -16580 106026 -16535
rect 105963 -16629 105970 -16618
rect 105974 -16629 105979 -16580
rect 105974 -16663 106015 -16629
rect 106019 -16663 106026 -16618
rect 105963 -16697 105970 -16671
rect 105974 -16713 105979 -16663
rect 105883 -16777 105924 -16743
rect 104611 -16853 104616 -16819
rect 104620 -16853 104661 -16819
rect 104728 -16870 104769 -16836
rect 104773 -16870 104780 -16825
rect 104873 -16832 104880 -16821
rect 104884 -16866 104925 -16832
rect 105432 -16856 105473 -16822
rect 105477 -16856 105484 -16814
rect 105577 -16822 105584 -16814
rect 105588 -16856 105629 -16822
rect 106005 -16845 106012 -16697
rect 106028 -16713 106031 -16363
rect 106062 -16679 106065 -16363
rect 106119 -16379 106126 -16371
rect 106068 -16413 106109 -16379
rect 106130 -16413 106181 -16379
rect 106840 -16422 106845 -16406
rect 106863 -16422 106870 -16414
rect 106874 -16422 106879 -16406
rect 107176 -16408 107211 -16374
rect 107221 -16408 107222 -16363
rect 107321 -16374 107322 -16363
rect 107332 -16408 107367 -16374
rect 107377 -16408 107378 -16363
rect 107477 -16374 107478 -16363
rect 108053 -16367 108088 -16333
rect 108230 -16367 108265 -16333
rect 108823 -16336 108824 -16328
rect 108923 -16336 108924 -16328
rect 107488 -16408 107523 -16374
rect 108219 -16417 108220 -16406
rect 108424 -16410 108459 -16376
rect 108469 -16410 108470 -16365
rect 108569 -16376 108570 -16365
rect 108750 -16370 108813 -16336
rect 108822 -16370 108857 -16336
rect 108934 -16370 108969 -16336
rect 109659 -16360 109694 -16326
rect 109755 -16360 109790 -16326
rect 109851 -16360 109886 -16326
rect 109947 -16360 109982 -16326
rect 110043 -16360 110078 -16326
rect 110139 -16360 110174 -16326
rect 110235 -16360 110270 -16326
rect 111563 -16333 111564 -16322
rect 111740 -16327 111803 -16293
rect 111812 -16327 111847 -16293
rect 111924 -16327 111959 -16293
rect 112455 -16317 112490 -16283
rect 112551 -16317 112586 -16283
rect 112647 -16317 112682 -16283
rect 112743 -16317 112778 -16283
rect 112839 -16317 112874 -16283
rect 113864 -16324 113899 -16290
rect 113909 -16324 113910 -16279
rect 114009 -16290 114010 -16279
rect 114020 -16324 114055 -16290
rect 114065 -16324 114066 -16279
rect 114165 -16290 114166 -16279
rect 114344 -16284 114379 -16250
rect 114416 -16284 114451 -16250
rect 114488 -16284 114523 -16250
rect 114632 -16284 114667 -16250
rect 114704 -16284 114739 -16250
rect 114741 -16284 114811 -16250
rect 114848 -16284 114883 -16250
rect 114918 -16284 114953 -16250
rect 115445 -16274 115480 -16240
rect 115541 -16274 115576 -16240
rect 115637 -16274 115672 -16240
rect 117144 -16241 117179 -16207
rect 117208 -16241 117251 -16207
rect 117253 -16241 117254 -16199
rect 117353 -16207 117354 -16199
rect 117288 -16241 117323 -16207
rect 117364 -16241 117399 -16207
rect 117409 -16241 117410 -16199
rect 117509 -16207 117510 -16199
rect 117458 -16241 117493 -16207
rect 117520 -16241 117565 -16207
rect 118435 -16231 118470 -16197
rect 118531 -16231 118566 -16197
rect 118627 -16231 118662 -16197
rect 118251 -16250 118252 -16242
rect 114176 -16324 114211 -16290
rect 115157 -16293 115158 -16285
rect 115257 -16293 115258 -16285
rect 108580 -16410 108615 -16376
rect 106119 -16462 106126 -16451
rect 106300 -16456 106341 -16422
rect 106372 -16456 106413 -16422
rect 106444 -16456 106485 -16422
rect 106588 -16456 106629 -16422
rect 106660 -16456 106773 -16422
rect 106804 -16456 106845 -16422
rect 106130 -16496 106171 -16462
rect 106119 -16546 106126 -16535
rect 106697 -16539 106738 -16505
rect 106130 -16580 106171 -16546
rect 106119 -16629 106126 -16618
rect 106130 -16663 106171 -16629
rect 106362 -16689 106403 -16655
rect 106407 -16689 106414 -16644
rect 106484 -16706 106489 -16588
rect 106507 -16655 106514 -16644
rect 106518 -16655 106523 -16622
rect 106554 -16655 106559 -16622
rect 106518 -16689 106559 -16655
rect 106563 -16689 106570 -16644
rect 106518 -16740 106523 -16689
rect 106554 -16740 106559 -16689
rect 106588 -16706 106593 -16589
rect 106697 -16623 106738 -16589
rect 106697 -16706 106738 -16672
rect 106840 -16706 106845 -16456
rect 106874 -16456 106915 -16422
rect 106863 -16505 106870 -16494
rect 106874 -16505 106879 -16456
rect 107176 -16491 107211 -16457
rect 107221 -16491 107222 -16446
rect 107321 -16457 107322 -16446
rect 107332 -16491 107367 -16457
rect 107377 -16491 107378 -16446
rect 107477 -16457 107478 -16446
rect 108053 -16451 108088 -16417
rect 108230 -16451 108265 -16417
rect 107488 -16491 107523 -16457
rect 106874 -16539 106915 -16505
rect 106863 -16589 106870 -16578
rect 106874 -16589 106879 -16539
rect 107023 -16565 107138 -16499
rect 107321 -16525 107322 -16499
rect 107718 -16517 107753 -16483
rect 107763 -16517 107764 -16472
rect 107863 -16483 107864 -16472
rect 107874 -16517 107909 -16483
rect 107919 -16517 107920 -16472
rect 108219 -16500 108220 -16489
rect 108424 -16494 108459 -16460
rect 108469 -16494 108470 -16449
rect 108569 -16460 108570 -16449
rect 108778 -16453 108813 -16419
rect 108823 -16453 108824 -16408
rect 108923 -16419 108924 -16408
rect 109104 -16413 109139 -16379
rect 109168 -16413 109211 -16379
rect 109213 -16413 109214 -16371
rect 109313 -16379 109314 -16371
rect 109248 -16413 109283 -16379
rect 109324 -16413 109359 -16379
rect 109369 -16413 109370 -16371
rect 109469 -16379 109470 -16371
rect 109418 -16413 109453 -16379
rect 109480 -16413 109525 -16379
rect 110520 -16408 110555 -16374
rect 110565 -16408 110566 -16363
rect 110665 -16374 110666 -16363
rect 110676 -16408 110711 -16374
rect 110721 -16408 110722 -16363
rect 110821 -16374 110822 -16363
rect 111397 -16367 111432 -16333
rect 111574 -16367 111609 -16333
rect 112167 -16336 112168 -16328
rect 112267 -16336 112268 -16328
rect 110832 -16408 110867 -16374
rect 108934 -16453 108969 -16419
rect 110213 -16422 110214 -16414
rect 111563 -16417 111564 -16406
rect 111768 -16410 111803 -16376
rect 111813 -16410 111814 -16365
rect 111913 -16376 111914 -16365
rect 112094 -16370 112157 -16336
rect 112166 -16370 112201 -16336
rect 112278 -16370 112313 -16336
rect 113003 -16360 113038 -16326
rect 113099 -16360 113134 -16326
rect 113195 -16360 113230 -16326
rect 113291 -16360 113326 -16326
rect 113387 -16360 113422 -16326
rect 113483 -16360 113518 -16326
rect 113579 -16360 113614 -16326
rect 114907 -16333 114908 -16322
rect 115084 -16327 115147 -16293
rect 115156 -16327 115191 -16293
rect 115268 -16327 115303 -16293
rect 115799 -16317 115834 -16283
rect 115895 -16317 115930 -16283
rect 115991 -16317 116026 -16283
rect 116087 -16317 116122 -16283
rect 116183 -16317 116218 -16283
rect 117208 -16324 117243 -16290
rect 117253 -16324 117254 -16279
rect 117353 -16290 117354 -16279
rect 117364 -16324 117399 -16290
rect 117409 -16324 117410 -16279
rect 117509 -16290 117510 -16279
rect 117688 -16284 117723 -16250
rect 117760 -16284 117795 -16250
rect 117832 -16284 117867 -16250
rect 117976 -16284 118011 -16250
rect 118048 -16284 118083 -16250
rect 118085 -16284 118155 -16250
rect 118192 -16284 118227 -16250
rect 118262 -16284 118297 -16250
rect 118789 -16274 118824 -16240
rect 118885 -16274 118920 -16240
rect 118981 -16274 119016 -16240
rect 120488 -16241 120523 -16207
rect 120552 -16241 120595 -16207
rect 120597 -16241 120598 -16199
rect 120697 -16207 120698 -16199
rect 120632 -16241 120667 -16207
rect 120708 -16241 120743 -16207
rect 120753 -16241 120754 -16199
rect 120853 -16207 120854 -16199
rect 120802 -16241 120837 -16207
rect 120864 -16241 120909 -16207
rect 121779 -16231 121814 -16197
rect 121875 -16231 121910 -16197
rect 121971 -16231 122006 -16197
rect 121595 -16250 121596 -16242
rect 117520 -16324 117555 -16290
rect 118501 -16293 118502 -16285
rect 118601 -16293 118602 -16285
rect 111924 -16410 111959 -16376
rect 108580 -16494 108615 -16460
rect 106874 -16623 106915 -16589
rect 107241 -16605 107276 -16571
rect 106863 -16672 106870 -16661
rect 106874 -16672 106879 -16623
rect 106874 -16706 106915 -16672
rect 106874 -16740 106879 -16706
rect 107176 -16723 107211 -16689
rect 107221 -16723 107222 -16681
rect 104621 -16906 104662 -16872
rect 104693 -16906 104734 -16872
rect 104765 -16906 104806 -16872
rect 105078 -16913 105119 -16879
rect 105123 -16913 105130 -16868
rect 105223 -16879 105230 -16868
rect 105234 -16913 105275 -16879
rect 105818 -16895 105859 -16861
rect 105863 -16895 105870 -16853
rect 103712 -16959 104194 -16925
rect 105046 -16949 105087 -16915
rect 105118 -16949 105159 -16915
rect 105432 -16956 105473 -16922
rect 105477 -16956 105484 -16911
rect 105577 -16922 105584 -16911
rect 106005 -16913 106017 -16845
rect 106046 -16879 106051 -16811
rect 106091 -16843 106096 -16775
rect 106125 -16809 106130 -16743
rect 107363 -16753 107364 -16525
rect 108053 -16534 108088 -16500
rect 108230 -16534 108265 -16500
rect 108424 -16577 108459 -16543
rect 108469 -16577 108470 -16532
rect 108569 -16543 108570 -16532
rect 108778 -16537 108813 -16503
rect 108823 -16537 108824 -16492
rect 108923 -16503 108924 -16492
rect 109168 -16496 109203 -16462
rect 109213 -16496 109214 -16451
rect 109313 -16462 109314 -16451
rect 109324 -16496 109359 -16462
rect 109369 -16496 109370 -16451
rect 109469 -16462 109470 -16451
rect 109650 -16456 109685 -16422
rect 109722 -16456 109757 -16422
rect 109794 -16456 109829 -16422
rect 109938 -16456 109973 -16422
rect 110010 -16456 110045 -16422
rect 110047 -16456 110117 -16422
rect 110154 -16456 110189 -16422
rect 110224 -16456 110259 -16422
rect 109480 -16496 109515 -16462
rect 110520 -16491 110555 -16457
rect 110565 -16491 110566 -16446
rect 110665 -16457 110666 -16446
rect 110676 -16491 110711 -16457
rect 110721 -16491 110722 -16446
rect 110821 -16457 110822 -16446
rect 111397 -16451 111432 -16417
rect 111574 -16451 111609 -16417
rect 110832 -16491 110867 -16457
rect 108934 -16537 108969 -16503
rect 110213 -16505 110214 -16494
rect 108580 -16577 108615 -16543
rect 107493 -16621 107528 -16587
rect 107694 -16666 107729 -16632
rect 107817 -16637 107818 -16595
rect 108139 -16624 108174 -16590
rect 108778 -16620 108813 -16586
rect 108823 -16620 108824 -16575
rect 108923 -16586 108924 -16575
rect 109168 -16580 109203 -16546
rect 109213 -16580 109214 -16535
rect 109313 -16546 109314 -16535
rect 109324 -16580 109359 -16546
rect 109369 -16580 109370 -16535
rect 109469 -16546 109470 -16535
rect 110047 -16539 110082 -16505
rect 110224 -16539 110259 -16505
rect 109480 -16580 109515 -16546
rect 110367 -16565 110482 -16499
rect 110665 -16525 110666 -16499
rect 111062 -16517 111097 -16483
rect 111107 -16517 111108 -16472
rect 111207 -16483 111208 -16472
rect 111218 -16517 111253 -16483
rect 111263 -16517 111264 -16472
rect 111563 -16500 111564 -16489
rect 111768 -16494 111803 -16460
rect 111813 -16494 111814 -16449
rect 111913 -16460 111914 -16449
rect 112122 -16453 112157 -16419
rect 112167 -16453 112168 -16408
rect 112267 -16419 112268 -16408
rect 112448 -16413 112483 -16379
rect 112512 -16413 112555 -16379
rect 112557 -16413 112558 -16371
rect 112657 -16379 112658 -16371
rect 112592 -16413 112627 -16379
rect 112668 -16413 112703 -16379
rect 112713 -16413 112714 -16371
rect 112813 -16379 112814 -16371
rect 112762 -16413 112797 -16379
rect 112824 -16413 112869 -16379
rect 113864 -16408 113899 -16374
rect 113909 -16408 113910 -16363
rect 114009 -16374 114010 -16363
rect 114020 -16408 114055 -16374
rect 114065 -16408 114066 -16363
rect 114165 -16374 114166 -16363
rect 114741 -16367 114776 -16333
rect 114918 -16367 114953 -16333
rect 115511 -16336 115512 -16328
rect 115611 -16336 115612 -16328
rect 114176 -16408 114211 -16374
rect 112278 -16453 112313 -16419
rect 113557 -16422 113558 -16414
rect 114907 -16417 114908 -16406
rect 115112 -16410 115147 -16376
rect 115157 -16410 115158 -16365
rect 115257 -16376 115258 -16365
rect 115438 -16370 115501 -16336
rect 115510 -16370 115545 -16336
rect 115622 -16370 115657 -16336
rect 116347 -16360 116382 -16326
rect 116443 -16360 116478 -16326
rect 116539 -16360 116574 -16326
rect 116635 -16360 116670 -16326
rect 116731 -16360 116766 -16326
rect 116827 -16360 116862 -16326
rect 116923 -16360 116958 -16326
rect 118251 -16333 118252 -16322
rect 118428 -16327 118491 -16293
rect 118500 -16327 118535 -16293
rect 118612 -16327 118647 -16293
rect 119143 -16317 119178 -16283
rect 119239 -16317 119274 -16283
rect 119335 -16317 119370 -16283
rect 119431 -16317 119466 -16283
rect 119527 -16317 119562 -16283
rect 120552 -16324 120587 -16290
rect 120597 -16324 120598 -16279
rect 120697 -16290 120698 -16279
rect 120708 -16324 120743 -16290
rect 120753 -16324 120754 -16279
rect 120853 -16290 120854 -16279
rect 121032 -16284 121067 -16250
rect 121104 -16284 121139 -16250
rect 121176 -16284 121211 -16250
rect 121320 -16284 121355 -16250
rect 121392 -16284 121427 -16250
rect 121429 -16284 121499 -16250
rect 121536 -16284 121571 -16250
rect 121606 -16284 121641 -16250
rect 122133 -16274 122168 -16240
rect 122229 -16274 122264 -16240
rect 122325 -16274 122360 -16240
rect 123832 -16241 123867 -16207
rect 123896 -16241 123939 -16207
rect 123941 -16241 123942 -16199
rect 124041 -16207 124042 -16199
rect 123976 -16241 124011 -16207
rect 124052 -16241 124087 -16207
rect 124097 -16241 124098 -16199
rect 124197 -16207 124198 -16199
rect 124146 -16241 124181 -16207
rect 124208 -16241 124253 -16207
rect 125123 -16231 125158 -16197
rect 125219 -16231 125254 -16197
rect 125315 -16231 125350 -16197
rect 124939 -16250 124940 -16242
rect 120864 -16324 120899 -16290
rect 121845 -16293 121846 -16285
rect 121945 -16293 121946 -16285
rect 115268 -16410 115303 -16376
rect 111924 -16494 111959 -16460
rect 108934 -16620 108969 -16586
rect 110213 -16589 110214 -16578
rect 107463 -16689 107464 -16681
rect 107474 -16723 107509 -16689
rect 107694 -16734 107729 -16700
rect 106135 -16793 106176 -16759
rect 106338 -16838 106379 -16804
rect 106105 -16861 106112 -16853
rect 106116 -16895 106157 -16861
rect 106338 -16906 106379 -16872
rect 105588 -16956 105629 -16922
rect 103712 -16985 104181 -16959
rect 103716 -16993 103923 -16985
rect 103732 -17003 103907 -16993
rect 103458 -17140 103639 -17114
rect 102965 -17174 103006 -17140
rect 103061 -17174 103102 -17140
rect 103157 -17174 103198 -17140
rect 103253 -17174 103294 -17140
rect 103349 -17174 103390 -17140
rect 103445 -17174 103639 -17140
rect 103458 -17200 103639 -17174
rect 103658 -17174 103765 -17050
rect 103917 -17062 103923 -17051
rect 103536 -17870 103577 -17200
rect 103658 -17228 103667 -17174
rect 103343 -17936 103494 -17924
rect 103011 -17970 103494 -17936
rect 103343 -17971 103494 -17970
rect 103524 -17971 103577 -17870
rect 103670 -17971 103711 -17174
rect 103716 -17971 103722 -17174
rect 103928 -17971 103969 -17062
rect 104062 -17971 104103 -16985
rect 104315 -17002 104356 -16968
rect 104411 -17002 104452 -16968
rect 104507 -17002 104548 -16968
rect 104603 -17002 104644 -16968
rect 104699 -17002 104740 -16968
rect 104795 -17002 104836 -16968
rect 104891 -17002 104932 -16968
rect 105400 -16992 105441 -16958
rect 105472 -16992 105513 -16958
rect 105818 -16995 105859 -16961
rect 105863 -16995 105870 -16950
rect 106005 -17001 106012 -16913
rect 106387 -16922 106392 -16788
rect 106105 -16961 106112 -16950
rect 106421 -16956 106426 -16762
rect 106461 -16778 106468 -16767
rect 106457 -16809 106468 -16778
rect 106783 -16796 106824 -16762
rect 106116 -16995 106157 -16961
rect 105053 -17045 105094 -17011
rect 105149 -17045 105190 -17011
rect 105245 -17045 105286 -17011
rect 105754 -17035 105795 -17001
rect 105826 -17035 105867 -17001
rect 105898 -17035 105939 -17001
rect 105970 -17029 106012 -17001
rect 106316 -17025 106357 -16991
rect 106361 -17025 106368 -16980
rect 106457 -16992 106462 -16809
rect 106491 -16995 106496 -16812
rect 105970 -17035 106011 -17029
rect 105407 -17088 105448 -17054
rect 105503 -17088 105544 -17054
rect 105599 -17088 105640 -17054
rect 106503 -17076 106510 -16809
rect 107138 -16819 107525 -16753
rect 106519 -16860 106560 -16826
rect 106868 -16830 106885 -16819
rect 106868 -16832 106874 -16830
rect 106519 -16928 106560 -16894
rect 106571 -16995 106576 -16860
rect 106802 -16874 106874 -16832
rect 106936 -16874 107525 -16819
rect 107672 -16853 107707 -16819
rect 107717 -16853 107718 -16808
rect 106802 -16877 107525 -16874
rect 106605 -16980 106610 -16892
rect 106722 -16942 106763 -16908
rect 106767 -16942 106774 -16900
rect 106603 -16991 106610 -16980
rect 106605 -17025 106610 -16991
rect 106614 -17025 106655 -16991
rect 106722 -17042 106763 -17008
rect 106767 -17042 106774 -16997
rect 106615 -17078 106656 -17044
rect 106687 -17078 106728 -17044
rect 106759 -17078 106800 -17044
rect 105761 -17131 105802 -17097
rect 105857 -17131 105898 -17097
rect 105953 -17131 105994 -17097
rect 106049 -17131 106090 -17097
rect 106145 -17131 106186 -17097
rect 106802 -17114 106953 -16877
rect 107138 -16899 107525 -16877
rect 107062 -16925 107525 -16899
rect 107859 -16904 107860 -16637
rect 107875 -16688 107910 -16654
rect 108489 -16691 108524 -16657
rect 109168 -16663 109203 -16629
rect 109213 -16663 109214 -16618
rect 109313 -16629 109314 -16618
rect 109324 -16663 109359 -16629
rect 109369 -16663 109370 -16618
rect 109469 -16629 109470 -16618
rect 110047 -16623 110082 -16589
rect 110224 -16623 110259 -16589
rect 110585 -16605 110620 -16571
rect 109480 -16663 109515 -16629
rect 109313 -16697 109314 -16671
rect 109712 -16689 109747 -16655
rect 109757 -16689 109758 -16644
rect 109857 -16655 109858 -16644
rect 109868 -16689 109903 -16655
rect 109913 -16689 109914 -16644
rect 110213 -16672 110214 -16661
rect 107875 -16756 107910 -16722
rect 108078 -16770 108113 -16736
rect 108123 -16770 108124 -16728
rect 108223 -16740 108224 -16729
rect 108843 -16734 108878 -16700
rect 108234 -16774 108269 -16740
rect 107959 -16819 107960 -16808
rect 108428 -16813 108463 -16779
rect 108473 -16813 108474 -16771
rect 108573 -16779 108574 -16771
rect 109233 -16777 109268 -16743
rect 108584 -16813 108619 -16779
rect 107970 -16853 108005 -16819
rect 108078 -16870 108113 -16836
rect 108123 -16870 108124 -16825
rect 108223 -16832 108224 -16821
rect 108234 -16866 108269 -16832
rect 108782 -16856 108817 -16822
rect 108827 -16856 108828 -16814
rect 108927 -16822 108928 -16814
rect 108938 -16856 108973 -16822
rect 107971 -16906 108006 -16872
rect 108043 -16906 108078 -16872
rect 108115 -16906 108150 -16872
rect 108428 -16913 108463 -16879
rect 108473 -16913 108474 -16868
rect 108573 -16879 108574 -16868
rect 108584 -16913 108619 -16879
rect 109168 -16895 109203 -16861
rect 109213 -16895 109214 -16853
rect 107062 -16959 107538 -16925
rect 108396 -16949 108431 -16915
rect 108468 -16949 108503 -16915
rect 108782 -16956 108817 -16922
rect 108827 -16956 108828 -16911
rect 108927 -16922 108928 -16911
rect 108938 -16956 108973 -16922
rect 107062 -16969 107525 -16959
rect 107060 -16985 107525 -16969
rect 107060 -16993 107267 -16985
rect 107076 -17003 107251 -16993
rect 106802 -17140 106983 -17114
rect 106309 -17174 106350 -17140
rect 106405 -17174 106446 -17140
rect 106501 -17174 106542 -17140
rect 106597 -17174 106638 -17140
rect 106693 -17174 106734 -17140
rect 106789 -17174 106983 -17140
rect 106802 -17200 106983 -17174
rect 107002 -17174 107109 -17050
rect 107261 -17062 107267 -17051
rect 106880 -17870 106921 -17200
rect 107002 -17228 107011 -17174
rect 106687 -17936 106838 -17924
rect 106355 -17970 106838 -17936
rect 106687 -17971 106838 -17970
rect 106868 -17971 106921 -17870
rect 107014 -17971 107055 -17174
rect 107060 -17971 107066 -17174
rect 107272 -17971 107313 -17062
rect 107406 -17971 107447 -16985
rect 107665 -17002 107700 -16968
rect 107761 -17002 107796 -16968
rect 107857 -17002 107892 -16968
rect 107953 -17002 107988 -16968
rect 108049 -17002 108084 -16968
rect 108145 -17002 108180 -16968
rect 108241 -17002 108276 -16968
rect 108750 -16992 108785 -16958
rect 108822 -16992 108857 -16958
rect 109168 -16995 109203 -16961
rect 109213 -16995 109214 -16950
rect 109355 -17001 109356 -16697
rect 110047 -16706 110082 -16672
rect 110224 -16706 110259 -16672
rect 110520 -16723 110555 -16689
rect 110565 -16723 110566 -16681
rect 110707 -16753 110708 -16525
rect 111397 -16534 111432 -16500
rect 111574 -16534 111609 -16500
rect 111768 -16577 111803 -16543
rect 111813 -16577 111814 -16532
rect 111913 -16543 111914 -16532
rect 112122 -16537 112157 -16503
rect 112167 -16537 112168 -16492
rect 112267 -16503 112268 -16492
rect 112512 -16496 112547 -16462
rect 112557 -16496 112558 -16451
rect 112657 -16462 112658 -16451
rect 112668 -16496 112703 -16462
rect 112713 -16496 112714 -16451
rect 112813 -16462 112814 -16451
rect 112994 -16456 113029 -16422
rect 113066 -16456 113101 -16422
rect 113138 -16456 113173 -16422
rect 113282 -16456 113317 -16422
rect 113354 -16456 113389 -16422
rect 113391 -16456 113461 -16422
rect 113498 -16456 113533 -16422
rect 113568 -16456 113603 -16422
rect 112824 -16496 112859 -16462
rect 113864 -16491 113899 -16457
rect 113909 -16491 113910 -16446
rect 114009 -16457 114010 -16446
rect 114020 -16491 114055 -16457
rect 114065 -16491 114066 -16446
rect 114165 -16457 114166 -16446
rect 114741 -16451 114776 -16417
rect 114918 -16451 114953 -16417
rect 114176 -16491 114211 -16457
rect 112278 -16537 112313 -16503
rect 113557 -16505 113558 -16494
rect 111924 -16577 111959 -16543
rect 110837 -16621 110872 -16587
rect 111038 -16666 111073 -16632
rect 111161 -16637 111162 -16595
rect 111483 -16624 111518 -16590
rect 112122 -16620 112157 -16586
rect 112167 -16620 112168 -16575
rect 112267 -16586 112268 -16575
rect 112512 -16580 112547 -16546
rect 112557 -16580 112558 -16535
rect 112657 -16546 112658 -16535
rect 112668 -16580 112703 -16546
rect 112713 -16580 112714 -16535
rect 112813 -16546 112814 -16535
rect 113391 -16539 113426 -16505
rect 113568 -16539 113603 -16505
rect 112824 -16580 112859 -16546
rect 113711 -16565 113826 -16499
rect 114009 -16525 114010 -16499
rect 114406 -16517 114441 -16483
rect 114451 -16517 114452 -16472
rect 114551 -16483 114552 -16472
rect 114562 -16517 114597 -16483
rect 114607 -16517 114608 -16472
rect 114907 -16500 114908 -16489
rect 115112 -16494 115147 -16460
rect 115157 -16494 115158 -16449
rect 115257 -16460 115258 -16449
rect 115466 -16453 115501 -16419
rect 115511 -16453 115512 -16408
rect 115611 -16419 115612 -16408
rect 115792 -16413 115827 -16379
rect 115856 -16413 115899 -16379
rect 115901 -16413 115902 -16371
rect 116001 -16379 116002 -16371
rect 115936 -16413 115971 -16379
rect 116012 -16413 116047 -16379
rect 116057 -16413 116058 -16371
rect 116157 -16379 116158 -16371
rect 116106 -16413 116141 -16379
rect 116168 -16413 116213 -16379
rect 117208 -16408 117243 -16374
rect 117253 -16408 117254 -16363
rect 117353 -16374 117354 -16363
rect 117364 -16408 117399 -16374
rect 117409 -16408 117410 -16363
rect 117509 -16374 117510 -16363
rect 118085 -16367 118120 -16333
rect 118262 -16367 118297 -16333
rect 118855 -16336 118856 -16328
rect 118955 -16336 118956 -16328
rect 117520 -16408 117555 -16374
rect 115622 -16453 115657 -16419
rect 116901 -16422 116902 -16414
rect 118251 -16417 118252 -16406
rect 118456 -16410 118491 -16376
rect 118501 -16410 118502 -16365
rect 118601 -16376 118602 -16365
rect 118782 -16370 118845 -16336
rect 118854 -16370 118889 -16336
rect 118966 -16370 119001 -16336
rect 119691 -16360 119726 -16326
rect 119787 -16360 119822 -16326
rect 119883 -16360 119918 -16326
rect 119979 -16360 120014 -16326
rect 120075 -16360 120110 -16326
rect 120171 -16360 120206 -16326
rect 120267 -16360 120302 -16326
rect 121595 -16333 121596 -16322
rect 121772 -16327 121835 -16293
rect 121844 -16327 121879 -16293
rect 121956 -16327 121991 -16293
rect 122487 -16317 122522 -16283
rect 122583 -16317 122618 -16283
rect 122679 -16317 122714 -16283
rect 122775 -16317 122810 -16283
rect 122871 -16317 122906 -16283
rect 123896 -16324 123931 -16290
rect 123941 -16324 123942 -16279
rect 124041 -16290 124042 -16279
rect 124052 -16324 124087 -16290
rect 124097 -16324 124098 -16279
rect 124197 -16290 124198 -16279
rect 124376 -16284 124411 -16250
rect 124448 -16284 124483 -16250
rect 124520 -16284 124555 -16250
rect 124664 -16284 124699 -16250
rect 124736 -16284 124771 -16250
rect 124773 -16284 124843 -16250
rect 124880 -16284 124915 -16250
rect 124950 -16284 124985 -16250
rect 125477 -16274 125512 -16240
rect 125573 -16274 125608 -16240
rect 125669 -16274 125704 -16240
rect 127176 -16241 127211 -16207
rect 127240 -16241 127283 -16207
rect 127285 -16241 127286 -16199
rect 127385 -16207 127386 -16199
rect 127320 -16241 127355 -16207
rect 127396 -16241 127431 -16207
rect 127441 -16241 127442 -16199
rect 127541 -16207 127542 -16199
rect 127490 -16241 127525 -16207
rect 127552 -16241 127597 -16207
rect 128467 -16231 128502 -16197
rect 128563 -16231 128598 -16197
rect 128659 -16231 128694 -16197
rect 128283 -16250 128284 -16242
rect 124208 -16324 124243 -16290
rect 125189 -16293 125190 -16285
rect 125289 -16293 125290 -16285
rect 118612 -16410 118647 -16376
rect 115268 -16494 115303 -16460
rect 112278 -16620 112313 -16586
rect 113557 -16589 113558 -16578
rect 110807 -16689 110808 -16681
rect 110818 -16723 110853 -16689
rect 111038 -16734 111073 -16700
rect 109485 -16793 109520 -16759
rect 109688 -16838 109723 -16804
rect 109811 -16809 109812 -16767
rect 110133 -16796 110168 -16762
rect 109455 -16861 109456 -16853
rect 109466 -16895 109501 -16861
rect 109688 -16906 109723 -16872
rect 109455 -16961 109456 -16950
rect 109466 -16995 109501 -16961
rect 108403 -17045 108438 -17011
rect 108499 -17045 108534 -17011
rect 108595 -17045 108630 -17011
rect 109104 -17035 109139 -17001
rect 109176 -17035 109211 -17001
rect 109248 -17035 109283 -17001
rect 109320 -17029 109356 -17001
rect 109666 -17025 109701 -16991
rect 109711 -17025 109712 -16980
rect 109320 -17035 109355 -17029
rect 108757 -17088 108792 -17054
rect 108853 -17088 108888 -17054
rect 108949 -17088 108984 -17054
rect 109853 -17076 109854 -16809
rect 110482 -16819 110869 -16753
rect 109869 -16860 109904 -16826
rect 110218 -16832 110229 -16819
rect 110152 -16874 110229 -16832
rect 110280 -16874 110869 -16819
rect 111016 -16853 111051 -16819
rect 111061 -16853 111062 -16808
rect 110152 -16877 110869 -16874
rect 109869 -16928 109904 -16894
rect 110072 -16942 110107 -16908
rect 110117 -16942 110118 -16900
rect 109953 -16991 109954 -16980
rect 109964 -17025 109999 -16991
rect 110072 -17042 110107 -17008
rect 110117 -17042 110118 -16997
rect 109965 -17078 110000 -17044
rect 110037 -17078 110072 -17044
rect 110109 -17078 110144 -17044
rect 109111 -17131 109146 -17097
rect 109207 -17131 109242 -17097
rect 109303 -17131 109338 -17097
rect 109399 -17131 109434 -17097
rect 109495 -17131 109530 -17097
rect 110152 -17114 110297 -16877
rect 110482 -16899 110869 -16877
rect 110406 -16925 110869 -16899
rect 111203 -16904 111204 -16637
rect 111219 -16688 111254 -16654
rect 111833 -16691 111868 -16657
rect 112512 -16663 112547 -16629
rect 112557 -16663 112558 -16618
rect 112657 -16629 112658 -16618
rect 112668 -16663 112703 -16629
rect 112713 -16663 112714 -16618
rect 112813 -16629 112814 -16618
rect 113391 -16623 113426 -16589
rect 113568 -16623 113603 -16589
rect 113929 -16605 113964 -16571
rect 112824 -16663 112859 -16629
rect 112657 -16697 112658 -16671
rect 113056 -16689 113091 -16655
rect 113101 -16689 113102 -16644
rect 113201 -16655 113202 -16644
rect 113212 -16689 113247 -16655
rect 113257 -16689 113258 -16644
rect 113557 -16672 113558 -16661
rect 111219 -16756 111254 -16722
rect 111422 -16770 111457 -16736
rect 111467 -16770 111468 -16728
rect 111567 -16740 111568 -16729
rect 112187 -16734 112222 -16700
rect 111578 -16774 111613 -16740
rect 111303 -16819 111304 -16808
rect 111772 -16813 111807 -16779
rect 111817 -16813 111818 -16771
rect 111917 -16779 111918 -16771
rect 112577 -16777 112612 -16743
rect 111928 -16813 111963 -16779
rect 111314 -16853 111349 -16819
rect 111422 -16870 111457 -16836
rect 111467 -16870 111468 -16825
rect 111567 -16832 111568 -16821
rect 111578 -16866 111613 -16832
rect 112126 -16856 112161 -16822
rect 112171 -16856 112172 -16814
rect 112271 -16822 112272 -16814
rect 112282 -16856 112317 -16822
rect 111315 -16906 111350 -16872
rect 111387 -16906 111422 -16872
rect 111459 -16906 111494 -16872
rect 111772 -16913 111807 -16879
rect 111817 -16913 111818 -16868
rect 111917 -16879 111918 -16868
rect 111928 -16913 111963 -16879
rect 112512 -16895 112547 -16861
rect 112557 -16895 112558 -16853
rect 110406 -16959 110882 -16925
rect 111740 -16949 111775 -16915
rect 111812 -16949 111847 -16915
rect 112126 -16956 112161 -16922
rect 112171 -16956 112172 -16911
rect 112271 -16922 112272 -16911
rect 112282 -16956 112317 -16922
rect 110406 -16985 110869 -16959
rect 110410 -16993 110611 -16985
rect 110426 -17003 110595 -16993
rect 110152 -17140 110327 -17114
rect 109659 -17174 109694 -17140
rect 109755 -17174 109790 -17140
rect 109851 -17174 109886 -17140
rect 109947 -17174 109982 -17140
rect 110043 -17174 110078 -17140
rect 110139 -17174 110327 -17140
rect 110152 -17200 110327 -17174
rect 110352 -17174 110453 -17050
rect 110230 -17870 110265 -17200
rect 110352 -17228 110355 -17174
rect 110037 -17936 110182 -17924
rect 109705 -17970 110182 -17936
rect 110037 -17971 110182 -17970
rect 110218 -17971 110265 -17870
rect 110364 -17971 110399 -17174
rect 110622 -17971 110657 -17062
rect 110756 -17971 110791 -16985
rect 111009 -17002 111044 -16968
rect 111105 -17002 111140 -16968
rect 111201 -17002 111236 -16968
rect 111297 -17002 111332 -16968
rect 111393 -17002 111428 -16968
rect 111489 -17002 111524 -16968
rect 111585 -17002 111620 -16968
rect 112094 -16992 112129 -16958
rect 112166 -16992 112201 -16958
rect 112512 -16995 112547 -16961
rect 112557 -16995 112558 -16950
rect 112699 -17001 112700 -16697
rect 113391 -16706 113426 -16672
rect 113568 -16706 113603 -16672
rect 113864 -16723 113899 -16689
rect 113909 -16723 113910 -16681
rect 114051 -16753 114052 -16525
rect 114741 -16534 114776 -16500
rect 114918 -16534 114953 -16500
rect 115112 -16577 115147 -16543
rect 115157 -16577 115158 -16532
rect 115257 -16543 115258 -16532
rect 115466 -16537 115501 -16503
rect 115511 -16537 115512 -16492
rect 115611 -16503 115612 -16492
rect 115856 -16496 115891 -16462
rect 115901 -16496 115902 -16451
rect 116001 -16462 116002 -16451
rect 116012 -16496 116047 -16462
rect 116057 -16496 116058 -16451
rect 116157 -16462 116158 -16451
rect 116338 -16456 116373 -16422
rect 116410 -16456 116445 -16422
rect 116482 -16456 116517 -16422
rect 116626 -16456 116661 -16422
rect 116698 -16456 116733 -16422
rect 116735 -16456 116805 -16422
rect 116842 -16456 116877 -16422
rect 116912 -16456 116947 -16422
rect 116168 -16496 116203 -16462
rect 117208 -16491 117243 -16457
rect 117253 -16491 117254 -16446
rect 117353 -16457 117354 -16446
rect 117364 -16491 117399 -16457
rect 117409 -16491 117410 -16446
rect 117509 -16457 117510 -16446
rect 118085 -16451 118120 -16417
rect 118262 -16451 118297 -16417
rect 117520 -16491 117555 -16457
rect 115622 -16537 115657 -16503
rect 116901 -16505 116902 -16494
rect 115268 -16577 115303 -16543
rect 114181 -16621 114216 -16587
rect 114382 -16666 114417 -16632
rect 114505 -16637 114506 -16595
rect 114827 -16624 114862 -16590
rect 115466 -16620 115501 -16586
rect 115511 -16620 115512 -16575
rect 115611 -16586 115612 -16575
rect 115856 -16580 115891 -16546
rect 115901 -16580 115902 -16535
rect 116001 -16546 116002 -16535
rect 116012 -16580 116047 -16546
rect 116057 -16580 116058 -16535
rect 116157 -16546 116158 -16535
rect 116735 -16539 116770 -16505
rect 116912 -16539 116947 -16505
rect 116168 -16580 116203 -16546
rect 117055 -16565 117170 -16499
rect 117353 -16525 117354 -16499
rect 117750 -16517 117785 -16483
rect 117795 -16517 117796 -16472
rect 117895 -16483 117896 -16472
rect 117906 -16517 117941 -16483
rect 117951 -16517 117952 -16472
rect 118251 -16500 118252 -16489
rect 118456 -16494 118491 -16460
rect 118501 -16494 118502 -16449
rect 118601 -16460 118602 -16449
rect 118810 -16453 118845 -16419
rect 118855 -16453 118856 -16408
rect 118955 -16419 118956 -16408
rect 119136 -16413 119171 -16379
rect 119200 -16413 119243 -16379
rect 119245 -16413 119246 -16371
rect 119345 -16379 119346 -16371
rect 119280 -16413 119315 -16379
rect 119356 -16413 119391 -16379
rect 119401 -16413 119402 -16371
rect 119501 -16379 119502 -16371
rect 119450 -16413 119485 -16379
rect 119512 -16413 119557 -16379
rect 120552 -16408 120587 -16374
rect 120597 -16408 120598 -16363
rect 120697 -16374 120698 -16363
rect 120708 -16408 120743 -16374
rect 120753 -16408 120754 -16363
rect 120853 -16374 120854 -16363
rect 121429 -16367 121464 -16333
rect 121606 -16367 121641 -16333
rect 122199 -16336 122200 -16328
rect 122299 -16336 122300 -16328
rect 120864 -16408 120899 -16374
rect 118966 -16453 119001 -16419
rect 120245 -16422 120246 -16414
rect 121595 -16417 121596 -16406
rect 121800 -16410 121835 -16376
rect 121845 -16410 121846 -16365
rect 121945 -16376 121946 -16365
rect 122126 -16370 122189 -16336
rect 122198 -16370 122233 -16336
rect 122310 -16370 122345 -16336
rect 123035 -16360 123070 -16326
rect 123131 -16360 123166 -16326
rect 123227 -16360 123262 -16326
rect 123323 -16360 123358 -16326
rect 123419 -16360 123454 -16326
rect 123515 -16360 123550 -16326
rect 123611 -16360 123646 -16326
rect 124939 -16333 124940 -16322
rect 125116 -16327 125179 -16293
rect 125188 -16327 125223 -16293
rect 125300 -16327 125335 -16293
rect 125831 -16317 125866 -16283
rect 125927 -16317 125962 -16283
rect 126023 -16317 126058 -16283
rect 126119 -16317 126154 -16283
rect 126215 -16317 126250 -16283
rect 127240 -16324 127275 -16290
rect 127285 -16324 127286 -16279
rect 127385 -16290 127386 -16279
rect 127396 -16324 127431 -16290
rect 127441 -16324 127442 -16279
rect 127541 -16290 127542 -16279
rect 127720 -16284 127755 -16250
rect 127792 -16284 127827 -16250
rect 127864 -16284 127899 -16250
rect 128008 -16284 128043 -16250
rect 128080 -16284 128115 -16250
rect 128117 -16284 128187 -16250
rect 128224 -16284 128259 -16250
rect 128294 -16284 128329 -16250
rect 128821 -16274 128856 -16240
rect 128917 -16274 128952 -16240
rect 129013 -16274 129048 -16240
rect 130520 -16241 130555 -16207
rect 130584 -16241 130627 -16207
rect 130629 -16241 130630 -16199
rect 130729 -16207 130730 -16199
rect 130664 -16241 130699 -16207
rect 130740 -16241 130775 -16207
rect 130785 -16241 130786 -16199
rect 130885 -16207 130886 -16199
rect 130834 -16241 130869 -16207
rect 130896 -16241 130941 -16207
rect 131811 -16231 131846 -16197
rect 131907 -16231 131942 -16197
rect 132003 -16231 132038 -16197
rect 131627 -16250 131628 -16242
rect 127552 -16324 127587 -16290
rect 128533 -16293 128534 -16285
rect 128633 -16293 128634 -16285
rect 121956 -16410 121991 -16376
rect 118612 -16494 118647 -16460
rect 115622 -16620 115657 -16586
rect 116901 -16589 116902 -16578
rect 114151 -16689 114152 -16681
rect 114162 -16723 114197 -16689
rect 114382 -16734 114417 -16700
rect 112829 -16793 112864 -16759
rect 113032 -16838 113067 -16804
rect 113155 -16809 113156 -16767
rect 113477 -16796 113512 -16762
rect 112799 -16861 112800 -16853
rect 112810 -16895 112845 -16861
rect 113032 -16906 113067 -16872
rect 112799 -16961 112800 -16950
rect 112810 -16995 112845 -16961
rect 111747 -17045 111782 -17011
rect 111843 -17045 111878 -17011
rect 111939 -17045 111974 -17011
rect 112448 -17035 112483 -17001
rect 112520 -17035 112555 -17001
rect 112592 -17035 112627 -17001
rect 112664 -17029 112700 -17001
rect 113010 -17025 113045 -16991
rect 113055 -17025 113056 -16980
rect 112664 -17035 112699 -17029
rect 112101 -17088 112136 -17054
rect 112197 -17088 112232 -17054
rect 112293 -17088 112328 -17054
rect 113197 -17076 113198 -16809
rect 113826 -16819 114213 -16753
rect 113213 -16860 113248 -16826
rect 113562 -16832 113573 -16819
rect 113496 -16874 113573 -16832
rect 113624 -16874 114213 -16819
rect 114360 -16853 114395 -16819
rect 114405 -16853 114406 -16808
rect 113496 -16877 114213 -16874
rect 113213 -16928 113248 -16894
rect 113416 -16942 113451 -16908
rect 113461 -16942 113462 -16900
rect 113297 -16991 113298 -16980
rect 113308 -17025 113343 -16991
rect 113416 -17042 113451 -17008
rect 113461 -17042 113462 -16997
rect 113309 -17078 113344 -17044
rect 113381 -17078 113416 -17044
rect 113453 -17078 113488 -17044
rect 112455 -17131 112490 -17097
rect 112551 -17131 112586 -17097
rect 112647 -17131 112682 -17097
rect 112743 -17131 112778 -17097
rect 112839 -17131 112874 -17097
rect 113496 -17114 113641 -16877
rect 113826 -16899 114213 -16877
rect 113750 -16925 114213 -16899
rect 114547 -16904 114548 -16637
rect 114563 -16688 114598 -16654
rect 115177 -16691 115212 -16657
rect 115856 -16663 115891 -16629
rect 115901 -16663 115902 -16618
rect 116001 -16629 116002 -16618
rect 116012 -16663 116047 -16629
rect 116057 -16663 116058 -16618
rect 116157 -16629 116158 -16618
rect 116735 -16623 116770 -16589
rect 116912 -16623 116947 -16589
rect 117273 -16605 117308 -16571
rect 116168 -16663 116203 -16629
rect 116001 -16697 116002 -16671
rect 116400 -16689 116435 -16655
rect 116445 -16689 116446 -16644
rect 116545 -16655 116546 -16644
rect 116556 -16689 116591 -16655
rect 116601 -16689 116602 -16644
rect 116901 -16672 116902 -16661
rect 114563 -16756 114598 -16722
rect 114766 -16770 114801 -16736
rect 114811 -16770 114812 -16728
rect 114911 -16740 114912 -16729
rect 115531 -16734 115566 -16700
rect 114922 -16774 114957 -16740
rect 114647 -16819 114648 -16808
rect 115116 -16813 115151 -16779
rect 115161 -16813 115162 -16771
rect 115261 -16779 115262 -16771
rect 115921 -16777 115956 -16743
rect 115272 -16813 115307 -16779
rect 114658 -16853 114693 -16819
rect 114766 -16870 114801 -16836
rect 114811 -16870 114812 -16825
rect 114911 -16832 114912 -16821
rect 114922 -16866 114957 -16832
rect 115470 -16856 115505 -16822
rect 115515 -16856 115516 -16814
rect 115615 -16822 115616 -16814
rect 115626 -16856 115661 -16822
rect 114659 -16906 114694 -16872
rect 114731 -16906 114766 -16872
rect 114803 -16906 114838 -16872
rect 115116 -16913 115151 -16879
rect 115161 -16913 115162 -16868
rect 115261 -16879 115262 -16868
rect 115272 -16913 115307 -16879
rect 115856 -16895 115891 -16861
rect 115901 -16895 115902 -16853
rect 113750 -16959 114226 -16925
rect 115084 -16949 115119 -16915
rect 115156 -16949 115191 -16915
rect 115470 -16956 115505 -16922
rect 115515 -16956 115516 -16911
rect 115615 -16922 115616 -16911
rect 115626 -16956 115661 -16922
rect 113750 -16985 114213 -16959
rect 113754 -16993 113955 -16985
rect 113770 -17003 113939 -16993
rect 113496 -17140 113671 -17114
rect 113003 -17174 113038 -17140
rect 113099 -17174 113134 -17140
rect 113195 -17174 113230 -17140
rect 113291 -17174 113326 -17140
rect 113387 -17174 113422 -17140
rect 113483 -17174 113671 -17140
rect 113496 -17200 113671 -17174
rect 113696 -17174 113797 -17050
rect 113574 -17870 113609 -17200
rect 113696 -17228 113699 -17174
rect 113381 -17936 113526 -17924
rect 113049 -17970 113526 -17936
rect 113381 -17971 113526 -17970
rect 113562 -17971 113609 -17870
rect 113708 -17971 113743 -17174
rect 113966 -17971 114001 -17062
rect 114100 -17971 114135 -16985
rect 114353 -17002 114388 -16968
rect 114449 -17002 114484 -16968
rect 114545 -17002 114580 -16968
rect 114641 -17002 114676 -16968
rect 114737 -17002 114772 -16968
rect 114833 -17002 114868 -16968
rect 114929 -17002 114964 -16968
rect 115438 -16992 115473 -16958
rect 115510 -16992 115545 -16958
rect 115856 -16995 115891 -16961
rect 115901 -16995 115902 -16950
rect 116043 -17001 116044 -16697
rect 116735 -16706 116770 -16672
rect 116912 -16706 116947 -16672
rect 117208 -16723 117243 -16689
rect 117253 -16723 117254 -16681
rect 117395 -16753 117396 -16525
rect 118085 -16534 118120 -16500
rect 118262 -16534 118297 -16500
rect 118456 -16577 118491 -16543
rect 118501 -16577 118502 -16532
rect 118601 -16543 118602 -16532
rect 118810 -16537 118845 -16503
rect 118855 -16537 118856 -16492
rect 118955 -16503 118956 -16492
rect 119200 -16496 119235 -16462
rect 119245 -16496 119246 -16451
rect 119345 -16462 119346 -16451
rect 119356 -16496 119391 -16462
rect 119401 -16496 119402 -16451
rect 119501 -16462 119502 -16451
rect 119682 -16456 119717 -16422
rect 119754 -16456 119789 -16422
rect 119826 -16456 119861 -16422
rect 119970 -16456 120005 -16422
rect 120042 -16456 120077 -16422
rect 120079 -16456 120149 -16422
rect 120186 -16456 120221 -16422
rect 120256 -16456 120291 -16422
rect 119512 -16496 119547 -16462
rect 120552 -16491 120587 -16457
rect 120597 -16491 120598 -16446
rect 120697 -16457 120698 -16446
rect 120708 -16491 120743 -16457
rect 120753 -16491 120754 -16446
rect 120853 -16457 120854 -16446
rect 121429 -16451 121464 -16417
rect 121606 -16451 121641 -16417
rect 120864 -16491 120899 -16457
rect 118966 -16537 119001 -16503
rect 120245 -16505 120246 -16494
rect 118612 -16577 118647 -16543
rect 117525 -16621 117560 -16587
rect 117726 -16666 117761 -16632
rect 117849 -16637 117850 -16595
rect 118171 -16624 118206 -16590
rect 118810 -16620 118845 -16586
rect 118855 -16620 118856 -16575
rect 118955 -16586 118956 -16575
rect 119200 -16580 119235 -16546
rect 119245 -16580 119246 -16535
rect 119345 -16546 119346 -16535
rect 119356 -16580 119391 -16546
rect 119401 -16580 119402 -16535
rect 119501 -16546 119502 -16535
rect 120079 -16539 120114 -16505
rect 120256 -16539 120291 -16505
rect 119512 -16580 119547 -16546
rect 120399 -16565 120514 -16499
rect 120697 -16525 120698 -16499
rect 121094 -16517 121129 -16483
rect 121139 -16517 121140 -16472
rect 121239 -16483 121240 -16472
rect 121250 -16517 121285 -16483
rect 121295 -16517 121296 -16472
rect 121595 -16500 121596 -16489
rect 121800 -16494 121835 -16460
rect 121845 -16494 121846 -16449
rect 121945 -16460 121946 -16449
rect 122154 -16453 122189 -16419
rect 122199 -16453 122200 -16408
rect 122299 -16419 122300 -16408
rect 122480 -16413 122515 -16379
rect 122544 -16413 122587 -16379
rect 122589 -16413 122590 -16371
rect 122689 -16379 122690 -16371
rect 122624 -16413 122659 -16379
rect 122700 -16413 122735 -16379
rect 122745 -16413 122746 -16371
rect 122845 -16379 122846 -16371
rect 122794 -16413 122829 -16379
rect 122856 -16413 122901 -16379
rect 123896 -16408 123931 -16374
rect 123941 -16408 123942 -16363
rect 124041 -16374 124042 -16363
rect 124052 -16408 124087 -16374
rect 124097 -16408 124098 -16363
rect 124197 -16374 124198 -16363
rect 124773 -16367 124808 -16333
rect 124950 -16367 124985 -16333
rect 125543 -16336 125544 -16328
rect 125643 -16336 125644 -16328
rect 124208 -16408 124243 -16374
rect 122310 -16453 122345 -16419
rect 123589 -16422 123590 -16414
rect 124939 -16417 124940 -16406
rect 125144 -16410 125179 -16376
rect 125189 -16410 125190 -16365
rect 125289 -16376 125290 -16365
rect 125470 -16370 125533 -16336
rect 125542 -16370 125577 -16336
rect 125654 -16370 125689 -16336
rect 126379 -16360 126414 -16326
rect 126475 -16360 126510 -16326
rect 126571 -16360 126606 -16326
rect 126667 -16360 126702 -16326
rect 126763 -16360 126798 -16326
rect 126859 -16360 126894 -16326
rect 126955 -16360 126990 -16326
rect 128283 -16333 128284 -16322
rect 128460 -16327 128523 -16293
rect 128532 -16327 128567 -16293
rect 128644 -16327 128679 -16293
rect 129175 -16317 129210 -16283
rect 129271 -16317 129306 -16283
rect 129367 -16317 129402 -16283
rect 129463 -16317 129498 -16283
rect 129559 -16317 129594 -16283
rect 130584 -16324 130619 -16290
rect 130629 -16324 130630 -16279
rect 130729 -16290 130730 -16279
rect 130740 -16324 130775 -16290
rect 130785 -16324 130786 -16279
rect 130885 -16290 130886 -16279
rect 131064 -16284 131099 -16250
rect 131136 -16284 131171 -16250
rect 131208 -16284 131243 -16250
rect 131352 -16284 131387 -16250
rect 131424 -16284 131459 -16250
rect 131461 -16284 131531 -16250
rect 131568 -16284 131603 -16250
rect 131638 -16284 131673 -16250
rect 132165 -16274 132200 -16240
rect 132261 -16274 132296 -16240
rect 132357 -16274 132392 -16240
rect 133864 -16241 133899 -16207
rect 133928 -16241 133971 -16207
rect 133973 -16241 133974 -16199
rect 134073 -16207 134074 -16199
rect 134008 -16241 134043 -16207
rect 134084 -16241 134119 -16207
rect 134129 -16241 134130 -16199
rect 134229 -16207 134230 -16199
rect 134178 -16241 134213 -16207
rect 134240 -16241 134285 -16207
rect 135155 -16231 135190 -16197
rect 135251 -16231 135286 -16197
rect 135347 -16231 135382 -16197
rect 134971 -16250 134972 -16242
rect 130896 -16324 130931 -16290
rect 131877 -16293 131878 -16285
rect 131977 -16293 131978 -16285
rect 125300 -16410 125335 -16376
rect 121956 -16494 121991 -16460
rect 118966 -16620 119001 -16586
rect 120245 -16589 120246 -16578
rect 117495 -16689 117496 -16681
rect 117506 -16723 117541 -16689
rect 117726 -16734 117761 -16700
rect 116173 -16793 116208 -16759
rect 116376 -16838 116411 -16804
rect 116499 -16809 116500 -16767
rect 116821 -16796 116856 -16762
rect 116143 -16861 116144 -16853
rect 116154 -16895 116189 -16861
rect 116376 -16906 116411 -16872
rect 116143 -16961 116144 -16950
rect 116154 -16995 116189 -16961
rect 115091 -17045 115126 -17011
rect 115187 -17045 115222 -17011
rect 115283 -17045 115318 -17011
rect 115792 -17035 115827 -17001
rect 115864 -17035 115899 -17001
rect 115936 -17035 115971 -17001
rect 116008 -17029 116044 -17001
rect 116354 -17025 116389 -16991
rect 116399 -17025 116400 -16980
rect 116008 -17035 116043 -17029
rect 115445 -17088 115480 -17054
rect 115541 -17088 115576 -17054
rect 115637 -17088 115672 -17054
rect 116541 -17076 116542 -16809
rect 117170 -16819 117557 -16753
rect 116557 -16860 116592 -16826
rect 116906 -16832 116917 -16819
rect 116840 -16874 116917 -16832
rect 116968 -16874 117557 -16819
rect 117704 -16853 117739 -16819
rect 117749 -16853 117750 -16808
rect 116840 -16877 117557 -16874
rect 116557 -16928 116592 -16894
rect 116760 -16942 116795 -16908
rect 116805 -16942 116806 -16900
rect 116641 -16991 116642 -16980
rect 116652 -17025 116687 -16991
rect 116760 -17042 116795 -17008
rect 116805 -17042 116806 -16997
rect 116653 -17078 116688 -17044
rect 116725 -17078 116760 -17044
rect 116797 -17078 116832 -17044
rect 115799 -17131 115834 -17097
rect 115895 -17131 115930 -17097
rect 115991 -17131 116026 -17097
rect 116087 -17131 116122 -17097
rect 116183 -17131 116218 -17097
rect 116840 -17114 116985 -16877
rect 117170 -16899 117557 -16877
rect 117094 -16925 117557 -16899
rect 117891 -16904 117892 -16637
rect 117907 -16688 117942 -16654
rect 118521 -16691 118556 -16657
rect 119200 -16663 119235 -16629
rect 119245 -16663 119246 -16618
rect 119345 -16629 119346 -16618
rect 119356 -16663 119391 -16629
rect 119401 -16663 119402 -16618
rect 119501 -16629 119502 -16618
rect 120079 -16623 120114 -16589
rect 120256 -16623 120291 -16589
rect 120617 -16605 120652 -16571
rect 119512 -16663 119547 -16629
rect 119345 -16697 119346 -16671
rect 119744 -16689 119779 -16655
rect 119789 -16689 119790 -16644
rect 119889 -16655 119890 -16644
rect 119900 -16689 119935 -16655
rect 119945 -16689 119946 -16644
rect 120245 -16672 120246 -16661
rect 117907 -16756 117942 -16722
rect 118110 -16770 118145 -16736
rect 118155 -16770 118156 -16728
rect 118255 -16740 118256 -16729
rect 118875 -16734 118910 -16700
rect 118266 -16774 118301 -16740
rect 117991 -16819 117992 -16808
rect 118460 -16813 118495 -16779
rect 118505 -16813 118506 -16771
rect 118605 -16779 118606 -16771
rect 119265 -16777 119300 -16743
rect 118616 -16813 118651 -16779
rect 118002 -16853 118037 -16819
rect 118110 -16870 118145 -16836
rect 118155 -16870 118156 -16825
rect 118255 -16832 118256 -16821
rect 118266 -16866 118301 -16832
rect 118814 -16856 118849 -16822
rect 118859 -16856 118860 -16814
rect 118959 -16822 118960 -16814
rect 118970 -16856 119005 -16822
rect 118003 -16906 118038 -16872
rect 118075 -16906 118110 -16872
rect 118147 -16906 118182 -16872
rect 118460 -16913 118495 -16879
rect 118505 -16913 118506 -16868
rect 118605 -16879 118606 -16868
rect 118616 -16913 118651 -16879
rect 119200 -16895 119235 -16861
rect 119245 -16895 119246 -16853
rect 117094 -16959 117570 -16925
rect 118428 -16949 118463 -16915
rect 118500 -16949 118535 -16915
rect 118814 -16956 118849 -16922
rect 118859 -16956 118860 -16911
rect 118959 -16922 118960 -16911
rect 118970 -16956 119005 -16922
rect 117094 -16985 117557 -16959
rect 117098 -16993 117299 -16985
rect 117114 -17003 117283 -16993
rect 116840 -17140 117015 -17114
rect 116347 -17174 116382 -17140
rect 116443 -17174 116478 -17140
rect 116539 -17174 116574 -17140
rect 116635 -17174 116670 -17140
rect 116731 -17174 116766 -17140
rect 116827 -17174 117015 -17140
rect 116840 -17200 117015 -17174
rect 117040 -17174 117141 -17050
rect 116918 -17870 116953 -17200
rect 117040 -17228 117043 -17174
rect 116725 -17936 116870 -17924
rect 116393 -17970 116870 -17936
rect 116725 -17971 116870 -17970
rect 116906 -17971 116953 -17870
rect 117052 -17971 117087 -17174
rect 117310 -17971 117345 -17062
rect 117444 -17971 117479 -16985
rect 117697 -17002 117732 -16968
rect 117793 -17002 117828 -16968
rect 117889 -17002 117924 -16968
rect 117985 -17002 118020 -16968
rect 118081 -17002 118116 -16968
rect 118177 -17002 118212 -16968
rect 118273 -17002 118308 -16968
rect 118782 -16992 118817 -16958
rect 118854 -16992 118889 -16958
rect 119200 -16995 119235 -16961
rect 119245 -16995 119246 -16950
rect 119387 -17001 119388 -16697
rect 120079 -16706 120114 -16672
rect 120256 -16706 120291 -16672
rect 120552 -16723 120587 -16689
rect 120597 -16723 120598 -16681
rect 120739 -16753 120740 -16525
rect 121429 -16534 121464 -16500
rect 121606 -16534 121641 -16500
rect 121800 -16577 121835 -16543
rect 121845 -16577 121846 -16532
rect 121945 -16543 121946 -16532
rect 122154 -16537 122189 -16503
rect 122199 -16537 122200 -16492
rect 122299 -16503 122300 -16492
rect 122544 -16496 122579 -16462
rect 122589 -16496 122590 -16451
rect 122689 -16462 122690 -16451
rect 122700 -16496 122735 -16462
rect 122745 -16496 122746 -16451
rect 122845 -16462 122846 -16451
rect 123026 -16456 123061 -16422
rect 123098 -16456 123133 -16422
rect 123170 -16456 123205 -16422
rect 123314 -16456 123349 -16422
rect 123386 -16456 123421 -16422
rect 123423 -16456 123493 -16422
rect 123530 -16456 123565 -16422
rect 123600 -16456 123635 -16422
rect 122856 -16496 122891 -16462
rect 123896 -16491 123931 -16457
rect 123941 -16491 123942 -16446
rect 124041 -16457 124042 -16446
rect 124052 -16491 124087 -16457
rect 124097 -16491 124098 -16446
rect 124197 -16457 124198 -16446
rect 124773 -16451 124808 -16417
rect 124950 -16451 124985 -16417
rect 124208 -16491 124243 -16457
rect 122310 -16537 122345 -16503
rect 123589 -16505 123590 -16494
rect 121956 -16577 121991 -16543
rect 120869 -16621 120904 -16587
rect 121070 -16666 121105 -16632
rect 121193 -16637 121194 -16595
rect 121515 -16624 121550 -16590
rect 122154 -16620 122189 -16586
rect 122199 -16620 122200 -16575
rect 122299 -16586 122300 -16575
rect 122544 -16580 122579 -16546
rect 122589 -16580 122590 -16535
rect 122689 -16546 122690 -16535
rect 122700 -16580 122735 -16546
rect 122745 -16580 122746 -16535
rect 122845 -16546 122846 -16535
rect 123423 -16539 123458 -16505
rect 123600 -16539 123635 -16505
rect 122856 -16580 122891 -16546
rect 123743 -16565 123858 -16499
rect 124041 -16525 124042 -16499
rect 124438 -16517 124473 -16483
rect 124483 -16517 124484 -16472
rect 124583 -16483 124584 -16472
rect 124594 -16517 124629 -16483
rect 124639 -16517 124640 -16472
rect 124939 -16500 124940 -16489
rect 125144 -16494 125179 -16460
rect 125189 -16494 125190 -16449
rect 125289 -16460 125290 -16449
rect 125498 -16453 125533 -16419
rect 125543 -16453 125544 -16408
rect 125643 -16419 125644 -16408
rect 125824 -16413 125859 -16379
rect 125888 -16413 125931 -16379
rect 125933 -16413 125934 -16371
rect 126033 -16379 126034 -16371
rect 125968 -16413 126003 -16379
rect 126044 -16413 126079 -16379
rect 126089 -16413 126090 -16371
rect 126189 -16379 126190 -16371
rect 126138 -16413 126173 -16379
rect 126200 -16413 126245 -16379
rect 127240 -16408 127275 -16374
rect 127285 -16408 127286 -16363
rect 127385 -16374 127386 -16363
rect 127396 -16408 127431 -16374
rect 127441 -16408 127442 -16363
rect 127541 -16374 127542 -16363
rect 128117 -16367 128152 -16333
rect 128294 -16367 128329 -16333
rect 128887 -16336 128888 -16328
rect 128987 -16336 128988 -16328
rect 127552 -16408 127587 -16374
rect 125654 -16453 125689 -16419
rect 126933 -16422 126934 -16414
rect 128283 -16417 128284 -16406
rect 128488 -16410 128523 -16376
rect 128533 -16410 128534 -16365
rect 128633 -16376 128634 -16365
rect 128814 -16370 128877 -16336
rect 128886 -16370 128921 -16336
rect 128998 -16370 129033 -16336
rect 129723 -16360 129758 -16326
rect 129819 -16360 129854 -16326
rect 129915 -16360 129950 -16326
rect 130011 -16360 130046 -16326
rect 130107 -16360 130142 -16326
rect 130203 -16360 130238 -16326
rect 130299 -16360 130334 -16326
rect 131627 -16333 131628 -16322
rect 131804 -16327 131867 -16293
rect 131876 -16327 131911 -16293
rect 131988 -16327 132023 -16293
rect 132519 -16317 132554 -16283
rect 132615 -16317 132650 -16283
rect 132711 -16317 132746 -16283
rect 132807 -16317 132842 -16283
rect 132903 -16317 132938 -16283
rect 133928 -16324 133963 -16290
rect 133973 -16324 133974 -16279
rect 134073 -16290 134074 -16279
rect 134084 -16324 134119 -16290
rect 134129 -16324 134130 -16279
rect 134229 -16290 134230 -16279
rect 134408 -16284 134443 -16250
rect 134480 -16284 134515 -16250
rect 134552 -16284 134587 -16250
rect 134696 -16284 134731 -16250
rect 134768 -16284 134803 -16250
rect 134805 -16284 134875 -16250
rect 134912 -16284 134947 -16250
rect 134982 -16284 135017 -16250
rect 135509 -16274 135544 -16240
rect 135605 -16274 135640 -16240
rect 135701 -16274 135736 -16240
rect 137208 -16241 137243 -16207
rect 137272 -16241 137315 -16207
rect 137317 -16241 137318 -16199
rect 137417 -16207 137418 -16199
rect 137352 -16241 137387 -16207
rect 137428 -16241 137463 -16207
rect 137473 -16241 137474 -16199
rect 137573 -16207 137574 -16199
rect 137522 -16241 137557 -16207
rect 137584 -16241 137629 -16207
rect 138499 -16231 138534 -16197
rect 138595 -16231 138630 -16197
rect 138691 -16231 138726 -16197
rect 138315 -16250 138316 -16242
rect 134240 -16324 134275 -16290
rect 135221 -16293 135222 -16285
rect 135321 -16293 135322 -16285
rect 128644 -16410 128679 -16376
rect 125300 -16494 125335 -16460
rect 122310 -16620 122345 -16586
rect 123589 -16589 123590 -16578
rect 120839 -16689 120840 -16681
rect 120850 -16723 120885 -16689
rect 121070 -16734 121105 -16700
rect 119517 -16793 119552 -16759
rect 119720 -16838 119755 -16804
rect 119843 -16809 119844 -16767
rect 120165 -16796 120200 -16762
rect 119487 -16861 119488 -16853
rect 119498 -16895 119533 -16861
rect 119720 -16906 119755 -16872
rect 119487 -16961 119488 -16950
rect 119498 -16995 119533 -16961
rect 118435 -17045 118470 -17011
rect 118531 -17045 118566 -17011
rect 118627 -17045 118662 -17011
rect 119136 -17035 119171 -17001
rect 119208 -17035 119243 -17001
rect 119280 -17035 119315 -17001
rect 119352 -17029 119388 -17001
rect 119698 -17025 119733 -16991
rect 119743 -17025 119744 -16980
rect 119352 -17035 119387 -17029
rect 118789 -17088 118824 -17054
rect 118885 -17088 118920 -17054
rect 118981 -17088 119016 -17054
rect 119885 -17076 119886 -16809
rect 120514 -16819 120901 -16753
rect 119901 -16860 119936 -16826
rect 120250 -16832 120261 -16819
rect 120184 -16874 120261 -16832
rect 120312 -16874 120901 -16819
rect 121048 -16853 121083 -16819
rect 121093 -16853 121094 -16808
rect 120184 -16877 120901 -16874
rect 119901 -16928 119936 -16894
rect 120104 -16942 120139 -16908
rect 120149 -16942 120150 -16900
rect 119985 -16991 119986 -16980
rect 119996 -17025 120031 -16991
rect 120104 -17042 120139 -17008
rect 120149 -17042 120150 -16997
rect 119997 -17078 120032 -17044
rect 120069 -17078 120104 -17044
rect 120141 -17078 120176 -17044
rect 119143 -17131 119178 -17097
rect 119239 -17131 119274 -17097
rect 119335 -17131 119370 -17097
rect 119431 -17131 119466 -17097
rect 119527 -17131 119562 -17097
rect 120184 -17114 120329 -16877
rect 120514 -16899 120901 -16877
rect 120438 -16925 120901 -16899
rect 121235 -16904 121236 -16637
rect 121251 -16688 121286 -16654
rect 121865 -16691 121900 -16657
rect 122544 -16663 122579 -16629
rect 122589 -16663 122590 -16618
rect 122689 -16629 122690 -16618
rect 122700 -16663 122735 -16629
rect 122745 -16663 122746 -16618
rect 122845 -16629 122846 -16618
rect 123423 -16623 123458 -16589
rect 123600 -16623 123635 -16589
rect 123961 -16605 123996 -16571
rect 122856 -16663 122891 -16629
rect 122689 -16697 122690 -16671
rect 123088 -16689 123123 -16655
rect 123133 -16689 123134 -16644
rect 123233 -16655 123234 -16644
rect 123244 -16689 123279 -16655
rect 123289 -16689 123290 -16644
rect 123589 -16672 123590 -16661
rect 121251 -16756 121286 -16722
rect 121454 -16770 121489 -16736
rect 121499 -16770 121500 -16728
rect 121599 -16740 121600 -16729
rect 122219 -16734 122254 -16700
rect 121610 -16774 121645 -16740
rect 121335 -16819 121336 -16808
rect 121804 -16813 121839 -16779
rect 121849 -16813 121850 -16771
rect 121949 -16779 121950 -16771
rect 122609 -16777 122644 -16743
rect 121960 -16813 121995 -16779
rect 121346 -16853 121381 -16819
rect 121454 -16870 121489 -16836
rect 121499 -16870 121500 -16825
rect 121599 -16832 121600 -16821
rect 121610 -16866 121645 -16832
rect 122158 -16856 122193 -16822
rect 122203 -16856 122204 -16814
rect 122303 -16822 122304 -16814
rect 122314 -16856 122349 -16822
rect 121347 -16906 121382 -16872
rect 121419 -16906 121454 -16872
rect 121491 -16906 121526 -16872
rect 121804 -16913 121839 -16879
rect 121849 -16913 121850 -16868
rect 121949 -16879 121950 -16868
rect 121960 -16913 121995 -16879
rect 122544 -16895 122579 -16861
rect 122589 -16895 122590 -16853
rect 120438 -16959 120914 -16925
rect 121772 -16949 121807 -16915
rect 121844 -16949 121879 -16915
rect 122158 -16956 122193 -16922
rect 122203 -16956 122204 -16911
rect 122303 -16922 122304 -16911
rect 122314 -16956 122349 -16922
rect 120438 -16985 120901 -16959
rect 120442 -16993 120643 -16985
rect 120458 -17003 120627 -16993
rect 120184 -17140 120359 -17114
rect 119691 -17174 119726 -17140
rect 119787 -17174 119822 -17140
rect 119883 -17174 119918 -17140
rect 119979 -17174 120014 -17140
rect 120075 -17174 120110 -17140
rect 120171 -17174 120359 -17140
rect 120184 -17200 120359 -17174
rect 120384 -17174 120485 -17050
rect 120262 -17870 120297 -17200
rect 120384 -17228 120387 -17174
rect 120069 -17936 120214 -17924
rect 119737 -17970 120214 -17936
rect 120069 -17971 120214 -17970
rect 120250 -17971 120297 -17870
rect 120396 -17971 120431 -17174
rect 120654 -17971 120689 -17062
rect 120788 -17971 120823 -16985
rect 121041 -17002 121076 -16968
rect 121137 -17002 121172 -16968
rect 121233 -17002 121268 -16968
rect 121329 -17002 121364 -16968
rect 121425 -17002 121460 -16968
rect 121521 -17002 121556 -16968
rect 121617 -17002 121652 -16968
rect 122126 -16992 122161 -16958
rect 122198 -16992 122233 -16958
rect 122544 -16995 122579 -16961
rect 122589 -16995 122590 -16950
rect 122731 -17001 122732 -16697
rect 123423 -16706 123458 -16672
rect 123600 -16706 123635 -16672
rect 123896 -16723 123931 -16689
rect 123941 -16723 123942 -16681
rect 124083 -16753 124084 -16525
rect 124773 -16534 124808 -16500
rect 124950 -16534 124985 -16500
rect 125144 -16577 125179 -16543
rect 125189 -16577 125190 -16532
rect 125289 -16543 125290 -16532
rect 125498 -16537 125533 -16503
rect 125543 -16537 125544 -16492
rect 125643 -16503 125644 -16492
rect 125888 -16496 125923 -16462
rect 125933 -16496 125934 -16451
rect 126033 -16462 126034 -16451
rect 126044 -16496 126079 -16462
rect 126089 -16496 126090 -16451
rect 126189 -16462 126190 -16451
rect 126370 -16456 126405 -16422
rect 126442 -16456 126477 -16422
rect 126514 -16456 126549 -16422
rect 126658 -16456 126693 -16422
rect 126730 -16456 126765 -16422
rect 126767 -16456 126837 -16422
rect 126874 -16456 126909 -16422
rect 126944 -16456 126979 -16422
rect 126200 -16496 126235 -16462
rect 127240 -16491 127275 -16457
rect 127285 -16491 127286 -16446
rect 127385 -16457 127386 -16446
rect 127396 -16491 127431 -16457
rect 127441 -16491 127442 -16446
rect 127541 -16457 127542 -16446
rect 128117 -16451 128152 -16417
rect 128294 -16451 128329 -16417
rect 127552 -16491 127587 -16457
rect 125654 -16537 125689 -16503
rect 126933 -16505 126934 -16494
rect 125300 -16577 125335 -16543
rect 124213 -16621 124248 -16587
rect 124414 -16666 124449 -16632
rect 124537 -16637 124538 -16595
rect 124859 -16624 124894 -16590
rect 125498 -16620 125533 -16586
rect 125543 -16620 125544 -16575
rect 125643 -16586 125644 -16575
rect 125888 -16580 125923 -16546
rect 125933 -16580 125934 -16535
rect 126033 -16546 126034 -16535
rect 126044 -16580 126079 -16546
rect 126089 -16580 126090 -16535
rect 126189 -16546 126190 -16535
rect 126767 -16539 126802 -16505
rect 126944 -16539 126979 -16505
rect 126200 -16580 126235 -16546
rect 127087 -16565 127202 -16499
rect 127385 -16525 127386 -16499
rect 127782 -16517 127817 -16483
rect 127827 -16517 127828 -16472
rect 127927 -16483 127928 -16472
rect 127938 -16517 127973 -16483
rect 127983 -16517 127984 -16472
rect 128283 -16500 128284 -16489
rect 128488 -16494 128523 -16460
rect 128533 -16494 128534 -16449
rect 128633 -16460 128634 -16449
rect 128842 -16453 128877 -16419
rect 128887 -16453 128888 -16408
rect 128987 -16419 128988 -16408
rect 129168 -16413 129203 -16379
rect 129232 -16413 129275 -16379
rect 129277 -16413 129278 -16371
rect 129377 -16379 129378 -16371
rect 129312 -16413 129347 -16379
rect 129388 -16413 129423 -16379
rect 129433 -16413 129434 -16371
rect 129533 -16379 129534 -16371
rect 129482 -16413 129517 -16379
rect 129544 -16413 129589 -16379
rect 130584 -16408 130619 -16374
rect 130629 -16408 130630 -16363
rect 130729 -16374 130730 -16363
rect 130740 -16408 130775 -16374
rect 130785 -16408 130786 -16363
rect 130885 -16374 130886 -16363
rect 131461 -16367 131496 -16333
rect 131638 -16367 131673 -16333
rect 132231 -16336 132232 -16328
rect 132331 -16336 132332 -16328
rect 130896 -16408 130931 -16374
rect 128998 -16453 129033 -16419
rect 130277 -16422 130278 -16414
rect 131627 -16417 131628 -16406
rect 131832 -16410 131867 -16376
rect 131877 -16410 131878 -16365
rect 131977 -16376 131978 -16365
rect 132158 -16370 132221 -16336
rect 132230 -16370 132265 -16336
rect 132342 -16370 132377 -16336
rect 133067 -16360 133102 -16326
rect 133163 -16360 133198 -16326
rect 133259 -16360 133294 -16326
rect 133355 -16360 133390 -16326
rect 133451 -16360 133486 -16326
rect 133547 -16360 133582 -16326
rect 133643 -16360 133678 -16326
rect 134971 -16333 134972 -16322
rect 135148 -16327 135211 -16293
rect 135220 -16327 135255 -16293
rect 135332 -16327 135367 -16293
rect 135863 -16317 135898 -16283
rect 135959 -16317 135994 -16283
rect 136055 -16317 136090 -16283
rect 136151 -16317 136186 -16283
rect 136247 -16317 136282 -16283
rect 137272 -16324 137307 -16290
rect 137317 -16324 137318 -16279
rect 137417 -16290 137418 -16279
rect 137428 -16324 137463 -16290
rect 137473 -16324 137474 -16279
rect 137573 -16290 137574 -16279
rect 137752 -16284 137787 -16250
rect 137824 -16284 137859 -16250
rect 137896 -16284 137931 -16250
rect 138040 -16284 138075 -16250
rect 138112 -16284 138147 -16250
rect 138149 -16284 138219 -16250
rect 138256 -16284 138291 -16250
rect 138326 -16284 138361 -16250
rect 138853 -16274 138888 -16240
rect 138949 -16274 138984 -16240
rect 139045 -16274 139080 -16240
rect 140552 -16241 140587 -16207
rect 140616 -16241 140659 -16207
rect 140661 -16241 140662 -16199
rect 140761 -16207 140762 -16199
rect 140696 -16241 140731 -16207
rect 140772 -16241 140807 -16207
rect 140817 -16241 140818 -16199
rect 140917 -16207 140918 -16199
rect 140866 -16241 140901 -16207
rect 140928 -16241 140973 -16207
rect 141843 -16231 141878 -16197
rect 141939 -16231 141974 -16197
rect 142035 -16231 142070 -16197
rect 141659 -16250 141660 -16242
rect 137584 -16324 137619 -16290
rect 138565 -16293 138566 -16285
rect 138665 -16293 138666 -16285
rect 131988 -16410 132023 -16376
rect 128644 -16494 128679 -16460
rect 125654 -16620 125689 -16586
rect 126933 -16589 126934 -16578
rect 124183 -16689 124184 -16681
rect 124194 -16723 124229 -16689
rect 124414 -16734 124449 -16700
rect 122861 -16793 122896 -16759
rect 123064 -16838 123099 -16804
rect 123187 -16809 123188 -16767
rect 123509 -16796 123544 -16762
rect 122831 -16861 122832 -16853
rect 122842 -16895 122877 -16861
rect 123064 -16906 123099 -16872
rect 122831 -16961 122832 -16950
rect 122842 -16995 122877 -16961
rect 121779 -17045 121814 -17011
rect 121875 -17045 121910 -17011
rect 121971 -17045 122006 -17011
rect 122480 -17035 122515 -17001
rect 122552 -17035 122587 -17001
rect 122624 -17035 122659 -17001
rect 122696 -17029 122732 -17001
rect 123042 -17025 123077 -16991
rect 123087 -17025 123088 -16980
rect 122696 -17035 122731 -17029
rect 122133 -17088 122168 -17054
rect 122229 -17088 122264 -17054
rect 122325 -17088 122360 -17054
rect 123229 -17076 123230 -16809
rect 123858 -16819 124245 -16753
rect 123245 -16860 123280 -16826
rect 123594 -16832 123605 -16819
rect 123528 -16874 123605 -16832
rect 123656 -16874 124245 -16819
rect 124392 -16853 124427 -16819
rect 124437 -16853 124438 -16808
rect 123528 -16877 124245 -16874
rect 123245 -16928 123280 -16894
rect 123448 -16942 123483 -16908
rect 123493 -16942 123494 -16900
rect 123329 -16991 123330 -16980
rect 123340 -17025 123375 -16991
rect 123448 -17042 123483 -17008
rect 123493 -17042 123494 -16997
rect 123341 -17078 123376 -17044
rect 123413 -17078 123448 -17044
rect 123485 -17078 123520 -17044
rect 122487 -17131 122522 -17097
rect 122583 -17131 122618 -17097
rect 122679 -17131 122714 -17097
rect 122775 -17131 122810 -17097
rect 122871 -17131 122906 -17097
rect 123528 -17114 123673 -16877
rect 123858 -16899 124245 -16877
rect 123782 -16925 124245 -16899
rect 124579 -16904 124580 -16637
rect 124595 -16688 124630 -16654
rect 125209 -16691 125244 -16657
rect 125888 -16663 125923 -16629
rect 125933 -16663 125934 -16618
rect 126033 -16629 126034 -16618
rect 126044 -16663 126079 -16629
rect 126089 -16663 126090 -16618
rect 126189 -16629 126190 -16618
rect 126767 -16623 126802 -16589
rect 126944 -16623 126979 -16589
rect 127305 -16605 127340 -16571
rect 126200 -16663 126235 -16629
rect 126033 -16697 126034 -16671
rect 126432 -16689 126467 -16655
rect 126477 -16689 126478 -16644
rect 126577 -16655 126578 -16644
rect 126588 -16689 126623 -16655
rect 126633 -16689 126634 -16644
rect 126933 -16672 126934 -16661
rect 124595 -16756 124630 -16722
rect 124798 -16770 124833 -16736
rect 124843 -16770 124844 -16728
rect 124943 -16740 124944 -16729
rect 125563 -16734 125598 -16700
rect 124954 -16774 124989 -16740
rect 124679 -16819 124680 -16808
rect 125148 -16813 125183 -16779
rect 125193 -16813 125194 -16771
rect 125293 -16779 125294 -16771
rect 125953 -16777 125988 -16743
rect 125304 -16813 125339 -16779
rect 124690 -16853 124725 -16819
rect 124798 -16870 124833 -16836
rect 124843 -16870 124844 -16825
rect 124943 -16832 124944 -16821
rect 124954 -16866 124989 -16832
rect 125502 -16856 125537 -16822
rect 125547 -16856 125548 -16814
rect 125647 -16822 125648 -16814
rect 125658 -16856 125693 -16822
rect 124691 -16906 124726 -16872
rect 124763 -16906 124798 -16872
rect 124835 -16906 124870 -16872
rect 125148 -16913 125183 -16879
rect 125193 -16913 125194 -16868
rect 125293 -16879 125294 -16868
rect 125304 -16913 125339 -16879
rect 125888 -16895 125923 -16861
rect 125933 -16895 125934 -16853
rect 123782 -16959 124258 -16925
rect 125116 -16949 125151 -16915
rect 125188 -16949 125223 -16915
rect 125502 -16956 125537 -16922
rect 125547 -16956 125548 -16911
rect 125647 -16922 125648 -16911
rect 125658 -16956 125693 -16922
rect 123782 -16985 124245 -16959
rect 123786 -16993 123987 -16985
rect 123802 -17003 123971 -16993
rect 123528 -17140 123703 -17114
rect 123035 -17174 123070 -17140
rect 123131 -17174 123166 -17140
rect 123227 -17174 123262 -17140
rect 123323 -17174 123358 -17140
rect 123419 -17174 123454 -17140
rect 123515 -17174 123703 -17140
rect 123528 -17200 123703 -17174
rect 123728 -17174 123829 -17050
rect 123606 -17870 123641 -17200
rect 123728 -17228 123731 -17174
rect 123413 -17936 123558 -17924
rect 123081 -17970 123558 -17936
rect 123413 -17971 123558 -17970
rect 123594 -17971 123641 -17870
rect 123740 -17971 123775 -17174
rect 123998 -17971 124033 -17062
rect 124132 -17971 124167 -16985
rect 124385 -17002 124420 -16968
rect 124481 -17002 124516 -16968
rect 124577 -17002 124612 -16968
rect 124673 -17002 124708 -16968
rect 124769 -17002 124804 -16968
rect 124865 -17002 124900 -16968
rect 124961 -17002 124996 -16968
rect 125470 -16992 125505 -16958
rect 125542 -16992 125577 -16958
rect 125888 -16995 125923 -16961
rect 125933 -16995 125934 -16950
rect 126075 -17001 126076 -16697
rect 126767 -16706 126802 -16672
rect 126944 -16706 126979 -16672
rect 127240 -16723 127275 -16689
rect 127285 -16723 127286 -16681
rect 127427 -16753 127428 -16525
rect 128117 -16534 128152 -16500
rect 128294 -16534 128329 -16500
rect 128488 -16577 128523 -16543
rect 128533 -16577 128534 -16532
rect 128633 -16543 128634 -16532
rect 128842 -16537 128877 -16503
rect 128887 -16537 128888 -16492
rect 128987 -16503 128988 -16492
rect 129232 -16496 129267 -16462
rect 129277 -16496 129278 -16451
rect 129377 -16462 129378 -16451
rect 129388 -16496 129423 -16462
rect 129433 -16496 129434 -16451
rect 129533 -16462 129534 -16451
rect 129714 -16456 129749 -16422
rect 129786 -16456 129821 -16422
rect 129858 -16456 129893 -16422
rect 130002 -16456 130037 -16422
rect 130074 -16456 130109 -16422
rect 130111 -16456 130181 -16422
rect 130218 -16456 130253 -16422
rect 130288 -16456 130323 -16422
rect 129544 -16496 129579 -16462
rect 130584 -16491 130619 -16457
rect 130629 -16491 130630 -16446
rect 130729 -16457 130730 -16446
rect 130740 -16491 130775 -16457
rect 130785 -16491 130786 -16446
rect 130885 -16457 130886 -16446
rect 131461 -16451 131496 -16417
rect 131638 -16451 131673 -16417
rect 130896 -16491 130931 -16457
rect 128998 -16537 129033 -16503
rect 130277 -16505 130278 -16494
rect 128644 -16577 128679 -16543
rect 127557 -16621 127592 -16587
rect 127758 -16666 127793 -16632
rect 127881 -16637 127882 -16595
rect 128203 -16624 128238 -16590
rect 128842 -16620 128877 -16586
rect 128887 -16620 128888 -16575
rect 128987 -16586 128988 -16575
rect 129232 -16580 129267 -16546
rect 129277 -16580 129278 -16535
rect 129377 -16546 129378 -16535
rect 129388 -16580 129423 -16546
rect 129433 -16580 129434 -16535
rect 129533 -16546 129534 -16535
rect 130111 -16539 130146 -16505
rect 130288 -16539 130323 -16505
rect 129544 -16580 129579 -16546
rect 130431 -16565 130546 -16499
rect 130729 -16525 130730 -16499
rect 131126 -16517 131161 -16483
rect 131171 -16517 131172 -16472
rect 131271 -16483 131272 -16472
rect 131282 -16517 131317 -16483
rect 131327 -16517 131328 -16472
rect 131627 -16500 131628 -16489
rect 131832 -16494 131867 -16460
rect 131877 -16494 131878 -16449
rect 131977 -16460 131978 -16449
rect 132186 -16453 132221 -16419
rect 132231 -16453 132232 -16408
rect 132331 -16419 132332 -16408
rect 132512 -16413 132547 -16379
rect 132576 -16413 132619 -16379
rect 132621 -16413 132622 -16371
rect 132721 -16379 132722 -16371
rect 132656 -16413 132691 -16379
rect 132732 -16413 132767 -16379
rect 132777 -16413 132778 -16371
rect 132877 -16379 132878 -16371
rect 132826 -16413 132861 -16379
rect 132888 -16413 132933 -16379
rect 133928 -16408 133963 -16374
rect 133973 -16408 133974 -16363
rect 134073 -16374 134074 -16363
rect 134084 -16408 134119 -16374
rect 134129 -16408 134130 -16363
rect 134229 -16374 134230 -16363
rect 134805 -16367 134840 -16333
rect 134982 -16367 135017 -16333
rect 135575 -16336 135576 -16328
rect 135675 -16336 135676 -16328
rect 134240 -16408 134275 -16374
rect 132342 -16453 132377 -16419
rect 133621 -16422 133622 -16414
rect 134971 -16417 134972 -16406
rect 135176 -16410 135211 -16376
rect 135221 -16410 135222 -16365
rect 135321 -16376 135322 -16365
rect 135502 -16370 135565 -16336
rect 135574 -16370 135609 -16336
rect 135686 -16370 135721 -16336
rect 136411 -16360 136446 -16326
rect 136507 -16360 136542 -16326
rect 136603 -16360 136638 -16326
rect 136699 -16360 136734 -16326
rect 136795 -16360 136830 -16326
rect 136891 -16360 136926 -16326
rect 136987 -16360 137022 -16326
rect 138315 -16333 138316 -16322
rect 138492 -16327 138555 -16293
rect 138564 -16327 138599 -16293
rect 138676 -16327 138711 -16293
rect 139207 -16317 139242 -16283
rect 139303 -16317 139338 -16283
rect 139399 -16317 139434 -16283
rect 139495 -16317 139530 -16283
rect 139591 -16317 139626 -16283
rect 140616 -16324 140651 -16290
rect 140661 -16324 140662 -16279
rect 140761 -16290 140762 -16279
rect 140772 -16324 140807 -16290
rect 140817 -16324 140818 -16279
rect 140917 -16290 140918 -16279
rect 141096 -16284 141131 -16250
rect 141168 -16284 141203 -16250
rect 141240 -16284 141275 -16250
rect 141384 -16284 141419 -16250
rect 141456 -16284 141491 -16250
rect 141493 -16284 141563 -16250
rect 141600 -16284 141635 -16250
rect 141670 -16284 141705 -16250
rect 142197 -16274 142232 -16240
rect 142293 -16274 142328 -16240
rect 142389 -16274 142424 -16240
rect 143896 -16241 143931 -16207
rect 143960 -16241 144003 -16207
rect 144005 -16241 144006 -16199
rect 144105 -16207 144106 -16199
rect 144040 -16241 144075 -16207
rect 144116 -16241 144151 -16207
rect 144161 -16241 144162 -16199
rect 144261 -16207 144262 -16199
rect 144210 -16241 144245 -16207
rect 144272 -16241 144317 -16207
rect 145187 -16231 145222 -16197
rect 145283 -16231 145318 -16197
rect 145379 -16231 145414 -16197
rect 145003 -16250 145004 -16242
rect 140928 -16324 140963 -16290
rect 141909 -16293 141910 -16285
rect 142009 -16293 142010 -16285
rect 135332 -16410 135367 -16376
rect 131988 -16494 132023 -16460
rect 128998 -16620 129033 -16586
rect 130277 -16589 130278 -16578
rect 127527 -16689 127528 -16681
rect 127538 -16723 127573 -16689
rect 127758 -16734 127793 -16700
rect 126205 -16793 126240 -16759
rect 126408 -16838 126443 -16804
rect 126531 -16809 126532 -16767
rect 126853 -16796 126888 -16762
rect 126175 -16861 126176 -16853
rect 126186 -16895 126221 -16861
rect 126408 -16906 126443 -16872
rect 126175 -16961 126176 -16950
rect 126186 -16995 126221 -16961
rect 125123 -17045 125158 -17011
rect 125219 -17045 125254 -17011
rect 125315 -17045 125350 -17011
rect 125824 -17035 125859 -17001
rect 125896 -17035 125931 -17001
rect 125968 -17035 126003 -17001
rect 126040 -17029 126076 -17001
rect 126386 -17025 126421 -16991
rect 126431 -17025 126432 -16980
rect 126040 -17035 126075 -17029
rect 125477 -17088 125512 -17054
rect 125573 -17088 125608 -17054
rect 125669 -17088 125704 -17054
rect 126573 -17076 126574 -16809
rect 127202 -16819 127589 -16753
rect 126589 -16860 126624 -16826
rect 126938 -16832 126949 -16819
rect 126872 -16874 126949 -16832
rect 127000 -16874 127589 -16819
rect 127736 -16853 127771 -16819
rect 127781 -16853 127782 -16808
rect 126872 -16877 127589 -16874
rect 126589 -16928 126624 -16894
rect 126792 -16942 126827 -16908
rect 126837 -16942 126838 -16900
rect 126673 -16991 126674 -16980
rect 126684 -17025 126719 -16991
rect 126792 -17042 126827 -17008
rect 126837 -17042 126838 -16997
rect 126685 -17078 126720 -17044
rect 126757 -17078 126792 -17044
rect 126829 -17078 126864 -17044
rect 125831 -17131 125866 -17097
rect 125927 -17131 125962 -17097
rect 126023 -17131 126058 -17097
rect 126119 -17131 126154 -17097
rect 126215 -17131 126250 -17097
rect 126872 -17114 127017 -16877
rect 127202 -16899 127589 -16877
rect 127126 -16925 127589 -16899
rect 127923 -16904 127924 -16637
rect 127939 -16688 127974 -16654
rect 128553 -16691 128588 -16657
rect 129232 -16663 129267 -16629
rect 129277 -16663 129278 -16618
rect 129377 -16629 129378 -16618
rect 129388 -16663 129423 -16629
rect 129433 -16663 129434 -16618
rect 129533 -16629 129534 -16618
rect 130111 -16623 130146 -16589
rect 130288 -16623 130323 -16589
rect 130649 -16605 130684 -16571
rect 129544 -16663 129579 -16629
rect 129377 -16697 129378 -16671
rect 129776 -16689 129811 -16655
rect 129821 -16689 129822 -16644
rect 129921 -16655 129922 -16644
rect 129932 -16689 129967 -16655
rect 129977 -16689 129978 -16644
rect 130277 -16672 130278 -16661
rect 127939 -16756 127974 -16722
rect 128142 -16770 128177 -16736
rect 128187 -16770 128188 -16728
rect 128287 -16740 128288 -16729
rect 128907 -16734 128942 -16700
rect 128298 -16774 128333 -16740
rect 128023 -16819 128024 -16808
rect 128492 -16813 128527 -16779
rect 128537 -16813 128538 -16771
rect 128637 -16779 128638 -16771
rect 129297 -16777 129332 -16743
rect 128648 -16813 128683 -16779
rect 128034 -16853 128069 -16819
rect 128142 -16870 128177 -16836
rect 128187 -16870 128188 -16825
rect 128287 -16832 128288 -16821
rect 128298 -16866 128333 -16832
rect 128846 -16856 128881 -16822
rect 128891 -16856 128892 -16814
rect 128991 -16822 128992 -16814
rect 129002 -16856 129037 -16822
rect 128035 -16906 128070 -16872
rect 128107 -16906 128142 -16872
rect 128179 -16906 128214 -16872
rect 128492 -16913 128527 -16879
rect 128537 -16913 128538 -16868
rect 128637 -16879 128638 -16868
rect 128648 -16913 128683 -16879
rect 129232 -16895 129267 -16861
rect 129277 -16895 129278 -16853
rect 127126 -16959 127602 -16925
rect 128460 -16949 128495 -16915
rect 128532 -16949 128567 -16915
rect 128846 -16956 128881 -16922
rect 128891 -16956 128892 -16911
rect 128991 -16922 128992 -16911
rect 129002 -16956 129037 -16922
rect 127126 -16985 127589 -16959
rect 127130 -16993 127331 -16985
rect 127146 -17003 127315 -16993
rect 126872 -17140 127047 -17114
rect 126379 -17174 126414 -17140
rect 126475 -17174 126510 -17140
rect 126571 -17174 126606 -17140
rect 126667 -17174 126702 -17140
rect 126763 -17174 126798 -17140
rect 126859 -17174 127047 -17140
rect 126872 -17200 127047 -17174
rect 127072 -17174 127173 -17050
rect 126950 -17870 126985 -17200
rect 127072 -17228 127075 -17174
rect 126757 -17936 126902 -17924
rect 126425 -17970 126902 -17936
rect 126757 -17971 126902 -17970
rect 126938 -17971 126985 -17870
rect 127084 -17971 127119 -17174
rect 127342 -17971 127377 -17062
rect 127476 -17971 127511 -16985
rect 127729 -17002 127764 -16968
rect 127825 -17002 127860 -16968
rect 127921 -17002 127956 -16968
rect 128017 -17002 128052 -16968
rect 128113 -17002 128148 -16968
rect 128209 -17002 128244 -16968
rect 128305 -17002 128340 -16968
rect 128814 -16992 128849 -16958
rect 128886 -16992 128921 -16958
rect 129232 -16995 129267 -16961
rect 129277 -16995 129278 -16950
rect 129419 -17001 129420 -16697
rect 130111 -16706 130146 -16672
rect 130288 -16706 130323 -16672
rect 130584 -16723 130619 -16689
rect 130629 -16723 130630 -16681
rect 130771 -16753 130772 -16525
rect 131461 -16534 131496 -16500
rect 131638 -16534 131673 -16500
rect 131832 -16577 131867 -16543
rect 131877 -16577 131878 -16532
rect 131977 -16543 131978 -16532
rect 132186 -16537 132221 -16503
rect 132231 -16537 132232 -16492
rect 132331 -16503 132332 -16492
rect 132576 -16496 132611 -16462
rect 132621 -16496 132622 -16451
rect 132721 -16462 132722 -16451
rect 132732 -16496 132767 -16462
rect 132777 -16496 132778 -16451
rect 132877 -16462 132878 -16451
rect 133058 -16456 133093 -16422
rect 133130 -16456 133165 -16422
rect 133202 -16456 133237 -16422
rect 133346 -16456 133381 -16422
rect 133418 -16456 133453 -16422
rect 133455 -16456 133525 -16422
rect 133562 -16456 133597 -16422
rect 133632 -16456 133667 -16422
rect 132888 -16496 132923 -16462
rect 133928 -16491 133963 -16457
rect 133973 -16491 133974 -16446
rect 134073 -16457 134074 -16446
rect 134084 -16491 134119 -16457
rect 134129 -16491 134130 -16446
rect 134229 -16457 134230 -16446
rect 134805 -16451 134840 -16417
rect 134982 -16451 135017 -16417
rect 134240 -16491 134275 -16457
rect 132342 -16537 132377 -16503
rect 133621 -16505 133622 -16494
rect 131988 -16577 132023 -16543
rect 130901 -16621 130936 -16587
rect 131102 -16666 131137 -16632
rect 131225 -16637 131226 -16595
rect 131547 -16624 131582 -16590
rect 132186 -16620 132221 -16586
rect 132231 -16620 132232 -16575
rect 132331 -16586 132332 -16575
rect 132576 -16580 132611 -16546
rect 132621 -16580 132622 -16535
rect 132721 -16546 132722 -16535
rect 132732 -16580 132767 -16546
rect 132777 -16580 132778 -16535
rect 132877 -16546 132878 -16535
rect 133455 -16539 133490 -16505
rect 133632 -16539 133667 -16505
rect 132888 -16580 132923 -16546
rect 133775 -16565 133890 -16499
rect 134073 -16525 134074 -16499
rect 134470 -16517 134505 -16483
rect 134515 -16517 134516 -16472
rect 134615 -16483 134616 -16472
rect 134626 -16517 134661 -16483
rect 134671 -16517 134672 -16472
rect 134971 -16500 134972 -16489
rect 135176 -16494 135211 -16460
rect 135221 -16494 135222 -16449
rect 135321 -16460 135322 -16449
rect 135530 -16453 135565 -16419
rect 135575 -16453 135576 -16408
rect 135675 -16419 135676 -16408
rect 135856 -16413 135891 -16379
rect 135920 -16413 135963 -16379
rect 135965 -16413 135966 -16371
rect 136065 -16379 136066 -16371
rect 136000 -16413 136035 -16379
rect 136076 -16413 136111 -16379
rect 136121 -16413 136122 -16371
rect 136221 -16379 136222 -16371
rect 136170 -16413 136205 -16379
rect 136232 -16413 136277 -16379
rect 137272 -16408 137307 -16374
rect 137317 -16408 137318 -16363
rect 137417 -16374 137418 -16363
rect 137428 -16408 137463 -16374
rect 137473 -16408 137474 -16363
rect 137573 -16374 137574 -16363
rect 138149 -16367 138184 -16333
rect 138326 -16367 138361 -16333
rect 138919 -16336 138920 -16328
rect 139019 -16336 139020 -16328
rect 137584 -16408 137619 -16374
rect 135686 -16453 135721 -16419
rect 136965 -16422 136966 -16414
rect 138315 -16417 138316 -16406
rect 138520 -16410 138555 -16376
rect 138565 -16410 138566 -16365
rect 138665 -16376 138666 -16365
rect 138846 -16370 138909 -16336
rect 138918 -16370 138953 -16336
rect 139030 -16370 139065 -16336
rect 139755 -16360 139790 -16326
rect 139851 -16360 139886 -16326
rect 139947 -16360 139982 -16326
rect 140043 -16360 140078 -16326
rect 140139 -16360 140174 -16326
rect 140235 -16360 140270 -16326
rect 140331 -16360 140366 -16326
rect 141659 -16333 141660 -16322
rect 141836 -16327 141899 -16293
rect 141908 -16327 141943 -16293
rect 142020 -16327 142055 -16293
rect 142551 -16317 142586 -16283
rect 142647 -16317 142682 -16283
rect 142743 -16317 142778 -16283
rect 142839 -16317 142874 -16283
rect 142935 -16317 142970 -16283
rect 143960 -16324 143995 -16290
rect 144005 -16324 144006 -16279
rect 144105 -16290 144106 -16279
rect 144116 -16324 144151 -16290
rect 144161 -16324 144162 -16279
rect 144261 -16290 144262 -16279
rect 144440 -16284 144475 -16250
rect 144512 -16284 144547 -16250
rect 144584 -16284 144619 -16250
rect 144728 -16284 144763 -16250
rect 144800 -16284 144835 -16250
rect 144837 -16284 144907 -16250
rect 144944 -16284 144979 -16250
rect 145014 -16284 145049 -16250
rect 145541 -16274 145576 -16240
rect 145637 -16274 145672 -16240
rect 145733 -16274 145768 -16240
rect 147240 -16241 147275 -16207
rect 147304 -16241 147347 -16207
rect 147349 -16241 147350 -16199
rect 147449 -16207 147450 -16199
rect 147384 -16241 147419 -16207
rect 147460 -16241 147495 -16207
rect 147505 -16241 147506 -16199
rect 147605 -16207 147606 -16199
rect 147554 -16241 147589 -16207
rect 147616 -16241 147661 -16207
rect 148531 -16231 148566 -16197
rect 148627 -16231 148662 -16197
rect 148723 -16231 148758 -16197
rect 148347 -16250 148348 -16242
rect 144272 -16324 144307 -16290
rect 145253 -16293 145254 -16285
rect 145353 -16293 145354 -16285
rect 138676 -16410 138711 -16376
rect 135332 -16494 135367 -16460
rect 132342 -16620 132377 -16586
rect 133621 -16589 133622 -16578
rect 130871 -16689 130872 -16681
rect 130882 -16723 130917 -16689
rect 131102 -16734 131137 -16700
rect 129549 -16793 129584 -16759
rect 129752 -16838 129787 -16804
rect 129875 -16809 129876 -16767
rect 130197 -16796 130232 -16762
rect 129519 -16861 129520 -16853
rect 129530 -16895 129565 -16861
rect 129752 -16906 129787 -16872
rect 129519 -16961 129520 -16950
rect 129530 -16995 129565 -16961
rect 128467 -17045 128502 -17011
rect 128563 -17045 128598 -17011
rect 128659 -17045 128694 -17011
rect 129168 -17035 129203 -17001
rect 129240 -17035 129275 -17001
rect 129312 -17035 129347 -17001
rect 129384 -17029 129420 -17001
rect 129730 -17025 129765 -16991
rect 129775 -17025 129776 -16980
rect 129384 -17035 129419 -17029
rect 128821 -17088 128856 -17054
rect 128917 -17088 128952 -17054
rect 129013 -17088 129048 -17054
rect 129917 -17076 129918 -16809
rect 130546 -16819 130933 -16753
rect 129933 -16860 129968 -16826
rect 130282 -16832 130293 -16819
rect 130216 -16874 130293 -16832
rect 130344 -16874 130933 -16819
rect 131080 -16853 131115 -16819
rect 131125 -16853 131126 -16808
rect 130216 -16877 130933 -16874
rect 129933 -16928 129968 -16894
rect 130136 -16942 130171 -16908
rect 130181 -16942 130182 -16900
rect 130017 -16991 130018 -16980
rect 130028 -17025 130063 -16991
rect 130136 -17042 130171 -17008
rect 130181 -17042 130182 -16997
rect 130029 -17078 130064 -17044
rect 130101 -17078 130136 -17044
rect 130173 -17078 130208 -17044
rect 129175 -17131 129210 -17097
rect 129271 -17131 129306 -17097
rect 129367 -17131 129402 -17097
rect 129463 -17131 129498 -17097
rect 129559 -17131 129594 -17097
rect 130216 -17114 130361 -16877
rect 130546 -16899 130933 -16877
rect 130470 -16925 130933 -16899
rect 131267 -16904 131268 -16637
rect 131283 -16688 131318 -16654
rect 131897 -16691 131932 -16657
rect 132576 -16663 132611 -16629
rect 132621 -16663 132622 -16618
rect 132721 -16629 132722 -16618
rect 132732 -16663 132767 -16629
rect 132777 -16663 132778 -16618
rect 132877 -16629 132878 -16618
rect 133455 -16623 133490 -16589
rect 133632 -16623 133667 -16589
rect 133993 -16605 134028 -16571
rect 132888 -16663 132923 -16629
rect 132721 -16697 132722 -16671
rect 133120 -16689 133155 -16655
rect 133165 -16689 133166 -16644
rect 133265 -16655 133266 -16644
rect 133276 -16689 133311 -16655
rect 133321 -16689 133322 -16644
rect 133621 -16672 133622 -16661
rect 131283 -16756 131318 -16722
rect 131486 -16770 131521 -16736
rect 131531 -16770 131532 -16728
rect 131631 -16740 131632 -16729
rect 132251 -16734 132286 -16700
rect 131642 -16774 131677 -16740
rect 131367 -16819 131368 -16808
rect 131836 -16813 131871 -16779
rect 131881 -16813 131882 -16771
rect 131981 -16779 131982 -16771
rect 132641 -16777 132676 -16743
rect 131992 -16813 132027 -16779
rect 131378 -16853 131413 -16819
rect 131486 -16870 131521 -16836
rect 131531 -16870 131532 -16825
rect 131631 -16832 131632 -16821
rect 131642 -16866 131677 -16832
rect 132190 -16856 132225 -16822
rect 132235 -16856 132236 -16814
rect 132335 -16822 132336 -16814
rect 132346 -16856 132381 -16822
rect 131379 -16906 131414 -16872
rect 131451 -16906 131486 -16872
rect 131523 -16906 131558 -16872
rect 131836 -16913 131871 -16879
rect 131881 -16913 131882 -16868
rect 131981 -16879 131982 -16868
rect 131992 -16913 132027 -16879
rect 132576 -16895 132611 -16861
rect 132621 -16895 132622 -16853
rect 130470 -16959 130946 -16925
rect 131804 -16949 131839 -16915
rect 131876 -16949 131911 -16915
rect 132190 -16956 132225 -16922
rect 132235 -16956 132236 -16911
rect 132335 -16922 132336 -16911
rect 132346 -16956 132381 -16922
rect 130470 -16985 130933 -16959
rect 130474 -16993 130675 -16985
rect 130490 -17003 130659 -16993
rect 130216 -17140 130391 -17114
rect 129723 -17174 129758 -17140
rect 129819 -17174 129854 -17140
rect 129915 -17174 129950 -17140
rect 130011 -17174 130046 -17140
rect 130107 -17174 130142 -17140
rect 130203 -17174 130391 -17140
rect 130216 -17200 130391 -17174
rect 130416 -17174 130517 -17050
rect 130294 -17870 130329 -17200
rect 130416 -17228 130419 -17174
rect 130101 -17936 130246 -17924
rect 129769 -17970 130246 -17936
rect 130101 -17971 130246 -17970
rect 130282 -17971 130329 -17870
rect 130428 -17971 130463 -17174
rect 130686 -17971 130721 -17062
rect 130820 -17971 130855 -16985
rect 131073 -17002 131108 -16968
rect 131169 -17002 131204 -16968
rect 131265 -17002 131300 -16968
rect 131361 -17002 131396 -16968
rect 131457 -17002 131492 -16968
rect 131553 -17002 131588 -16968
rect 131649 -17002 131684 -16968
rect 132158 -16992 132193 -16958
rect 132230 -16992 132265 -16958
rect 132576 -16995 132611 -16961
rect 132621 -16995 132622 -16950
rect 132763 -17001 132764 -16697
rect 133455 -16706 133490 -16672
rect 133632 -16706 133667 -16672
rect 133928 -16723 133963 -16689
rect 133973 -16723 133974 -16681
rect 134115 -16753 134116 -16525
rect 134805 -16534 134840 -16500
rect 134982 -16534 135017 -16500
rect 135176 -16577 135211 -16543
rect 135221 -16577 135222 -16532
rect 135321 -16543 135322 -16532
rect 135530 -16537 135565 -16503
rect 135575 -16537 135576 -16492
rect 135675 -16503 135676 -16492
rect 135920 -16496 135955 -16462
rect 135965 -16496 135966 -16451
rect 136065 -16462 136066 -16451
rect 136076 -16496 136111 -16462
rect 136121 -16496 136122 -16451
rect 136221 -16462 136222 -16451
rect 136402 -16456 136437 -16422
rect 136474 -16456 136509 -16422
rect 136546 -16456 136581 -16422
rect 136690 -16456 136725 -16422
rect 136762 -16456 136797 -16422
rect 136799 -16456 136869 -16422
rect 136906 -16456 136941 -16422
rect 136976 -16456 137011 -16422
rect 136232 -16496 136267 -16462
rect 137272 -16491 137307 -16457
rect 137317 -16491 137318 -16446
rect 137417 -16457 137418 -16446
rect 137428 -16491 137463 -16457
rect 137473 -16491 137474 -16446
rect 137573 -16457 137574 -16446
rect 138149 -16451 138184 -16417
rect 138326 -16451 138361 -16417
rect 137584 -16491 137619 -16457
rect 135686 -16537 135721 -16503
rect 136965 -16505 136966 -16494
rect 135332 -16577 135367 -16543
rect 134245 -16621 134280 -16587
rect 134446 -16666 134481 -16632
rect 134569 -16637 134570 -16595
rect 134891 -16624 134926 -16590
rect 135530 -16620 135565 -16586
rect 135575 -16620 135576 -16575
rect 135675 -16586 135676 -16575
rect 135920 -16580 135955 -16546
rect 135965 -16580 135966 -16535
rect 136065 -16546 136066 -16535
rect 136076 -16580 136111 -16546
rect 136121 -16580 136122 -16535
rect 136221 -16546 136222 -16535
rect 136799 -16539 136834 -16505
rect 136976 -16539 137011 -16505
rect 136232 -16580 136267 -16546
rect 137119 -16565 137234 -16499
rect 137417 -16525 137418 -16499
rect 137814 -16517 137849 -16483
rect 137859 -16517 137860 -16472
rect 137959 -16483 137960 -16472
rect 137970 -16517 138005 -16483
rect 138015 -16517 138016 -16472
rect 138315 -16500 138316 -16489
rect 138520 -16494 138555 -16460
rect 138565 -16494 138566 -16449
rect 138665 -16460 138666 -16449
rect 138874 -16453 138909 -16419
rect 138919 -16453 138920 -16408
rect 139019 -16419 139020 -16408
rect 139200 -16413 139235 -16379
rect 139264 -16413 139307 -16379
rect 139309 -16413 139310 -16371
rect 139409 -16379 139410 -16371
rect 139344 -16413 139379 -16379
rect 139420 -16413 139455 -16379
rect 139465 -16413 139466 -16371
rect 139565 -16379 139566 -16371
rect 139514 -16413 139549 -16379
rect 139576 -16413 139621 -16379
rect 140616 -16408 140651 -16374
rect 140661 -16408 140662 -16363
rect 140761 -16374 140762 -16363
rect 140772 -16408 140807 -16374
rect 140817 -16408 140818 -16363
rect 140917 -16374 140918 -16363
rect 141493 -16367 141528 -16333
rect 141670 -16367 141705 -16333
rect 142263 -16336 142264 -16328
rect 142363 -16336 142364 -16328
rect 140928 -16408 140963 -16374
rect 139030 -16453 139065 -16419
rect 140309 -16422 140310 -16414
rect 141659 -16417 141660 -16406
rect 141864 -16410 141899 -16376
rect 141909 -16410 141910 -16365
rect 142009 -16376 142010 -16365
rect 142190 -16370 142253 -16336
rect 142262 -16370 142297 -16336
rect 142374 -16370 142409 -16336
rect 143099 -16360 143134 -16326
rect 143195 -16360 143230 -16326
rect 143291 -16360 143326 -16326
rect 143387 -16360 143422 -16326
rect 143483 -16360 143518 -16326
rect 143579 -16360 143614 -16326
rect 143675 -16360 143710 -16326
rect 145003 -16333 145004 -16322
rect 145180 -16327 145243 -16293
rect 145252 -16327 145287 -16293
rect 145364 -16327 145399 -16293
rect 145895 -16317 145930 -16283
rect 145991 -16317 146026 -16283
rect 146087 -16317 146122 -16283
rect 146183 -16317 146218 -16283
rect 146279 -16317 146314 -16283
rect 147304 -16324 147339 -16290
rect 147349 -16324 147350 -16279
rect 147449 -16290 147450 -16279
rect 147460 -16324 147495 -16290
rect 147505 -16324 147506 -16279
rect 147605 -16290 147606 -16279
rect 147784 -16284 147819 -16250
rect 147856 -16284 147891 -16250
rect 147928 -16284 147963 -16250
rect 148072 -16284 148107 -16250
rect 148144 -16284 148179 -16250
rect 148181 -16284 148251 -16250
rect 148288 -16284 148323 -16250
rect 148358 -16284 148393 -16250
rect 148885 -16274 148920 -16240
rect 148981 -16274 149016 -16240
rect 149077 -16274 149112 -16240
rect 150584 -16241 150619 -16207
rect 150648 -16241 150691 -16207
rect 150693 -16241 150694 -16199
rect 150793 -16207 150794 -16199
rect 150728 -16241 150763 -16207
rect 150804 -16241 150839 -16207
rect 150849 -16241 150850 -16199
rect 150949 -16207 150950 -16199
rect 150898 -16241 150933 -16207
rect 150960 -16241 151005 -16207
rect 151875 -16231 151910 -16197
rect 151971 -16231 152006 -16197
rect 152067 -16231 152102 -16197
rect 151691 -16250 151692 -16242
rect 147616 -16324 147651 -16290
rect 148597 -16293 148598 -16285
rect 148697 -16293 148698 -16285
rect 142020 -16410 142055 -16376
rect 138676 -16494 138711 -16460
rect 135686 -16620 135721 -16586
rect 136965 -16589 136966 -16578
rect 134215 -16689 134216 -16681
rect 134226 -16723 134261 -16689
rect 134446 -16734 134481 -16700
rect 132893 -16793 132928 -16759
rect 133096 -16838 133131 -16804
rect 133219 -16809 133220 -16767
rect 133541 -16796 133576 -16762
rect 132863 -16861 132864 -16853
rect 132874 -16895 132909 -16861
rect 133096 -16906 133131 -16872
rect 132863 -16961 132864 -16950
rect 132874 -16995 132909 -16961
rect 131811 -17045 131846 -17011
rect 131907 -17045 131942 -17011
rect 132003 -17045 132038 -17011
rect 132512 -17035 132547 -17001
rect 132584 -17035 132619 -17001
rect 132656 -17035 132691 -17001
rect 132728 -17029 132764 -17001
rect 133074 -17025 133109 -16991
rect 133119 -17025 133120 -16980
rect 132728 -17035 132763 -17029
rect 132165 -17088 132200 -17054
rect 132261 -17088 132296 -17054
rect 132357 -17088 132392 -17054
rect 133261 -17076 133262 -16809
rect 133890 -16819 134277 -16753
rect 133277 -16860 133312 -16826
rect 133626 -16832 133637 -16819
rect 133560 -16874 133637 -16832
rect 133688 -16874 134277 -16819
rect 134424 -16853 134459 -16819
rect 134469 -16853 134470 -16808
rect 133560 -16877 134277 -16874
rect 133277 -16928 133312 -16894
rect 133480 -16942 133515 -16908
rect 133525 -16942 133526 -16900
rect 133361 -16991 133362 -16980
rect 133372 -17025 133407 -16991
rect 133480 -17042 133515 -17008
rect 133525 -17042 133526 -16997
rect 133373 -17078 133408 -17044
rect 133445 -17078 133480 -17044
rect 133517 -17078 133552 -17044
rect 132519 -17131 132554 -17097
rect 132615 -17131 132650 -17097
rect 132711 -17131 132746 -17097
rect 132807 -17131 132842 -17097
rect 132903 -17131 132938 -17097
rect 133560 -17114 133705 -16877
rect 133890 -16899 134277 -16877
rect 133814 -16925 134277 -16899
rect 134611 -16904 134612 -16637
rect 134627 -16688 134662 -16654
rect 135241 -16691 135276 -16657
rect 135920 -16663 135955 -16629
rect 135965 -16663 135966 -16618
rect 136065 -16629 136066 -16618
rect 136076 -16663 136111 -16629
rect 136121 -16663 136122 -16618
rect 136221 -16629 136222 -16618
rect 136799 -16623 136834 -16589
rect 136976 -16623 137011 -16589
rect 137337 -16605 137372 -16571
rect 136232 -16663 136267 -16629
rect 136065 -16697 136066 -16671
rect 136464 -16689 136499 -16655
rect 136509 -16689 136510 -16644
rect 136609 -16655 136610 -16644
rect 136620 -16689 136655 -16655
rect 136665 -16689 136666 -16644
rect 136965 -16672 136966 -16661
rect 134627 -16756 134662 -16722
rect 134830 -16770 134865 -16736
rect 134875 -16770 134876 -16728
rect 134975 -16740 134976 -16729
rect 135595 -16734 135630 -16700
rect 134986 -16774 135021 -16740
rect 134711 -16819 134712 -16808
rect 135180 -16813 135215 -16779
rect 135225 -16813 135226 -16771
rect 135325 -16779 135326 -16771
rect 135985 -16777 136020 -16743
rect 135336 -16813 135371 -16779
rect 134722 -16853 134757 -16819
rect 134830 -16870 134865 -16836
rect 134875 -16870 134876 -16825
rect 134975 -16832 134976 -16821
rect 134986 -16866 135021 -16832
rect 135534 -16856 135569 -16822
rect 135579 -16856 135580 -16814
rect 135679 -16822 135680 -16814
rect 135690 -16856 135725 -16822
rect 134723 -16906 134758 -16872
rect 134795 -16906 134830 -16872
rect 134867 -16906 134902 -16872
rect 135180 -16913 135215 -16879
rect 135225 -16913 135226 -16868
rect 135325 -16879 135326 -16868
rect 135336 -16913 135371 -16879
rect 135920 -16895 135955 -16861
rect 135965 -16895 135966 -16853
rect 133814 -16959 134290 -16925
rect 135148 -16949 135183 -16915
rect 135220 -16949 135255 -16915
rect 135534 -16956 135569 -16922
rect 135579 -16956 135580 -16911
rect 135679 -16922 135680 -16911
rect 135690 -16956 135725 -16922
rect 133814 -16985 134277 -16959
rect 133818 -16993 134019 -16985
rect 133834 -17003 134003 -16993
rect 133560 -17140 133735 -17114
rect 133067 -17174 133102 -17140
rect 133163 -17174 133198 -17140
rect 133259 -17174 133294 -17140
rect 133355 -17174 133390 -17140
rect 133451 -17174 133486 -17140
rect 133547 -17174 133735 -17140
rect 133560 -17200 133735 -17174
rect 133760 -17174 133861 -17050
rect 133638 -17870 133673 -17200
rect 133760 -17228 133763 -17174
rect 133445 -17936 133590 -17924
rect 133113 -17970 133590 -17936
rect 133445 -17971 133590 -17970
rect 133626 -17971 133673 -17870
rect 133772 -17971 133807 -17174
rect 134030 -17971 134065 -17062
rect 134164 -17971 134199 -16985
rect 134417 -17002 134452 -16968
rect 134513 -17002 134548 -16968
rect 134609 -17002 134644 -16968
rect 134705 -17002 134740 -16968
rect 134801 -17002 134836 -16968
rect 134897 -17002 134932 -16968
rect 134993 -17002 135028 -16968
rect 135502 -16992 135537 -16958
rect 135574 -16992 135609 -16958
rect 135920 -16995 135955 -16961
rect 135965 -16995 135966 -16950
rect 136107 -17001 136108 -16697
rect 136799 -16706 136834 -16672
rect 136976 -16706 137011 -16672
rect 137272 -16723 137307 -16689
rect 137317 -16723 137318 -16681
rect 137459 -16753 137460 -16525
rect 138149 -16534 138184 -16500
rect 138326 -16534 138361 -16500
rect 138520 -16577 138555 -16543
rect 138565 -16577 138566 -16532
rect 138665 -16543 138666 -16532
rect 138874 -16537 138909 -16503
rect 138919 -16537 138920 -16492
rect 139019 -16503 139020 -16492
rect 139264 -16496 139299 -16462
rect 139309 -16496 139310 -16451
rect 139409 -16462 139410 -16451
rect 139420 -16496 139455 -16462
rect 139465 -16496 139466 -16451
rect 139565 -16462 139566 -16451
rect 139746 -16456 139781 -16422
rect 139818 -16456 139853 -16422
rect 139890 -16456 139925 -16422
rect 140034 -16456 140069 -16422
rect 140106 -16456 140141 -16422
rect 140143 -16456 140213 -16422
rect 140250 -16456 140285 -16422
rect 140320 -16456 140355 -16422
rect 139576 -16496 139611 -16462
rect 140616 -16491 140651 -16457
rect 140661 -16491 140662 -16446
rect 140761 -16457 140762 -16446
rect 140772 -16491 140807 -16457
rect 140817 -16491 140818 -16446
rect 140917 -16457 140918 -16446
rect 141493 -16451 141528 -16417
rect 141670 -16451 141705 -16417
rect 140928 -16491 140963 -16457
rect 139030 -16537 139065 -16503
rect 140309 -16505 140310 -16494
rect 138676 -16577 138711 -16543
rect 137589 -16621 137624 -16587
rect 137790 -16666 137825 -16632
rect 137913 -16637 137914 -16595
rect 138235 -16624 138270 -16590
rect 138874 -16620 138909 -16586
rect 138919 -16620 138920 -16575
rect 139019 -16586 139020 -16575
rect 139264 -16580 139299 -16546
rect 139309 -16580 139310 -16535
rect 139409 -16546 139410 -16535
rect 139420 -16580 139455 -16546
rect 139465 -16580 139466 -16535
rect 139565 -16546 139566 -16535
rect 140143 -16539 140178 -16505
rect 140320 -16539 140355 -16505
rect 139576 -16580 139611 -16546
rect 140463 -16565 140578 -16499
rect 140761 -16525 140762 -16499
rect 141158 -16517 141193 -16483
rect 141203 -16517 141204 -16472
rect 141303 -16483 141304 -16472
rect 141314 -16517 141349 -16483
rect 141359 -16517 141360 -16472
rect 141659 -16500 141660 -16489
rect 141864 -16494 141899 -16460
rect 141909 -16494 141910 -16449
rect 142009 -16460 142010 -16449
rect 142218 -16453 142253 -16419
rect 142263 -16453 142264 -16408
rect 142363 -16419 142364 -16408
rect 142544 -16413 142579 -16379
rect 142608 -16413 142651 -16379
rect 142653 -16413 142654 -16371
rect 142753 -16379 142754 -16371
rect 142688 -16413 142723 -16379
rect 142764 -16413 142799 -16379
rect 142809 -16413 142810 -16371
rect 142909 -16379 142910 -16371
rect 142858 -16413 142893 -16379
rect 142920 -16413 142965 -16379
rect 143960 -16408 143995 -16374
rect 144005 -16408 144006 -16363
rect 144105 -16374 144106 -16363
rect 144116 -16408 144151 -16374
rect 144161 -16408 144162 -16363
rect 144261 -16374 144262 -16363
rect 144837 -16367 144872 -16333
rect 145014 -16367 145049 -16333
rect 145607 -16336 145608 -16328
rect 145707 -16336 145708 -16328
rect 144272 -16408 144307 -16374
rect 142374 -16453 142409 -16419
rect 143653 -16422 143654 -16414
rect 145003 -16417 145004 -16406
rect 145208 -16410 145243 -16376
rect 145253 -16410 145254 -16365
rect 145353 -16376 145354 -16365
rect 145534 -16370 145597 -16336
rect 145606 -16370 145641 -16336
rect 145718 -16370 145753 -16336
rect 146443 -16360 146478 -16326
rect 146539 -16360 146574 -16326
rect 146635 -16360 146670 -16326
rect 146731 -16360 146766 -16326
rect 146827 -16360 146862 -16326
rect 146923 -16360 146958 -16326
rect 147019 -16360 147054 -16326
rect 148347 -16333 148348 -16322
rect 148524 -16327 148587 -16293
rect 148596 -16327 148631 -16293
rect 148708 -16327 148743 -16293
rect 149239 -16317 149274 -16283
rect 149335 -16317 149370 -16283
rect 149431 -16317 149466 -16283
rect 149527 -16317 149562 -16283
rect 149623 -16317 149658 -16283
rect 150648 -16324 150683 -16290
rect 150693 -16324 150694 -16279
rect 150793 -16290 150794 -16279
rect 150804 -16324 150839 -16290
rect 150849 -16324 150850 -16279
rect 150949 -16290 150950 -16279
rect 151128 -16284 151163 -16250
rect 151200 -16284 151235 -16250
rect 151272 -16284 151307 -16250
rect 151416 -16284 151451 -16250
rect 151488 -16284 151523 -16250
rect 151525 -16284 151595 -16250
rect 151632 -16284 151667 -16250
rect 151702 -16284 151737 -16250
rect 152229 -16274 152264 -16240
rect 152325 -16274 152360 -16240
rect 152421 -16274 152456 -16240
rect 153928 -16241 153963 -16207
rect 153992 -16241 154035 -16207
rect 154037 -16241 154038 -16199
rect 154137 -16207 154138 -16199
rect 154072 -16241 154107 -16207
rect 154148 -16241 154183 -16207
rect 154193 -16241 154194 -16199
rect 154293 -16207 154294 -16199
rect 154242 -16241 154277 -16207
rect 154304 -16241 154349 -16207
rect 155219 -16231 155254 -16197
rect 155315 -16231 155350 -16197
rect 155411 -16231 155446 -16197
rect 155035 -16250 155036 -16242
rect 150960 -16324 150995 -16290
rect 151941 -16293 151942 -16285
rect 152041 -16293 152042 -16285
rect 145364 -16410 145399 -16376
rect 142020 -16494 142055 -16460
rect 139030 -16620 139065 -16586
rect 140309 -16589 140310 -16578
rect 137559 -16689 137560 -16681
rect 137570 -16723 137605 -16689
rect 137790 -16734 137825 -16700
rect 136237 -16793 136272 -16759
rect 136440 -16838 136475 -16804
rect 136563 -16809 136564 -16767
rect 136885 -16796 136920 -16762
rect 136207 -16861 136208 -16853
rect 136218 -16895 136253 -16861
rect 136440 -16906 136475 -16872
rect 136207 -16961 136208 -16950
rect 136218 -16995 136253 -16961
rect 135155 -17045 135190 -17011
rect 135251 -17045 135286 -17011
rect 135347 -17045 135382 -17011
rect 135856 -17035 135891 -17001
rect 135928 -17035 135963 -17001
rect 136000 -17035 136035 -17001
rect 136072 -17029 136108 -17001
rect 136418 -17025 136453 -16991
rect 136463 -17025 136464 -16980
rect 136072 -17035 136107 -17029
rect 135509 -17088 135544 -17054
rect 135605 -17088 135640 -17054
rect 135701 -17088 135736 -17054
rect 136605 -17076 136606 -16809
rect 137234 -16819 137621 -16753
rect 136621 -16860 136656 -16826
rect 136970 -16832 136981 -16819
rect 136904 -16874 136981 -16832
rect 137032 -16874 137621 -16819
rect 137768 -16853 137803 -16819
rect 137813 -16853 137814 -16808
rect 136904 -16877 137621 -16874
rect 136621 -16928 136656 -16894
rect 136824 -16942 136859 -16908
rect 136869 -16942 136870 -16900
rect 136705 -16991 136706 -16980
rect 136716 -17025 136751 -16991
rect 136824 -17042 136859 -17008
rect 136869 -17042 136870 -16997
rect 136717 -17078 136752 -17044
rect 136789 -17078 136824 -17044
rect 136861 -17078 136896 -17044
rect 135863 -17131 135898 -17097
rect 135959 -17131 135994 -17097
rect 136055 -17131 136090 -17097
rect 136151 -17131 136186 -17097
rect 136247 -17131 136282 -17097
rect 136904 -17114 137049 -16877
rect 137234 -16899 137621 -16877
rect 137158 -16925 137621 -16899
rect 137955 -16904 137956 -16637
rect 137971 -16688 138006 -16654
rect 138585 -16691 138620 -16657
rect 139264 -16663 139299 -16629
rect 139309 -16663 139310 -16618
rect 139409 -16629 139410 -16618
rect 139420 -16663 139455 -16629
rect 139465 -16663 139466 -16618
rect 139565 -16629 139566 -16618
rect 140143 -16623 140178 -16589
rect 140320 -16623 140355 -16589
rect 140681 -16605 140716 -16571
rect 139576 -16663 139611 -16629
rect 139409 -16697 139410 -16671
rect 139808 -16689 139843 -16655
rect 139853 -16689 139854 -16644
rect 139953 -16655 139954 -16644
rect 139964 -16689 139999 -16655
rect 140009 -16689 140010 -16644
rect 140309 -16672 140310 -16661
rect 137971 -16756 138006 -16722
rect 138174 -16770 138209 -16736
rect 138219 -16770 138220 -16728
rect 138319 -16740 138320 -16729
rect 138939 -16734 138974 -16700
rect 138330 -16774 138365 -16740
rect 138055 -16819 138056 -16808
rect 138524 -16813 138559 -16779
rect 138569 -16813 138570 -16771
rect 138669 -16779 138670 -16771
rect 139329 -16777 139364 -16743
rect 138680 -16813 138715 -16779
rect 138066 -16853 138101 -16819
rect 138174 -16870 138209 -16836
rect 138219 -16870 138220 -16825
rect 138319 -16832 138320 -16821
rect 138330 -16866 138365 -16832
rect 138878 -16856 138913 -16822
rect 138923 -16856 138924 -16814
rect 139023 -16822 139024 -16814
rect 139034 -16856 139069 -16822
rect 138067 -16906 138102 -16872
rect 138139 -16906 138174 -16872
rect 138211 -16906 138246 -16872
rect 138524 -16913 138559 -16879
rect 138569 -16913 138570 -16868
rect 138669 -16879 138670 -16868
rect 138680 -16913 138715 -16879
rect 139264 -16895 139299 -16861
rect 139309 -16895 139310 -16853
rect 137158 -16959 137634 -16925
rect 138492 -16949 138527 -16915
rect 138564 -16949 138599 -16915
rect 138878 -16956 138913 -16922
rect 138923 -16956 138924 -16911
rect 139023 -16922 139024 -16911
rect 139034 -16956 139069 -16922
rect 137158 -16985 137621 -16959
rect 137162 -16993 137363 -16985
rect 137178 -17003 137347 -16993
rect 136904 -17140 137079 -17114
rect 136411 -17174 136446 -17140
rect 136507 -17174 136542 -17140
rect 136603 -17174 136638 -17140
rect 136699 -17174 136734 -17140
rect 136795 -17174 136830 -17140
rect 136891 -17174 137079 -17140
rect 136904 -17200 137079 -17174
rect 137104 -17174 137205 -17050
rect 136982 -17870 137017 -17200
rect 137104 -17228 137107 -17174
rect 136789 -17936 136934 -17924
rect 136457 -17970 136934 -17936
rect 136789 -17971 136934 -17970
rect 136970 -17971 137017 -17870
rect 137116 -17971 137151 -17174
rect 137374 -17971 137409 -17062
rect 137508 -17971 137543 -16985
rect 137761 -17002 137796 -16968
rect 137857 -17002 137892 -16968
rect 137953 -17002 137988 -16968
rect 138049 -17002 138084 -16968
rect 138145 -17002 138180 -16968
rect 138241 -17002 138276 -16968
rect 138337 -17002 138372 -16968
rect 138846 -16992 138881 -16958
rect 138918 -16992 138953 -16958
rect 139264 -16995 139299 -16961
rect 139309 -16995 139310 -16950
rect 139451 -17001 139452 -16697
rect 140143 -16706 140178 -16672
rect 140320 -16706 140355 -16672
rect 140616 -16723 140651 -16689
rect 140661 -16723 140662 -16681
rect 140803 -16753 140804 -16525
rect 141493 -16534 141528 -16500
rect 141670 -16534 141705 -16500
rect 141864 -16577 141899 -16543
rect 141909 -16577 141910 -16532
rect 142009 -16543 142010 -16532
rect 142218 -16537 142253 -16503
rect 142263 -16537 142264 -16492
rect 142363 -16503 142364 -16492
rect 142608 -16496 142643 -16462
rect 142653 -16496 142654 -16451
rect 142753 -16462 142754 -16451
rect 142764 -16496 142799 -16462
rect 142809 -16496 142810 -16451
rect 142909 -16462 142910 -16451
rect 143090 -16456 143125 -16422
rect 143162 -16456 143197 -16422
rect 143234 -16456 143269 -16422
rect 143378 -16456 143413 -16422
rect 143450 -16456 143485 -16422
rect 143487 -16456 143557 -16422
rect 143594 -16456 143629 -16422
rect 143664 -16456 143699 -16422
rect 142920 -16496 142955 -16462
rect 143960 -16491 143995 -16457
rect 144005 -16491 144006 -16446
rect 144105 -16457 144106 -16446
rect 144116 -16491 144151 -16457
rect 144161 -16491 144162 -16446
rect 144261 -16457 144262 -16446
rect 144837 -16451 144872 -16417
rect 145014 -16451 145049 -16417
rect 144272 -16491 144307 -16457
rect 142374 -16537 142409 -16503
rect 143653 -16505 143654 -16494
rect 142020 -16577 142055 -16543
rect 140933 -16621 140968 -16587
rect 141134 -16666 141169 -16632
rect 141257 -16637 141258 -16595
rect 141579 -16624 141614 -16590
rect 142218 -16620 142253 -16586
rect 142263 -16620 142264 -16575
rect 142363 -16586 142364 -16575
rect 142608 -16580 142643 -16546
rect 142653 -16580 142654 -16535
rect 142753 -16546 142754 -16535
rect 142764 -16580 142799 -16546
rect 142809 -16580 142810 -16535
rect 142909 -16546 142910 -16535
rect 143487 -16539 143522 -16505
rect 143664 -16539 143699 -16505
rect 142920 -16580 142955 -16546
rect 143807 -16565 143922 -16499
rect 144105 -16525 144106 -16499
rect 144502 -16517 144537 -16483
rect 144547 -16517 144548 -16472
rect 144647 -16483 144648 -16472
rect 144658 -16517 144693 -16483
rect 144703 -16517 144704 -16472
rect 145003 -16500 145004 -16489
rect 145208 -16494 145243 -16460
rect 145253 -16494 145254 -16449
rect 145353 -16460 145354 -16449
rect 145562 -16453 145597 -16419
rect 145607 -16453 145608 -16408
rect 145707 -16419 145708 -16408
rect 145888 -16413 145923 -16379
rect 145952 -16413 145995 -16379
rect 145997 -16413 145998 -16371
rect 146097 -16379 146098 -16371
rect 146032 -16413 146067 -16379
rect 146108 -16413 146143 -16379
rect 146153 -16413 146154 -16371
rect 146253 -16379 146254 -16371
rect 146202 -16413 146237 -16379
rect 146264 -16413 146309 -16379
rect 147304 -16408 147339 -16374
rect 147349 -16408 147350 -16363
rect 147449 -16374 147450 -16363
rect 147460 -16408 147495 -16374
rect 147505 -16408 147506 -16363
rect 147605 -16374 147606 -16363
rect 148181 -16367 148216 -16333
rect 148358 -16367 148393 -16333
rect 148951 -16336 148952 -16328
rect 149051 -16336 149052 -16328
rect 147616 -16408 147651 -16374
rect 145718 -16453 145753 -16419
rect 146997 -16422 146998 -16414
rect 148347 -16417 148348 -16406
rect 148552 -16410 148587 -16376
rect 148597 -16410 148598 -16365
rect 148697 -16376 148698 -16365
rect 148878 -16370 148941 -16336
rect 148950 -16370 148985 -16336
rect 149062 -16370 149097 -16336
rect 149787 -16360 149822 -16326
rect 149883 -16360 149918 -16326
rect 149979 -16360 150014 -16326
rect 150075 -16360 150110 -16326
rect 150171 -16360 150206 -16326
rect 150267 -16360 150302 -16326
rect 150363 -16360 150398 -16326
rect 151691 -16333 151692 -16322
rect 151868 -16327 151931 -16293
rect 151940 -16327 151975 -16293
rect 152052 -16327 152087 -16293
rect 152583 -16317 152618 -16283
rect 152679 -16317 152714 -16283
rect 152775 -16317 152810 -16283
rect 152871 -16317 152906 -16283
rect 152967 -16317 153002 -16283
rect 153992 -16324 154027 -16290
rect 154037 -16324 154038 -16279
rect 154137 -16290 154138 -16279
rect 154148 -16324 154183 -16290
rect 154193 -16324 154194 -16279
rect 154293 -16290 154294 -16279
rect 154472 -16284 154507 -16250
rect 154544 -16284 154579 -16250
rect 154616 -16284 154651 -16250
rect 154760 -16284 154795 -16250
rect 154832 -16284 154867 -16250
rect 154869 -16284 154939 -16250
rect 154976 -16284 155011 -16250
rect 155046 -16284 155081 -16250
rect 155573 -16274 155608 -16240
rect 155669 -16274 155704 -16240
rect 155765 -16274 155800 -16240
rect 157272 -16241 157307 -16207
rect 157336 -16241 157379 -16207
rect 157381 -16241 157382 -16199
rect 157481 -16207 157482 -16199
rect 157416 -16241 157451 -16207
rect 157492 -16241 157527 -16207
rect 157537 -16241 157538 -16199
rect 157637 -16207 157638 -16199
rect 157586 -16241 157621 -16207
rect 157648 -16241 157693 -16207
rect 158563 -16231 158598 -16197
rect 158659 -16231 158694 -16197
rect 158755 -16231 158790 -16197
rect 158379 -16250 158380 -16242
rect 154304 -16324 154339 -16290
rect 155285 -16293 155286 -16285
rect 155385 -16293 155386 -16285
rect 148708 -16410 148743 -16376
rect 145364 -16494 145399 -16460
rect 142374 -16620 142409 -16586
rect 143653 -16589 143654 -16578
rect 140903 -16689 140904 -16681
rect 140914 -16723 140949 -16689
rect 141134 -16734 141169 -16700
rect 139581 -16793 139616 -16759
rect 139784 -16838 139819 -16804
rect 139907 -16809 139908 -16767
rect 140229 -16796 140264 -16762
rect 139551 -16861 139552 -16853
rect 139562 -16895 139597 -16861
rect 139784 -16906 139819 -16872
rect 139551 -16961 139552 -16950
rect 139562 -16995 139597 -16961
rect 138499 -17045 138534 -17011
rect 138595 -17045 138630 -17011
rect 138691 -17045 138726 -17011
rect 139200 -17035 139235 -17001
rect 139272 -17035 139307 -17001
rect 139344 -17035 139379 -17001
rect 139416 -17029 139452 -17001
rect 139762 -17025 139797 -16991
rect 139807 -17025 139808 -16980
rect 139416 -17035 139451 -17029
rect 138853 -17088 138888 -17054
rect 138949 -17088 138984 -17054
rect 139045 -17088 139080 -17054
rect 139949 -17076 139950 -16809
rect 140578 -16819 140965 -16753
rect 139965 -16860 140000 -16826
rect 140314 -16832 140325 -16819
rect 140248 -16874 140325 -16832
rect 140376 -16874 140965 -16819
rect 141112 -16853 141147 -16819
rect 141157 -16853 141158 -16808
rect 140248 -16877 140965 -16874
rect 139965 -16928 140000 -16894
rect 140168 -16942 140203 -16908
rect 140213 -16942 140214 -16900
rect 140049 -16991 140050 -16980
rect 140060 -17025 140095 -16991
rect 140168 -17042 140203 -17008
rect 140213 -17042 140214 -16997
rect 140061 -17078 140096 -17044
rect 140133 -17078 140168 -17044
rect 140205 -17078 140240 -17044
rect 139207 -17131 139242 -17097
rect 139303 -17131 139338 -17097
rect 139399 -17131 139434 -17097
rect 139495 -17131 139530 -17097
rect 139591 -17131 139626 -17097
rect 140248 -17114 140393 -16877
rect 140578 -16899 140965 -16877
rect 140502 -16925 140965 -16899
rect 141299 -16904 141300 -16637
rect 141315 -16688 141350 -16654
rect 141929 -16691 141964 -16657
rect 142608 -16663 142643 -16629
rect 142653 -16663 142654 -16618
rect 142753 -16629 142754 -16618
rect 142764 -16663 142799 -16629
rect 142809 -16663 142810 -16618
rect 142909 -16629 142910 -16618
rect 143487 -16623 143522 -16589
rect 143664 -16623 143699 -16589
rect 144025 -16605 144060 -16571
rect 142920 -16663 142955 -16629
rect 142753 -16697 142754 -16671
rect 143152 -16689 143187 -16655
rect 143197 -16689 143198 -16644
rect 143297 -16655 143298 -16644
rect 143308 -16689 143343 -16655
rect 143353 -16689 143354 -16644
rect 143653 -16672 143654 -16661
rect 141315 -16756 141350 -16722
rect 141518 -16770 141553 -16736
rect 141563 -16770 141564 -16728
rect 141663 -16740 141664 -16729
rect 142283 -16734 142318 -16700
rect 141674 -16774 141709 -16740
rect 141399 -16819 141400 -16808
rect 141868 -16813 141903 -16779
rect 141913 -16813 141914 -16771
rect 142013 -16779 142014 -16771
rect 142673 -16777 142708 -16743
rect 142024 -16813 142059 -16779
rect 141410 -16853 141445 -16819
rect 141518 -16870 141553 -16836
rect 141563 -16870 141564 -16825
rect 141663 -16832 141664 -16821
rect 141674 -16866 141709 -16832
rect 142222 -16856 142257 -16822
rect 142267 -16856 142268 -16814
rect 142367 -16822 142368 -16814
rect 142378 -16856 142413 -16822
rect 141411 -16906 141446 -16872
rect 141483 -16906 141518 -16872
rect 141555 -16906 141590 -16872
rect 141868 -16913 141903 -16879
rect 141913 -16913 141914 -16868
rect 142013 -16879 142014 -16868
rect 142024 -16913 142059 -16879
rect 142608 -16895 142643 -16861
rect 142653 -16895 142654 -16853
rect 140502 -16959 140978 -16925
rect 141836 -16949 141871 -16915
rect 141908 -16949 141943 -16915
rect 142222 -16956 142257 -16922
rect 142267 -16956 142268 -16911
rect 142367 -16922 142368 -16911
rect 142378 -16956 142413 -16922
rect 140502 -16985 140965 -16959
rect 140506 -16993 140707 -16985
rect 140522 -17003 140691 -16993
rect 140248 -17140 140423 -17114
rect 139755 -17174 139790 -17140
rect 139851 -17174 139886 -17140
rect 139947 -17174 139982 -17140
rect 140043 -17174 140078 -17140
rect 140139 -17174 140174 -17140
rect 140235 -17174 140423 -17140
rect 140248 -17200 140423 -17174
rect 140448 -17174 140549 -17050
rect 140326 -17870 140361 -17200
rect 140448 -17228 140451 -17174
rect 140133 -17936 140278 -17924
rect 139801 -17970 140278 -17936
rect 140133 -17971 140278 -17970
rect 140314 -17971 140361 -17870
rect 140460 -17971 140495 -17174
rect 140718 -17971 140753 -17062
rect 140852 -17971 140887 -16985
rect 141105 -17002 141140 -16968
rect 141201 -17002 141236 -16968
rect 141297 -17002 141332 -16968
rect 141393 -17002 141428 -16968
rect 141489 -17002 141524 -16968
rect 141585 -17002 141620 -16968
rect 141681 -17002 141716 -16968
rect 142190 -16992 142225 -16958
rect 142262 -16992 142297 -16958
rect 142608 -16995 142643 -16961
rect 142653 -16995 142654 -16950
rect 142795 -17001 142796 -16697
rect 143487 -16706 143522 -16672
rect 143664 -16706 143699 -16672
rect 143960 -16723 143995 -16689
rect 144005 -16723 144006 -16681
rect 144147 -16753 144148 -16525
rect 144837 -16534 144872 -16500
rect 145014 -16534 145049 -16500
rect 145208 -16577 145243 -16543
rect 145253 -16577 145254 -16532
rect 145353 -16543 145354 -16532
rect 145562 -16537 145597 -16503
rect 145607 -16537 145608 -16492
rect 145707 -16503 145708 -16492
rect 145952 -16496 145987 -16462
rect 145997 -16496 145998 -16451
rect 146097 -16462 146098 -16451
rect 146108 -16496 146143 -16462
rect 146153 -16496 146154 -16451
rect 146253 -16462 146254 -16451
rect 146434 -16456 146469 -16422
rect 146506 -16456 146541 -16422
rect 146578 -16456 146613 -16422
rect 146722 -16456 146757 -16422
rect 146794 -16456 146829 -16422
rect 146831 -16456 146901 -16422
rect 146938 -16456 146973 -16422
rect 147008 -16456 147043 -16422
rect 146264 -16496 146299 -16462
rect 147304 -16491 147339 -16457
rect 147349 -16491 147350 -16446
rect 147449 -16457 147450 -16446
rect 147460 -16491 147495 -16457
rect 147505 -16491 147506 -16446
rect 147605 -16457 147606 -16446
rect 148181 -16451 148216 -16417
rect 148358 -16451 148393 -16417
rect 147616 -16491 147651 -16457
rect 145718 -16537 145753 -16503
rect 146997 -16505 146998 -16494
rect 145364 -16577 145399 -16543
rect 144277 -16621 144312 -16587
rect 144478 -16666 144513 -16632
rect 144601 -16637 144602 -16595
rect 144923 -16624 144958 -16590
rect 145562 -16620 145597 -16586
rect 145607 -16620 145608 -16575
rect 145707 -16586 145708 -16575
rect 145952 -16580 145987 -16546
rect 145997 -16580 145998 -16535
rect 146097 -16546 146098 -16535
rect 146108 -16580 146143 -16546
rect 146153 -16580 146154 -16535
rect 146253 -16546 146254 -16535
rect 146831 -16539 146866 -16505
rect 147008 -16539 147043 -16505
rect 146264 -16580 146299 -16546
rect 147151 -16565 147266 -16499
rect 147449 -16525 147450 -16499
rect 147846 -16517 147881 -16483
rect 147891 -16517 147892 -16472
rect 147991 -16483 147992 -16472
rect 148002 -16517 148037 -16483
rect 148047 -16517 148048 -16472
rect 148347 -16500 148348 -16489
rect 148552 -16494 148587 -16460
rect 148597 -16494 148598 -16449
rect 148697 -16460 148698 -16449
rect 148906 -16453 148941 -16419
rect 148951 -16453 148952 -16408
rect 149051 -16419 149052 -16408
rect 149232 -16413 149267 -16379
rect 149296 -16413 149339 -16379
rect 149341 -16413 149342 -16371
rect 149441 -16379 149442 -16371
rect 149376 -16413 149411 -16379
rect 149452 -16413 149487 -16379
rect 149497 -16413 149498 -16371
rect 149597 -16379 149598 -16371
rect 149546 -16413 149581 -16379
rect 149608 -16413 149653 -16379
rect 150648 -16408 150683 -16374
rect 150693 -16408 150694 -16363
rect 150793 -16374 150794 -16363
rect 150804 -16408 150839 -16374
rect 150849 -16408 150850 -16363
rect 150949 -16374 150950 -16363
rect 151525 -16367 151560 -16333
rect 151702 -16367 151737 -16333
rect 152295 -16336 152296 -16328
rect 152395 -16336 152396 -16328
rect 150960 -16408 150995 -16374
rect 149062 -16453 149097 -16419
rect 150341 -16422 150342 -16414
rect 151691 -16417 151692 -16406
rect 151896 -16410 151931 -16376
rect 151941 -16410 151942 -16365
rect 152041 -16376 152042 -16365
rect 152222 -16370 152285 -16336
rect 152294 -16370 152329 -16336
rect 152406 -16370 152441 -16336
rect 153131 -16360 153166 -16326
rect 153227 -16360 153262 -16326
rect 153323 -16360 153358 -16326
rect 153419 -16360 153454 -16326
rect 153515 -16360 153550 -16326
rect 153611 -16360 153646 -16326
rect 153707 -16360 153742 -16326
rect 155035 -16333 155036 -16322
rect 155212 -16327 155275 -16293
rect 155284 -16327 155319 -16293
rect 155396 -16327 155431 -16293
rect 155927 -16317 155962 -16283
rect 156023 -16317 156058 -16283
rect 156119 -16317 156154 -16283
rect 156215 -16317 156250 -16283
rect 156311 -16317 156346 -16283
rect 157336 -16324 157371 -16290
rect 157381 -16324 157382 -16279
rect 157481 -16290 157482 -16279
rect 157492 -16324 157527 -16290
rect 157537 -16324 157538 -16279
rect 157637 -16290 157638 -16279
rect 157816 -16284 157851 -16250
rect 157888 -16284 157923 -16250
rect 157960 -16284 157995 -16250
rect 158104 -16284 158139 -16250
rect 158176 -16284 158211 -16250
rect 158213 -16284 158283 -16250
rect 158320 -16284 158355 -16250
rect 158390 -16284 158425 -16250
rect 158917 -16274 158952 -16240
rect 159013 -16274 159048 -16240
rect 159109 -16274 159144 -16240
rect 160616 -16241 160651 -16207
rect 160680 -16241 160723 -16207
rect 160725 -16241 160726 -16199
rect 160825 -16207 160826 -16199
rect 160760 -16241 160795 -16207
rect 160836 -16241 160871 -16207
rect 160881 -16241 160882 -16199
rect 160981 -16207 160982 -16199
rect 160930 -16241 160965 -16207
rect 160992 -16241 161037 -16207
rect 161907 -16231 161942 -16197
rect 162003 -16231 162038 -16197
rect 162099 -16231 162134 -16197
rect 161723 -16250 161724 -16242
rect 157648 -16324 157683 -16290
rect 158629 -16293 158630 -16285
rect 158729 -16293 158730 -16285
rect 152052 -16410 152087 -16376
rect 148708 -16494 148743 -16460
rect 145718 -16620 145753 -16586
rect 146997 -16589 146998 -16578
rect 144247 -16689 144248 -16681
rect 144258 -16723 144293 -16689
rect 144478 -16734 144513 -16700
rect 142925 -16793 142960 -16759
rect 143128 -16838 143163 -16804
rect 143251 -16809 143252 -16767
rect 143573 -16796 143608 -16762
rect 142895 -16861 142896 -16853
rect 142906 -16895 142941 -16861
rect 143128 -16906 143163 -16872
rect 142895 -16961 142896 -16950
rect 142906 -16995 142941 -16961
rect 141843 -17045 141878 -17011
rect 141939 -17045 141974 -17011
rect 142035 -17045 142070 -17011
rect 142544 -17035 142579 -17001
rect 142616 -17035 142651 -17001
rect 142688 -17035 142723 -17001
rect 142760 -17029 142796 -17001
rect 143106 -17025 143141 -16991
rect 143151 -17025 143152 -16980
rect 142760 -17035 142795 -17029
rect 142197 -17088 142232 -17054
rect 142293 -17088 142328 -17054
rect 142389 -17088 142424 -17054
rect 143293 -17076 143294 -16809
rect 143922 -16819 144309 -16753
rect 143309 -16860 143344 -16826
rect 143658 -16832 143669 -16819
rect 143592 -16874 143669 -16832
rect 143720 -16874 144309 -16819
rect 144456 -16853 144491 -16819
rect 144501 -16853 144502 -16808
rect 143592 -16877 144309 -16874
rect 143309 -16928 143344 -16894
rect 143512 -16942 143547 -16908
rect 143557 -16942 143558 -16900
rect 143393 -16991 143394 -16980
rect 143404 -17025 143439 -16991
rect 143512 -17042 143547 -17008
rect 143557 -17042 143558 -16997
rect 143405 -17078 143440 -17044
rect 143477 -17078 143512 -17044
rect 143549 -17078 143584 -17044
rect 142551 -17131 142586 -17097
rect 142647 -17131 142682 -17097
rect 142743 -17131 142778 -17097
rect 142839 -17131 142874 -17097
rect 142935 -17131 142970 -17097
rect 143592 -17114 143737 -16877
rect 143922 -16899 144309 -16877
rect 143846 -16925 144309 -16899
rect 144643 -16904 144644 -16637
rect 144659 -16688 144694 -16654
rect 145273 -16691 145308 -16657
rect 145952 -16663 145987 -16629
rect 145997 -16663 145998 -16618
rect 146097 -16629 146098 -16618
rect 146108 -16663 146143 -16629
rect 146153 -16663 146154 -16618
rect 146253 -16629 146254 -16618
rect 146831 -16623 146866 -16589
rect 147008 -16623 147043 -16589
rect 147369 -16605 147404 -16571
rect 146264 -16663 146299 -16629
rect 146097 -16697 146098 -16671
rect 146496 -16689 146531 -16655
rect 146541 -16689 146542 -16644
rect 146641 -16655 146642 -16644
rect 146652 -16689 146687 -16655
rect 146697 -16689 146698 -16644
rect 146997 -16672 146998 -16661
rect 144659 -16756 144694 -16722
rect 144862 -16770 144897 -16736
rect 144907 -16770 144908 -16728
rect 145007 -16740 145008 -16729
rect 145627 -16734 145662 -16700
rect 145018 -16774 145053 -16740
rect 144743 -16819 144744 -16808
rect 145212 -16813 145247 -16779
rect 145257 -16813 145258 -16771
rect 145357 -16779 145358 -16771
rect 146017 -16777 146052 -16743
rect 145368 -16813 145403 -16779
rect 144754 -16853 144789 -16819
rect 144862 -16870 144897 -16836
rect 144907 -16870 144908 -16825
rect 145007 -16832 145008 -16821
rect 145018 -16866 145053 -16832
rect 145566 -16856 145601 -16822
rect 145611 -16856 145612 -16814
rect 145711 -16822 145712 -16814
rect 145722 -16856 145757 -16822
rect 144755 -16906 144790 -16872
rect 144827 -16906 144862 -16872
rect 144899 -16906 144934 -16872
rect 145212 -16913 145247 -16879
rect 145257 -16913 145258 -16868
rect 145357 -16879 145358 -16868
rect 145368 -16913 145403 -16879
rect 145952 -16895 145987 -16861
rect 145997 -16895 145998 -16853
rect 143846 -16959 144322 -16925
rect 145180 -16949 145215 -16915
rect 145252 -16949 145287 -16915
rect 145566 -16956 145601 -16922
rect 145611 -16956 145612 -16911
rect 145711 -16922 145712 -16911
rect 145722 -16956 145757 -16922
rect 143846 -16985 144309 -16959
rect 143850 -16993 144051 -16985
rect 143866 -17003 144035 -16993
rect 143592 -17140 143767 -17114
rect 143099 -17174 143134 -17140
rect 143195 -17174 143230 -17140
rect 143291 -17174 143326 -17140
rect 143387 -17174 143422 -17140
rect 143483 -17174 143518 -17140
rect 143579 -17174 143767 -17140
rect 143592 -17200 143767 -17174
rect 143792 -17174 143893 -17050
rect 143670 -17870 143705 -17200
rect 143792 -17228 143795 -17174
rect 143477 -17936 143622 -17924
rect 143145 -17970 143622 -17936
rect 143477 -17971 143622 -17970
rect 143658 -17971 143705 -17870
rect 143804 -17971 143839 -17174
rect 144062 -17971 144097 -17062
rect 144196 -17971 144231 -16985
rect 144449 -17002 144484 -16968
rect 144545 -17002 144580 -16968
rect 144641 -17002 144676 -16968
rect 144737 -17002 144772 -16968
rect 144833 -17002 144868 -16968
rect 144929 -17002 144964 -16968
rect 145025 -17002 145060 -16968
rect 145534 -16992 145569 -16958
rect 145606 -16992 145641 -16958
rect 145952 -16995 145987 -16961
rect 145997 -16995 145998 -16950
rect 146139 -17001 146140 -16697
rect 146831 -16706 146866 -16672
rect 147008 -16706 147043 -16672
rect 147304 -16723 147339 -16689
rect 147349 -16723 147350 -16681
rect 147491 -16753 147492 -16525
rect 148181 -16534 148216 -16500
rect 148358 -16534 148393 -16500
rect 148552 -16577 148587 -16543
rect 148597 -16577 148598 -16532
rect 148697 -16543 148698 -16532
rect 148906 -16537 148941 -16503
rect 148951 -16537 148952 -16492
rect 149051 -16503 149052 -16492
rect 149296 -16496 149331 -16462
rect 149341 -16496 149342 -16451
rect 149441 -16462 149442 -16451
rect 149452 -16496 149487 -16462
rect 149497 -16496 149498 -16451
rect 149597 -16462 149598 -16451
rect 149778 -16456 149813 -16422
rect 149850 -16456 149885 -16422
rect 149922 -16456 149957 -16422
rect 150066 -16456 150101 -16422
rect 150138 -16456 150173 -16422
rect 150175 -16456 150245 -16422
rect 150282 -16456 150317 -16422
rect 150352 -16456 150387 -16422
rect 149608 -16496 149643 -16462
rect 150648 -16491 150683 -16457
rect 150693 -16491 150694 -16446
rect 150793 -16457 150794 -16446
rect 150804 -16491 150839 -16457
rect 150849 -16491 150850 -16446
rect 150949 -16457 150950 -16446
rect 151525 -16451 151560 -16417
rect 151702 -16451 151737 -16417
rect 150960 -16491 150995 -16457
rect 149062 -16537 149097 -16503
rect 150341 -16505 150342 -16494
rect 148708 -16577 148743 -16543
rect 147621 -16621 147656 -16587
rect 147822 -16666 147857 -16632
rect 147945 -16637 147946 -16595
rect 148267 -16624 148302 -16590
rect 148906 -16620 148941 -16586
rect 148951 -16620 148952 -16575
rect 149051 -16586 149052 -16575
rect 149296 -16580 149331 -16546
rect 149341 -16580 149342 -16535
rect 149441 -16546 149442 -16535
rect 149452 -16580 149487 -16546
rect 149497 -16580 149498 -16535
rect 149597 -16546 149598 -16535
rect 150175 -16539 150210 -16505
rect 150352 -16539 150387 -16505
rect 149608 -16580 149643 -16546
rect 150495 -16565 150610 -16499
rect 150793 -16525 150794 -16499
rect 151190 -16517 151225 -16483
rect 151235 -16517 151236 -16472
rect 151335 -16483 151336 -16472
rect 151346 -16517 151381 -16483
rect 151391 -16517 151392 -16472
rect 151691 -16500 151692 -16489
rect 151896 -16494 151931 -16460
rect 151941 -16494 151942 -16449
rect 152041 -16460 152042 -16449
rect 152250 -16453 152285 -16419
rect 152295 -16453 152296 -16408
rect 152395 -16419 152396 -16408
rect 152576 -16413 152611 -16379
rect 152640 -16413 152683 -16379
rect 152685 -16413 152686 -16371
rect 152785 -16379 152786 -16371
rect 152720 -16413 152755 -16379
rect 152796 -16413 152831 -16379
rect 152841 -16413 152842 -16371
rect 152941 -16379 152942 -16371
rect 152890 -16413 152925 -16379
rect 152952 -16413 152997 -16379
rect 153992 -16408 154027 -16374
rect 154037 -16408 154038 -16363
rect 154137 -16374 154138 -16363
rect 154148 -16408 154183 -16374
rect 154193 -16408 154194 -16363
rect 154293 -16374 154294 -16363
rect 154869 -16367 154904 -16333
rect 155046 -16367 155081 -16333
rect 155639 -16336 155640 -16328
rect 155739 -16336 155740 -16328
rect 154304 -16408 154339 -16374
rect 152406 -16453 152441 -16419
rect 153685 -16422 153686 -16414
rect 155035 -16417 155036 -16406
rect 155240 -16410 155275 -16376
rect 155285 -16410 155286 -16365
rect 155385 -16376 155386 -16365
rect 155566 -16370 155629 -16336
rect 155638 -16370 155673 -16336
rect 155750 -16370 155785 -16336
rect 156475 -16360 156510 -16326
rect 156571 -16360 156606 -16326
rect 156667 -16360 156702 -16326
rect 156763 -16360 156798 -16326
rect 156859 -16360 156894 -16326
rect 156955 -16360 156990 -16326
rect 157051 -16360 157086 -16326
rect 158379 -16333 158380 -16322
rect 158556 -16327 158619 -16293
rect 158628 -16327 158663 -16293
rect 158740 -16327 158775 -16293
rect 159271 -16317 159306 -16283
rect 159367 -16317 159402 -16283
rect 159463 -16317 159498 -16283
rect 159559 -16317 159594 -16283
rect 159655 -16317 159690 -16283
rect 160680 -16324 160715 -16290
rect 160725 -16324 160726 -16279
rect 160825 -16290 160826 -16279
rect 160836 -16324 160871 -16290
rect 160881 -16324 160882 -16279
rect 160981 -16290 160982 -16279
rect 161160 -16284 161195 -16250
rect 161232 -16284 161267 -16250
rect 161304 -16284 161339 -16250
rect 161448 -16284 161483 -16250
rect 161520 -16284 161555 -16250
rect 161557 -16284 161627 -16250
rect 161664 -16284 161699 -16250
rect 161734 -16284 161769 -16250
rect 162261 -16274 162296 -16240
rect 162357 -16274 162392 -16240
rect 162453 -16274 162488 -16240
rect 163960 -16241 163995 -16207
rect 164024 -16241 164067 -16207
rect 164069 -16241 164070 -16199
rect 164169 -16207 164170 -16199
rect 164104 -16241 164139 -16207
rect 164180 -16241 164215 -16207
rect 164225 -16241 164226 -16199
rect 164325 -16207 164326 -16199
rect 164274 -16241 164309 -16207
rect 164336 -16241 164381 -16207
rect 165251 -16231 165286 -16197
rect 165347 -16231 165382 -16197
rect 165443 -16231 165478 -16197
rect 165067 -16250 165068 -16242
rect 160992 -16324 161027 -16290
rect 161973 -16293 161974 -16285
rect 162073 -16293 162074 -16285
rect 155396 -16410 155431 -16376
rect 152052 -16494 152087 -16460
rect 149062 -16620 149097 -16586
rect 150341 -16589 150342 -16578
rect 147591 -16689 147592 -16681
rect 147602 -16723 147637 -16689
rect 147822 -16734 147857 -16700
rect 146269 -16793 146304 -16759
rect 146472 -16838 146507 -16804
rect 146595 -16809 146596 -16767
rect 146917 -16796 146952 -16762
rect 146239 -16861 146240 -16853
rect 146250 -16895 146285 -16861
rect 146472 -16906 146507 -16872
rect 146239 -16961 146240 -16950
rect 146250 -16995 146285 -16961
rect 145187 -17045 145222 -17011
rect 145283 -17045 145318 -17011
rect 145379 -17045 145414 -17011
rect 145888 -17035 145923 -17001
rect 145960 -17035 145995 -17001
rect 146032 -17035 146067 -17001
rect 146104 -17029 146140 -17001
rect 146450 -17025 146485 -16991
rect 146495 -17025 146496 -16980
rect 146104 -17035 146139 -17029
rect 145541 -17088 145576 -17054
rect 145637 -17088 145672 -17054
rect 145733 -17088 145768 -17054
rect 146637 -17076 146638 -16809
rect 147266 -16819 147653 -16753
rect 146653 -16860 146688 -16826
rect 147002 -16832 147013 -16819
rect 146936 -16874 147013 -16832
rect 147064 -16874 147653 -16819
rect 147800 -16853 147835 -16819
rect 147845 -16853 147846 -16808
rect 146936 -16877 147653 -16874
rect 146653 -16928 146688 -16894
rect 146856 -16942 146891 -16908
rect 146901 -16942 146902 -16900
rect 146737 -16991 146738 -16980
rect 146748 -17025 146783 -16991
rect 146856 -17042 146891 -17008
rect 146901 -17042 146902 -16997
rect 146749 -17078 146784 -17044
rect 146821 -17078 146856 -17044
rect 146893 -17078 146928 -17044
rect 145895 -17131 145930 -17097
rect 145991 -17131 146026 -17097
rect 146087 -17131 146122 -17097
rect 146183 -17131 146218 -17097
rect 146279 -17131 146314 -17097
rect 146936 -17114 147081 -16877
rect 147266 -16899 147653 -16877
rect 147190 -16925 147653 -16899
rect 147987 -16904 147988 -16637
rect 148003 -16688 148038 -16654
rect 148617 -16691 148652 -16657
rect 149296 -16663 149331 -16629
rect 149341 -16663 149342 -16618
rect 149441 -16629 149442 -16618
rect 149452 -16663 149487 -16629
rect 149497 -16663 149498 -16618
rect 149597 -16629 149598 -16618
rect 150175 -16623 150210 -16589
rect 150352 -16623 150387 -16589
rect 150713 -16605 150748 -16571
rect 149608 -16663 149643 -16629
rect 149441 -16697 149442 -16671
rect 149840 -16689 149875 -16655
rect 149885 -16689 149886 -16644
rect 149985 -16655 149986 -16644
rect 149996 -16689 150031 -16655
rect 150041 -16689 150042 -16644
rect 150341 -16672 150342 -16661
rect 148003 -16756 148038 -16722
rect 148206 -16770 148241 -16736
rect 148251 -16770 148252 -16728
rect 148351 -16740 148352 -16729
rect 148971 -16734 149006 -16700
rect 148362 -16774 148397 -16740
rect 148087 -16819 148088 -16808
rect 148556 -16813 148591 -16779
rect 148601 -16813 148602 -16771
rect 148701 -16779 148702 -16771
rect 149361 -16777 149396 -16743
rect 148712 -16813 148747 -16779
rect 148098 -16853 148133 -16819
rect 148206 -16870 148241 -16836
rect 148251 -16870 148252 -16825
rect 148351 -16832 148352 -16821
rect 148362 -16866 148397 -16832
rect 148910 -16856 148945 -16822
rect 148955 -16856 148956 -16814
rect 149055 -16822 149056 -16814
rect 149066 -16856 149101 -16822
rect 148099 -16906 148134 -16872
rect 148171 -16906 148206 -16872
rect 148243 -16906 148278 -16872
rect 148556 -16913 148591 -16879
rect 148601 -16913 148602 -16868
rect 148701 -16879 148702 -16868
rect 148712 -16913 148747 -16879
rect 149296 -16895 149331 -16861
rect 149341 -16895 149342 -16853
rect 147190 -16959 147666 -16925
rect 148524 -16949 148559 -16915
rect 148596 -16949 148631 -16915
rect 148910 -16956 148945 -16922
rect 148955 -16956 148956 -16911
rect 149055 -16922 149056 -16911
rect 149066 -16956 149101 -16922
rect 147190 -16985 147653 -16959
rect 147194 -16993 147395 -16985
rect 147210 -17003 147379 -16993
rect 146936 -17140 147111 -17114
rect 146443 -17174 146478 -17140
rect 146539 -17174 146574 -17140
rect 146635 -17174 146670 -17140
rect 146731 -17174 146766 -17140
rect 146827 -17174 146862 -17140
rect 146923 -17174 147111 -17140
rect 146936 -17200 147111 -17174
rect 147136 -17174 147237 -17050
rect 147014 -17870 147049 -17200
rect 147136 -17228 147139 -17174
rect 146821 -17936 146966 -17924
rect 146489 -17970 146966 -17936
rect 146821 -17971 146966 -17970
rect 147002 -17971 147049 -17870
rect 147148 -17971 147183 -17174
rect 147406 -17971 147441 -17062
rect 147540 -17971 147575 -16985
rect 147793 -17002 147828 -16968
rect 147889 -17002 147924 -16968
rect 147985 -17002 148020 -16968
rect 148081 -17002 148116 -16968
rect 148177 -17002 148212 -16968
rect 148273 -17002 148308 -16968
rect 148369 -17002 148404 -16968
rect 148878 -16992 148913 -16958
rect 148950 -16992 148985 -16958
rect 149296 -16995 149331 -16961
rect 149341 -16995 149342 -16950
rect 149483 -17001 149484 -16697
rect 150175 -16706 150210 -16672
rect 150352 -16706 150387 -16672
rect 150648 -16723 150683 -16689
rect 150693 -16723 150694 -16681
rect 150835 -16753 150836 -16525
rect 151525 -16534 151560 -16500
rect 151702 -16534 151737 -16500
rect 151896 -16577 151931 -16543
rect 151941 -16577 151942 -16532
rect 152041 -16543 152042 -16532
rect 152250 -16537 152285 -16503
rect 152295 -16537 152296 -16492
rect 152395 -16503 152396 -16492
rect 152640 -16496 152675 -16462
rect 152685 -16496 152686 -16451
rect 152785 -16462 152786 -16451
rect 152796 -16496 152831 -16462
rect 152841 -16496 152842 -16451
rect 152941 -16462 152942 -16451
rect 153122 -16456 153157 -16422
rect 153194 -16456 153229 -16422
rect 153266 -16456 153301 -16422
rect 153410 -16456 153445 -16422
rect 153482 -16456 153517 -16422
rect 153519 -16456 153589 -16422
rect 153626 -16456 153661 -16422
rect 153696 -16456 153731 -16422
rect 152952 -16496 152987 -16462
rect 153992 -16491 154027 -16457
rect 154037 -16491 154038 -16446
rect 154137 -16457 154138 -16446
rect 154148 -16491 154183 -16457
rect 154193 -16491 154194 -16446
rect 154293 -16457 154294 -16446
rect 154869 -16451 154904 -16417
rect 155046 -16451 155081 -16417
rect 154304 -16491 154339 -16457
rect 152406 -16537 152441 -16503
rect 153685 -16505 153686 -16494
rect 152052 -16577 152087 -16543
rect 150965 -16621 151000 -16587
rect 151166 -16666 151201 -16632
rect 151289 -16637 151290 -16595
rect 151611 -16624 151646 -16590
rect 152250 -16620 152285 -16586
rect 152295 -16620 152296 -16575
rect 152395 -16586 152396 -16575
rect 152640 -16580 152675 -16546
rect 152685 -16580 152686 -16535
rect 152785 -16546 152786 -16535
rect 152796 -16580 152831 -16546
rect 152841 -16580 152842 -16535
rect 152941 -16546 152942 -16535
rect 153519 -16539 153554 -16505
rect 153696 -16539 153731 -16505
rect 152952 -16580 152987 -16546
rect 153839 -16565 153954 -16499
rect 154137 -16525 154138 -16499
rect 154534 -16517 154569 -16483
rect 154579 -16517 154580 -16472
rect 154679 -16483 154680 -16472
rect 154690 -16517 154725 -16483
rect 154735 -16517 154736 -16472
rect 155035 -16500 155036 -16489
rect 155240 -16494 155275 -16460
rect 155285 -16494 155286 -16449
rect 155385 -16460 155386 -16449
rect 155594 -16453 155629 -16419
rect 155639 -16453 155640 -16408
rect 155739 -16419 155740 -16408
rect 155920 -16413 155955 -16379
rect 155984 -16413 156027 -16379
rect 156029 -16413 156030 -16371
rect 156129 -16379 156130 -16371
rect 156064 -16413 156099 -16379
rect 156140 -16413 156175 -16379
rect 156185 -16413 156186 -16371
rect 156285 -16379 156286 -16371
rect 156234 -16413 156269 -16379
rect 156296 -16413 156341 -16379
rect 157336 -16408 157371 -16374
rect 157381 -16408 157382 -16363
rect 157481 -16374 157482 -16363
rect 157492 -16408 157527 -16374
rect 157537 -16408 157538 -16363
rect 157637 -16374 157638 -16363
rect 158213 -16367 158248 -16333
rect 158390 -16367 158425 -16333
rect 158983 -16336 158984 -16328
rect 159083 -16336 159084 -16328
rect 157648 -16408 157683 -16374
rect 155750 -16453 155785 -16419
rect 157029 -16422 157030 -16414
rect 158379 -16417 158380 -16406
rect 158584 -16410 158619 -16376
rect 158629 -16410 158630 -16365
rect 158729 -16376 158730 -16365
rect 158910 -16370 158973 -16336
rect 158982 -16370 159017 -16336
rect 159094 -16370 159129 -16336
rect 159819 -16360 159854 -16326
rect 159915 -16360 159950 -16326
rect 160011 -16360 160046 -16326
rect 160107 -16360 160142 -16326
rect 160203 -16360 160238 -16326
rect 160299 -16360 160334 -16326
rect 160395 -16360 160430 -16326
rect 161723 -16333 161724 -16322
rect 161900 -16327 161963 -16293
rect 161972 -16327 162007 -16293
rect 162084 -16327 162119 -16293
rect 162615 -16317 162650 -16283
rect 162711 -16317 162746 -16283
rect 162807 -16317 162842 -16283
rect 162903 -16317 162938 -16283
rect 162999 -16317 163034 -16283
rect 164024 -16324 164059 -16290
rect 164069 -16324 164070 -16279
rect 164169 -16290 164170 -16279
rect 164180 -16324 164215 -16290
rect 164225 -16324 164226 -16279
rect 164325 -16290 164326 -16279
rect 164504 -16284 164539 -16250
rect 164576 -16284 164611 -16250
rect 164648 -16284 164683 -16250
rect 164792 -16284 164827 -16250
rect 164864 -16284 164899 -16250
rect 164901 -16284 164971 -16250
rect 165008 -16284 165043 -16250
rect 165078 -16284 165113 -16250
rect 165605 -16274 165640 -16240
rect 165701 -16274 165736 -16240
rect 165797 -16274 165832 -16240
rect 167304 -16241 167339 -16207
rect 167368 -16241 167411 -16207
rect 167413 -16241 167414 -16199
rect 167513 -16207 167514 -16199
rect 167448 -16241 167483 -16207
rect 167524 -16241 167559 -16207
rect 167569 -16241 167570 -16199
rect 167669 -16207 167670 -16199
rect 167618 -16241 167653 -16207
rect 167680 -16241 167725 -16207
rect 168595 -16231 168630 -16197
rect 168691 -16231 168726 -16197
rect 168787 -16231 168822 -16197
rect 168411 -16250 168412 -16242
rect 164336 -16324 164371 -16290
rect 165317 -16293 165318 -16285
rect 165417 -16293 165418 -16285
rect 158740 -16410 158775 -16376
rect 155396 -16494 155431 -16460
rect 152406 -16620 152441 -16586
rect 153685 -16589 153686 -16578
rect 150935 -16689 150936 -16681
rect 150946 -16723 150981 -16689
rect 151166 -16734 151201 -16700
rect 149613 -16793 149648 -16759
rect 149816 -16838 149851 -16804
rect 149939 -16809 149940 -16767
rect 150261 -16796 150296 -16762
rect 149583 -16861 149584 -16853
rect 149594 -16895 149629 -16861
rect 149816 -16906 149851 -16872
rect 149583 -16961 149584 -16950
rect 149594 -16995 149629 -16961
rect 148531 -17045 148566 -17011
rect 148627 -17045 148662 -17011
rect 148723 -17045 148758 -17011
rect 149232 -17035 149267 -17001
rect 149304 -17035 149339 -17001
rect 149376 -17035 149411 -17001
rect 149448 -17029 149484 -17001
rect 149794 -17025 149829 -16991
rect 149839 -17025 149840 -16980
rect 149448 -17035 149483 -17029
rect 148885 -17088 148920 -17054
rect 148981 -17088 149016 -17054
rect 149077 -17088 149112 -17054
rect 149981 -17076 149982 -16809
rect 150610 -16819 150997 -16753
rect 149997 -16860 150032 -16826
rect 150346 -16832 150357 -16819
rect 150280 -16874 150357 -16832
rect 150408 -16874 150997 -16819
rect 151144 -16853 151179 -16819
rect 151189 -16853 151190 -16808
rect 150280 -16877 150997 -16874
rect 149997 -16928 150032 -16894
rect 150200 -16942 150235 -16908
rect 150245 -16942 150246 -16900
rect 150081 -16991 150082 -16980
rect 150092 -17025 150127 -16991
rect 150200 -17042 150235 -17008
rect 150245 -17042 150246 -16997
rect 150093 -17078 150128 -17044
rect 150165 -17078 150200 -17044
rect 150237 -17078 150272 -17044
rect 149239 -17131 149274 -17097
rect 149335 -17131 149370 -17097
rect 149431 -17131 149466 -17097
rect 149527 -17131 149562 -17097
rect 149623 -17131 149658 -17097
rect 150280 -17114 150425 -16877
rect 150610 -16899 150997 -16877
rect 150534 -16925 150997 -16899
rect 151331 -16904 151332 -16637
rect 151347 -16688 151382 -16654
rect 151961 -16691 151996 -16657
rect 152640 -16663 152675 -16629
rect 152685 -16663 152686 -16618
rect 152785 -16629 152786 -16618
rect 152796 -16663 152831 -16629
rect 152841 -16663 152842 -16618
rect 152941 -16629 152942 -16618
rect 153519 -16623 153554 -16589
rect 153696 -16623 153731 -16589
rect 154057 -16605 154092 -16571
rect 152952 -16663 152987 -16629
rect 152785 -16697 152786 -16671
rect 153184 -16689 153219 -16655
rect 153229 -16689 153230 -16644
rect 153329 -16655 153330 -16644
rect 153340 -16689 153375 -16655
rect 153385 -16689 153386 -16644
rect 153685 -16672 153686 -16661
rect 151347 -16756 151382 -16722
rect 151550 -16770 151585 -16736
rect 151595 -16770 151596 -16728
rect 151695 -16740 151696 -16729
rect 152315 -16734 152350 -16700
rect 151706 -16774 151741 -16740
rect 151431 -16819 151432 -16808
rect 151900 -16813 151935 -16779
rect 151945 -16813 151946 -16771
rect 152045 -16779 152046 -16771
rect 152705 -16777 152740 -16743
rect 152056 -16813 152091 -16779
rect 151442 -16853 151477 -16819
rect 151550 -16870 151585 -16836
rect 151595 -16870 151596 -16825
rect 151695 -16832 151696 -16821
rect 151706 -16866 151741 -16832
rect 152254 -16856 152289 -16822
rect 152299 -16856 152300 -16814
rect 152399 -16822 152400 -16814
rect 152410 -16856 152445 -16822
rect 151443 -16906 151478 -16872
rect 151515 -16906 151550 -16872
rect 151587 -16906 151622 -16872
rect 151900 -16913 151935 -16879
rect 151945 -16913 151946 -16868
rect 152045 -16879 152046 -16868
rect 152056 -16913 152091 -16879
rect 152640 -16895 152675 -16861
rect 152685 -16895 152686 -16853
rect 150534 -16959 151010 -16925
rect 151868 -16949 151903 -16915
rect 151940 -16949 151975 -16915
rect 152254 -16956 152289 -16922
rect 152299 -16956 152300 -16911
rect 152399 -16922 152400 -16911
rect 152410 -16956 152445 -16922
rect 150534 -16985 150997 -16959
rect 150538 -16993 150739 -16985
rect 150554 -17003 150723 -16993
rect 150280 -17140 150455 -17114
rect 149787 -17174 149822 -17140
rect 149883 -17174 149918 -17140
rect 149979 -17174 150014 -17140
rect 150075 -17174 150110 -17140
rect 150171 -17174 150206 -17140
rect 150267 -17174 150455 -17140
rect 150280 -17200 150455 -17174
rect 150480 -17174 150581 -17050
rect 150358 -17870 150393 -17200
rect 150480 -17228 150483 -17174
rect 150165 -17936 150310 -17924
rect 149833 -17970 150310 -17936
rect 150165 -17971 150310 -17970
rect 150346 -17971 150393 -17870
rect 150492 -17971 150527 -17174
rect 150750 -17971 150785 -17062
rect 150884 -17971 150919 -16985
rect 151137 -17002 151172 -16968
rect 151233 -17002 151268 -16968
rect 151329 -17002 151364 -16968
rect 151425 -17002 151460 -16968
rect 151521 -17002 151556 -16968
rect 151617 -17002 151652 -16968
rect 151713 -17002 151748 -16968
rect 152222 -16992 152257 -16958
rect 152294 -16992 152329 -16958
rect 152640 -16995 152675 -16961
rect 152685 -16995 152686 -16950
rect 152827 -17001 152828 -16697
rect 153519 -16706 153554 -16672
rect 153696 -16706 153731 -16672
rect 153992 -16723 154027 -16689
rect 154037 -16723 154038 -16681
rect 154179 -16753 154180 -16525
rect 154869 -16534 154904 -16500
rect 155046 -16534 155081 -16500
rect 155240 -16577 155275 -16543
rect 155285 -16577 155286 -16532
rect 155385 -16543 155386 -16532
rect 155594 -16537 155629 -16503
rect 155639 -16537 155640 -16492
rect 155739 -16503 155740 -16492
rect 155984 -16496 156019 -16462
rect 156029 -16496 156030 -16451
rect 156129 -16462 156130 -16451
rect 156140 -16496 156175 -16462
rect 156185 -16496 156186 -16451
rect 156285 -16462 156286 -16451
rect 156466 -16456 156501 -16422
rect 156538 -16456 156573 -16422
rect 156610 -16456 156645 -16422
rect 156754 -16456 156789 -16422
rect 156826 -16456 156861 -16422
rect 156863 -16456 156933 -16422
rect 156970 -16456 157005 -16422
rect 157040 -16456 157075 -16422
rect 156296 -16496 156331 -16462
rect 157336 -16491 157371 -16457
rect 157381 -16491 157382 -16446
rect 157481 -16457 157482 -16446
rect 157492 -16491 157527 -16457
rect 157537 -16491 157538 -16446
rect 157637 -16457 157638 -16446
rect 158213 -16451 158248 -16417
rect 158390 -16451 158425 -16417
rect 157648 -16491 157683 -16457
rect 155750 -16537 155785 -16503
rect 157029 -16505 157030 -16494
rect 155396 -16577 155431 -16543
rect 154309 -16621 154344 -16587
rect 154510 -16666 154545 -16632
rect 154633 -16637 154634 -16595
rect 154955 -16624 154990 -16590
rect 155594 -16620 155629 -16586
rect 155639 -16620 155640 -16575
rect 155739 -16586 155740 -16575
rect 155984 -16580 156019 -16546
rect 156029 -16580 156030 -16535
rect 156129 -16546 156130 -16535
rect 156140 -16580 156175 -16546
rect 156185 -16580 156186 -16535
rect 156285 -16546 156286 -16535
rect 156863 -16539 156898 -16505
rect 157040 -16539 157075 -16505
rect 156296 -16580 156331 -16546
rect 157183 -16565 157298 -16499
rect 157481 -16525 157482 -16499
rect 157878 -16517 157913 -16483
rect 157923 -16517 157924 -16472
rect 158023 -16483 158024 -16472
rect 158034 -16517 158069 -16483
rect 158079 -16517 158080 -16472
rect 158379 -16500 158380 -16489
rect 158584 -16494 158619 -16460
rect 158629 -16494 158630 -16449
rect 158729 -16460 158730 -16449
rect 158938 -16453 158973 -16419
rect 158983 -16453 158984 -16408
rect 159083 -16419 159084 -16408
rect 159264 -16413 159299 -16379
rect 159328 -16413 159371 -16379
rect 159373 -16413 159374 -16371
rect 159473 -16379 159474 -16371
rect 159408 -16413 159443 -16379
rect 159484 -16413 159519 -16379
rect 159529 -16413 159530 -16371
rect 159629 -16379 159630 -16371
rect 159578 -16413 159613 -16379
rect 159640 -16413 159685 -16379
rect 160680 -16408 160715 -16374
rect 160725 -16408 160726 -16363
rect 160825 -16374 160826 -16363
rect 160836 -16408 160871 -16374
rect 160881 -16408 160882 -16363
rect 160981 -16374 160982 -16363
rect 161557 -16367 161592 -16333
rect 161734 -16367 161769 -16333
rect 162327 -16336 162328 -16328
rect 162427 -16336 162428 -16328
rect 160992 -16408 161027 -16374
rect 159094 -16453 159129 -16419
rect 160373 -16422 160374 -16414
rect 161723 -16417 161724 -16406
rect 161928 -16410 161963 -16376
rect 161973 -16410 161974 -16365
rect 162073 -16376 162074 -16365
rect 162254 -16370 162317 -16336
rect 162326 -16370 162361 -16336
rect 162438 -16370 162473 -16336
rect 163163 -16360 163198 -16326
rect 163259 -16360 163294 -16326
rect 163355 -16360 163390 -16326
rect 163451 -16360 163486 -16326
rect 163547 -16360 163582 -16326
rect 163643 -16360 163678 -16326
rect 163739 -16360 163774 -16326
rect 165067 -16333 165068 -16322
rect 165244 -16327 165307 -16293
rect 165316 -16327 165351 -16293
rect 165428 -16327 165463 -16293
rect 165959 -16317 165994 -16283
rect 166055 -16317 166090 -16283
rect 166151 -16317 166186 -16283
rect 166247 -16317 166282 -16283
rect 166343 -16317 166378 -16283
rect 167368 -16324 167403 -16290
rect 167413 -16324 167414 -16279
rect 167513 -16290 167514 -16279
rect 167524 -16324 167559 -16290
rect 167569 -16324 167570 -16279
rect 167669 -16290 167670 -16279
rect 167848 -16284 167883 -16250
rect 167920 -16284 167955 -16250
rect 167992 -16284 168027 -16250
rect 168136 -16284 168171 -16250
rect 168208 -16284 168243 -16250
rect 168245 -16284 168315 -16250
rect 168352 -16284 168387 -16250
rect 168422 -16284 168457 -16250
rect 168949 -16274 168984 -16240
rect 169045 -16274 169080 -16240
rect 169141 -16274 169176 -16240
rect 170648 -16241 170683 -16207
rect 170712 -16241 170755 -16207
rect 170757 -16241 170758 -16199
rect 170857 -16207 170858 -16199
rect 170792 -16241 170827 -16207
rect 170868 -16241 170903 -16207
rect 170913 -16241 170914 -16199
rect 171013 -16207 171014 -16199
rect 170962 -16241 170997 -16207
rect 171024 -16241 171069 -16207
rect 171939 -16231 171974 -16197
rect 172035 -16231 172070 -16197
rect 172131 -16231 172166 -16197
rect 171755 -16250 171756 -16242
rect 167680 -16324 167715 -16290
rect 168661 -16293 168662 -16285
rect 168761 -16293 168762 -16285
rect 162084 -16410 162119 -16376
rect 158740 -16494 158775 -16460
rect 155750 -16620 155785 -16586
rect 157029 -16589 157030 -16578
rect 154279 -16689 154280 -16681
rect 154290 -16723 154325 -16689
rect 154510 -16734 154545 -16700
rect 152957 -16793 152992 -16759
rect 153160 -16838 153195 -16804
rect 153283 -16809 153284 -16767
rect 153605 -16796 153640 -16762
rect 152927 -16861 152928 -16853
rect 152938 -16895 152973 -16861
rect 153160 -16906 153195 -16872
rect 152927 -16961 152928 -16950
rect 152938 -16995 152973 -16961
rect 151875 -17045 151910 -17011
rect 151971 -17045 152006 -17011
rect 152067 -17045 152102 -17011
rect 152576 -17035 152611 -17001
rect 152648 -17035 152683 -17001
rect 152720 -17035 152755 -17001
rect 152792 -17029 152828 -17001
rect 153138 -17025 153173 -16991
rect 153183 -17025 153184 -16980
rect 152792 -17035 152827 -17029
rect 152229 -17088 152264 -17054
rect 152325 -17088 152360 -17054
rect 152421 -17088 152456 -17054
rect 153325 -17076 153326 -16809
rect 153954 -16819 154341 -16753
rect 153341 -16860 153376 -16826
rect 153690 -16832 153701 -16819
rect 153624 -16874 153701 -16832
rect 153752 -16874 154341 -16819
rect 154488 -16853 154523 -16819
rect 154533 -16853 154534 -16808
rect 153624 -16877 154341 -16874
rect 153341 -16928 153376 -16894
rect 153544 -16942 153579 -16908
rect 153589 -16942 153590 -16900
rect 153425 -16991 153426 -16980
rect 153436 -17025 153471 -16991
rect 153544 -17042 153579 -17008
rect 153589 -17042 153590 -16997
rect 153437 -17078 153472 -17044
rect 153509 -17078 153544 -17044
rect 153581 -17078 153616 -17044
rect 152583 -17131 152618 -17097
rect 152679 -17131 152714 -17097
rect 152775 -17131 152810 -17097
rect 152871 -17131 152906 -17097
rect 152967 -17131 153002 -17097
rect 153624 -17114 153769 -16877
rect 153954 -16899 154341 -16877
rect 153878 -16925 154341 -16899
rect 154675 -16904 154676 -16637
rect 154691 -16688 154726 -16654
rect 155305 -16691 155340 -16657
rect 155984 -16663 156019 -16629
rect 156029 -16663 156030 -16618
rect 156129 -16629 156130 -16618
rect 156140 -16663 156175 -16629
rect 156185 -16663 156186 -16618
rect 156285 -16629 156286 -16618
rect 156863 -16623 156898 -16589
rect 157040 -16623 157075 -16589
rect 157401 -16605 157436 -16571
rect 156296 -16663 156331 -16629
rect 156129 -16697 156130 -16671
rect 156528 -16689 156563 -16655
rect 156573 -16689 156574 -16644
rect 156673 -16655 156674 -16644
rect 156684 -16689 156719 -16655
rect 156729 -16689 156730 -16644
rect 157029 -16672 157030 -16661
rect 154691 -16756 154726 -16722
rect 154894 -16770 154929 -16736
rect 154939 -16770 154940 -16728
rect 155039 -16740 155040 -16729
rect 155659 -16734 155694 -16700
rect 155050 -16774 155085 -16740
rect 154775 -16819 154776 -16808
rect 155244 -16813 155279 -16779
rect 155289 -16813 155290 -16771
rect 155389 -16779 155390 -16771
rect 156049 -16777 156084 -16743
rect 155400 -16813 155435 -16779
rect 154786 -16853 154821 -16819
rect 154894 -16870 154929 -16836
rect 154939 -16870 154940 -16825
rect 155039 -16832 155040 -16821
rect 155050 -16866 155085 -16832
rect 155598 -16856 155633 -16822
rect 155643 -16856 155644 -16814
rect 155743 -16822 155744 -16814
rect 155754 -16856 155789 -16822
rect 154787 -16906 154822 -16872
rect 154859 -16906 154894 -16872
rect 154931 -16906 154966 -16872
rect 155244 -16913 155279 -16879
rect 155289 -16913 155290 -16868
rect 155389 -16879 155390 -16868
rect 155400 -16913 155435 -16879
rect 155984 -16895 156019 -16861
rect 156029 -16895 156030 -16853
rect 153878 -16959 154354 -16925
rect 155212 -16949 155247 -16915
rect 155284 -16949 155319 -16915
rect 155598 -16956 155633 -16922
rect 155643 -16956 155644 -16911
rect 155743 -16922 155744 -16911
rect 155754 -16956 155789 -16922
rect 153878 -16985 154341 -16959
rect 153882 -16993 154083 -16985
rect 153898 -17003 154067 -16993
rect 153624 -17140 153799 -17114
rect 153131 -17174 153166 -17140
rect 153227 -17174 153262 -17140
rect 153323 -17174 153358 -17140
rect 153419 -17174 153454 -17140
rect 153515 -17174 153550 -17140
rect 153611 -17174 153799 -17140
rect 153624 -17200 153799 -17174
rect 153824 -17174 153925 -17050
rect 153702 -17870 153737 -17200
rect 153824 -17228 153827 -17174
rect 153509 -17936 153654 -17924
rect 153177 -17970 153654 -17936
rect 153509 -17971 153654 -17970
rect 153690 -17971 153737 -17870
rect 153836 -17971 153871 -17174
rect 154094 -17971 154129 -17062
rect 154228 -17971 154263 -16985
rect 154481 -17002 154516 -16968
rect 154577 -17002 154612 -16968
rect 154673 -17002 154708 -16968
rect 154769 -17002 154804 -16968
rect 154865 -17002 154900 -16968
rect 154961 -17002 154996 -16968
rect 155057 -17002 155092 -16968
rect 155566 -16992 155601 -16958
rect 155638 -16992 155673 -16958
rect 155984 -16995 156019 -16961
rect 156029 -16995 156030 -16950
rect 156171 -17001 156172 -16697
rect 156863 -16706 156898 -16672
rect 157040 -16706 157075 -16672
rect 157336 -16723 157371 -16689
rect 157381 -16723 157382 -16681
rect 157523 -16753 157524 -16525
rect 158213 -16534 158248 -16500
rect 158390 -16534 158425 -16500
rect 158584 -16577 158619 -16543
rect 158629 -16577 158630 -16532
rect 158729 -16543 158730 -16532
rect 158938 -16537 158973 -16503
rect 158983 -16537 158984 -16492
rect 159083 -16503 159084 -16492
rect 159328 -16496 159363 -16462
rect 159373 -16496 159374 -16451
rect 159473 -16462 159474 -16451
rect 159484 -16496 159519 -16462
rect 159529 -16496 159530 -16451
rect 159629 -16462 159630 -16451
rect 159810 -16456 159845 -16422
rect 159882 -16456 159917 -16422
rect 159954 -16456 159989 -16422
rect 160098 -16456 160133 -16422
rect 160170 -16456 160205 -16422
rect 160207 -16456 160277 -16422
rect 160314 -16456 160349 -16422
rect 160384 -16456 160419 -16422
rect 159640 -16496 159675 -16462
rect 160680 -16491 160715 -16457
rect 160725 -16491 160726 -16446
rect 160825 -16457 160826 -16446
rect 160836 -16491 160871 -16457
rect 160881 -16491 160882 -16446
rect 160981 -16457 160982 -16446
rect 161557 -16451 161592 -16417
rect 161734 -16451 161769 -16417
rect 160992 -16491 161027 -16457
rect 159094 -16537 159129 -16503
rect 160373 -16505 160374 -16494
rect 158740 -16577 158775 -16543
rect 157653 -16621 157688 -16587
rect 157854 -16666 157889 -16632
rect 157977 -16637 157978 -16595
rect 158299 -16624 158334 -16590
rect 158938 -16620 158973 -16586
rect 158983 -16620 158984 -16575
rect 159083 -16586 159084 -16575
rect 159328 -16580 159363 -16546
rect 159373 -16580 159374 -16535
rect 159473 -16546 159474 -16535
rect 159484 -16580 159519 -16546
rect 159529 -16580 159530 -16535
rect 159629 -16546 159630 -16535
rect 160207 -16539 160242 -16505
rect 160384 -16539 160419 -16505
rect 159640 -16580 159675 -16546
rect 160527 -16565 160642 -16499
rect 160825 -16525 160826 -16499
rect 161222 -16517 161257 -16483
rect 161267 -16517 161268 -16472
rect 161367 -16483 161368 -16472
rect 161378 -16517 161413 -16483
rect 161423 -16517 161424 -16472
rect 161723 -16500 161724 -16489
rect 161928 -16494 161963 -16460
rect 161973 -16494 161974 -16449
rect 162073 -16460 162074 -16449
rect 162282 -16453 162317 -16419
rect 162327 -16453 162328 -16408
rect 162427 -16419 162428 -16408
rect 162608 -16413 162643 -16379
rect 162672 -16413 162715 -16379
rect 162717 -16413 162718 -16371
rect 162817 -16379 162818 -16371
rect 162752 -16413 162787 -16379
rect 162828 -16413 162863 -16379
rect 162873 -16413 162874 -16371
rect 162973 -16379 162974 -16371
rect 162922 -16413 162957 -16379
rect 162984 -16413 163029 -16379
rect 164024 -16408 164059 -16374
rect 164069 -16408 164070 -16363
rect 164169 -16374 164170 -16363
rect 164180 -16408 164215 -16374
rect 164225 -16408 164226 -16363
rect 164325 -16374 164326 -16363
rect 164901 -16367 164936 -16333
rect 165078 -16367 165113 -16333
rect 165671 -16336 165672 -16328
rect 165771 -16336 165772 -16328
rect 164336 -16408 164371 -16374
rect 162438 -16453 162473 -16419
rect 163717 -16422 163718 -16414
rect 165067 -16417 165068 -16406
rect 165272 -16410 165307 -16376
rect 165317 -16410 165318 -16365
rect 165417 -16376 165418 -16365
rect 165598 -16370 165661 -16336
rect 165670 -16370 165705 -16336
rect 165782 -16370 165817 -16336
rect 166507 -16360 166542 -16326
rect 166603 -16360 166638 -16326
rect 166699 -16360 166734 -16326
rect 166795 -16360 166830 -16326
rect 166891 -16360 166926 -16326
rect 166987 -16360 167022 -16326
rect 167083 -16360 167118 -16326
rect 168411 -16333 168412 -16322
rect 168588 -16327 168651 -16293
rect 168660 -16327 168695 -16293
rect 168772 -16327 168807 -16293
rect 169303 -16317 169338 -16283
rect 169399 -16317 169434 -16283
rect 169495 -16317 169530 -16283
rect 169591 -16317 169626 -16283
rect 169687 -16317 169722 -16283
rect 170712 -16324 170747 -16290
rect 170757 -16324 170758 -16279
rect 170857 -16290 170858 -16279
rect 170868 -16324 170903 -16290
rect 170913 -16324 170914 -16279
rect 171013 -16290 171014 -16279
rect 171192 -16284 171227 -16250
rect 171264 -16284 171299 -16250
rect 171336 -16284 171371 -16250
rect 171480 -16284 171515 -16250
rect 171552 -16284 171587 -16250
rect 171589 -16284 171659 -16250
rect 171696 -16284 171731 -16250
rect 171766 -16284 171801 -16250
rect 172293 -16274 172328 -16240
rect 172389 -16274 172424 -16240
rect 172485 -16274 172520 -16240
rect 173992 -16241 174027 -16207
rect 174056 -16241 174099 -16207
rect 174101 -16241 174102 -16199
rect 174201 -16207 174202 -16199
rect 174136 -16241 174171 -16207
rect 174212 -16241 174247 -16207
rect 174257 -16241 174258 -16199
rect 174357 -16207 174358 -16199
rect 174306 -16241 174341 -16207
rect 174368 -16241 174413 -16207
rect 175283 -16231 175318 -16197
rect 175379 -16231 175414 -16197
rect 175475 -16231 175510 -16197
rect 175099 -16250 175100 -16242
rect 171024 -16324 171059 -16290
rect 172005 -16293 172006 -16285
rect 172105 -16293 172106 -16285
rect 165428 -16410 165463 -16376
rect 162084 -16494 162119 -16460
rect 159094 -16620 159129 -16586
rect 160373 -16589 160374 -16578
rect 157623 -16689 157624 -16681
rect 157634 -16723 157669 -16689
rect 157854 -16734 157889 -16700
rect 156301 -16793 156336 -16759
rect 156504 -16838 156539 -16804
rect 156627 -16809 156628 -16767
rect 156949 -16796 156984 -16762
rect 156271 -16861 156272 -16853
rect 156282 -16895 156317 -16861
rect 156504 -16906 156539 -16872
rect 156271 -16961 156272 -16950
rect 156282 -16995 156317 -16961
rect 155219 -17045 155254 -17011
rect 155315 -17045 155350 -17011
rect 155411 -17045 155446 -17011
rect 155920 -17035 155955 -17001
rect 155992 -17035 156027 -17001
rect 156064 -17035 156099 -17001
rect 156136 -17029 156172 -17001
rect 156482 -17025 156517 -16991
rect 156527 -17025 156528 -16980
rect 156136 -17035 156171 -17029
rect 155573 -17088 155608 -17054
rect 155669 -17088 155704 -17054
rect 155765 -17088 155800 -17054
rect 156669 -17076 156670 -16809
rect 157298 -16819 157685 -16753
rect 156685 -16860 156720 -16826
rect 157034 -16832 157045 -16819
rect 156968 -16874 157045 -16832
rect 157096 -16874 157685 -16819
rect 157832 -16853 157867 -16819
rect 157877 -16853 157878 -16808
rect 156968 -16877 157685 -16874
rect 156685 -16928 156720 -16894
rect 156888 -16942 156923 -16908
rect 156933 -16942 156934 -16900
rect 156769 -16991 156770 -16980
rect 156780 -17025 156815 -16991
rect 156888 -17042 156923 -17008
rect 156933 -17042 156934 -16997
rect 156781 -17078 156816 -17044
rect 156853 -17078 156888 -17044
rect 156925 -17078 156960 -17044
rect 155927 -17131 155962 -17097
rect 156023 -17131 156058 -17097
rect 156119 -17131 156154 -17097
rect 156215 -17131 156250 -17097
rect 156311 -17131 156346 -17097
rect 156968 -17114 157113 -16877
rect 157298 -16899 157685 -16877
rect 157222 -16925 157685 -16899
rect 158019 -16904 158020 -16637
rect 158035 -16688 158070 -16654
rect 158649 -16691 158684 -16657
rect 159328 -16663 159363 -16629
rect 159373 -16663 159374 -16618
rect 159473 -16629 159474 -16618
rect 159484 -16663 159519 -16629
rect 159529 -16663 159530 -16618
rect 159629 -16629 159630 -16618
rect 160207 -16623 160242 -16589
rect 160384 -16623 160419 -16589
rect 160745 -16605 160780 -16571
rect 159640 -16663 159675 -16629
rect 159473 -16697 159474 -16671
rect 159872 -16689 159907 -16655
rect 159917 -16689 159918 -16644
rect 160017 -16655 160018 -16644
rect 160028 -16689 160063 -16655
rect 160073 -16689 160074 -16644
rect 160373 -16672 160374 -16661
rect 158035 -16756 158070 -16722
rect 158238 -16770 158273 -16736
rect 158283 -16770 158284 -16728
rect 158383 -16740 158384 -16729
rect 159003 -16734 159038 -16700
rect 158394 -16774 158429 -16740
rect 158119 -16819 158120 -16808
rect 158588 -16813 158623 -16779
rect 158633 -16813 158634 -16771
rect 158733 -16779 158734 -16771
rect 159393 -16777 159428 -16743
rect 158744 -16813 158779 -16779
rect 158130 -16853 158165 -16819
rect 158238 -16870 158273 -16836
rect 158283 -16870 158284 -16825
rect 158383 -16832 158384 -16821
rect 158394 -16866 158429 -16832
rect 158942 -16856 158977 -16822
rect 158987 -16856 158988 -16814
rect 159087 -16822 159088 -16814
rect 159098 -16856 159133 -16822
rect 158131 -16906 158166 -16872
rect 158203 -16906 158238 -16872
rect 158275 -16906 158310 -16872
rect 158588 -16913 158623 -16879
rect 158633 -16913 158634 -16868
rect 158733 -16879 158734 -16868
rect 158744 -16913 158779 -16879
rect 159328 -16895 159363 -16861
rect 159373 -16895 159374 -16853
rect 157222 -16959 157698 -16925
rect 158556 -16949 158591 -16915
rect 158628 -16949 158663 -16915
rect 158942 -16956 158977 -16922
rect 158987 -16956 158988 -16911
rect 159087 -16922 159088 -16911
rect 159098 -16956 159133 -16922
rect 157222 -16985 157685 -16959
rect 157226 -16993 157427 -16985
rect 157242 -17003 157411 -16993
rect 156968 -17140 157143 -17114
rect 156475 -17174 156510 -17140
rect 156571 -17174 156606 -17140
rect 156667 -17174 156702 -17140
rect 156763 -17174 156798 -17140
rect 156859 -17174 156894 -17140
rect 156955 -17174 157143 -17140
rect 156968 -17200 157143 -17174
rect 157168 -17174 157269 -17050
rect 157046 -17870 157081 -17200
rect 157168 -17228 157171 -17174
rect 156853 -17936 156998 -17924
rect 156521 -17970 156998 -17936
rect 156853 -17971 156998 -17970
rect 157034 -17971 157081 -17870
rect 157180 -17971 157215 -17174
rect 157438 -17971 157473 -17062
rect 157572 -17971 157607 -16985
rect 157825 -17002 157860 -16968
rect 157921 -17002 157956 -16968
rect 158017 -17002 158052 -16968
rect 158113 -17002 158148 -16968
rect 158209 -17002 158244 -16968
rect 158305 -17002 158340 -16968
rect 158401 -17002 158436 -16968
rect 158910 -16992 158945 -16958
rect 158982 -16992 159017 -16958
rect 159328 -16995 159363 -16961
rect 159373 -16995 159374 -16950
rect 159515 -17001 159516 -16697
rect 160207 -16706 160242 -16672
rect 160384 -16706 160419 -16672
rect 160680 -16723 160715 -16689
rect 160725 -16723 160726 -16681
rect 160867 -16753 160868 -16525
rect 161557 -16534 161592 -16500
rect 161734 -16534 161769 -16500
rect 161928 -16577 161963 -16543
rect 161973 -16577 161974 -16532
rect 162073 -16543 162074 -16532
rect 162282 -16537 162317 -16503
rect 162327 -16537 162328 -16492
rect 162427 -16503 162428 -16492
rect 162672 -16496 162707 -16462
rect 162717 -16496 162718 -16451
rect 162817 -16462 162818 -16451
rect 162828 -16496 162863 -16462
rect 162873 -16496 162874 -16451
rect 162973 -16462 162974 -16451
rect 163154 -16456 163189 -16422
rect 163226 -16456 163261 -16422
rect 163298 -16456 163333 -16422
rect 163442 -16456 163477 -16422
rect 163514 -16456 163549 -16422
rect 163551 -16456 163621 -16422
rect 163658 -16456 163693 -16422
rect 163728 -16456 163763 -16422
rect 162984 -16496 163019 -16462
rect 164024 -16491 164059 -16457
rect 164069 -16491 164070 -16446
rect 164169 -16457 164170 -16446
rect 164180 -16491 164215 -16457
rect 164225 -16491 164226 -16446
rect 164325 -16457 164326 -16446
rect 164901 -16451 164936 -16417
rect 165078 -16451 165113 -16417
rect 164336 -16491 164371 -16457
rect 162438 -16537 162473 -16503
rect 163717 -16505 163718 -16494
rect 162084 -16577 162119 -16543
rect 160997 -16621 161032 -16587
rect 161198 -16666 161233 -16632
rect 161321 -16637 161322 -16595
rect 161643 -16624 161678 -16590
rect 162282 -16620 162317 -16586
rect 162327 -16620 162328 -16575
rect 162427 -16586 162428 -16575
rect 162672 -16580 162707 -16546
rect 162717 -16580 162718 -16535
rect 162817 -16546 162818 -16535
rect 162828 -16580 162863 -16546
rect 162873 -16580 162874 -16535
rect 162973 -16546 162974 -16535
rect 163551 -16539 163586 -16505
rect 163728 -16539 163763 -16505
rect 162984 -16580 163019 -16546
rect 163871 -16565 163986 -16499
rect 164169 -16525 164170 -16499
rect 164566 -16517 164601 -16483
rect 164611 -16517 164612 -16472
rect 164711 -16483 164712 -16472
rect 164722 -16517 164757 -16483
rect 164767 -16517 164768 -16472
rect 165067 -16500 165068 -16489
rect 165272 -16494 165307 -16460
rect 165317 -16494 165318 -16449
rect 165417 -16460 165418 -16449
rect 165626 -16453 165661 -16419
rect 165671 -16453 165672 -16408
rect 165771 -16419 165772 -16408
rect 165952 -16413 165987 -16379
rect 166016 -16413 166059 -16379
rect 166061 -16413 166062 -16371
rect 166161 -16379 166162 -16371
rect 166096 -16413 166131 -16379
rect 166172 -16413 166207 -16379
rect 166217 -16413 166218 -16371
rect 166317 -16379 166318 -16371
rect 166266 -16413 166301 -16379
rect 166328 -16413 166373 -16379
rect 167368 -16408 167403 -16374
rect 167413 -16408 167414 -16363
rect 167513 -16374 167514 -16363
rect 167524 -16408 167559 -16374
rect 167569 -16408 167570 -16363
rect 167669 -16374 167670 -16363
rect 168245 -16367 168280 -16333
rect 168422 -16367 168457 -16333
rect 169015 -16336 169016 -16328
rect 169115 -16336 169116 -16328
rect 167680 -16408 167715 -16374
rect 165782 -16453 165817 -16419
rect 167061 -16422 167062 -16414
rect 168411 -16417 168412 -16406
rect 168616 -16410 168651 -16376
rect 168661 -16410 168662 -16365
rect 168761 -16376 168762 -16365
rect 168942 -16370 169005 -16336
rect 169014 -16370 169049 -16336
rect 169126 -16370 169161 -16336
rect 169851 -16360 169886 -16326
rect 169947 -16360 169982 -16326
rect 170043 -16360 170078 -16326
rect 170139 -16360 170174 -16326
rect 170235 -16360 170270 -16326
rect 170331 -16360 170366 -16326
rect 170427 -16360 170462 -16326
rect 171755 -16333 171756 -16322
rect 171932 -16327 171995 -16293
rect 172004 -16327 172039 -16293
rect 172116 -16327 172151 -16293
rect 172647 -16317 172682 -16283
rect 172743 -16317 172778 -16283
rect 172839 -16317 172874 -16283
rect 172935 -16317 172970 -16283
rect 173031 -16317 173066 -16283
rect 174056 -16324 174091 -16290
rect 174101 -16324 174102 -16279
rect 174201 -16290 174202 -16279
rect 174212 -16324 174247 -16290
rect 174257 -16324 174258 -16279
rect 174357 -16290 174358 -16279
rect 174536 -16284 174571 -16250
rect 174608 -16284 174643 -16250
rect 174680 -16284 174715 -16250
rect 174824 -16284 174859 -16250
rect 174896 -16284 174931 -16250
rect 174933 -16284 175003 -16250
rect 175040 -16284 175075 -16250
rect 175110 -16284 175145 -16250
rect 175637 -16274 175672 -16240
rect 175733 -16274 175768 -16240
rect 175829 -16274 175864 -16240
rect 177336 -16241 177371 -16207
rect 177400 -16241 177443 -16207
rect 177445 -16241 177446 -16199
rect 177545 -16207 177546 -16199
rect 177480 -16241 177515 -16207
rect 177556 -16241 177591 -16207
rect 177601 -16241 177602 -16199
rect 177701 -16207 177702 -16199
rect 177650 -16241 177685 -16207
rect 177712 -16241 177757 -16207
rect 178627 -16231 178662 -16197
rect 178723 -16231 178758 -16197
rect 178819 -16231 178854 -16197
rect 178443 -16250 178444 -16242
rect 174368 -16324 174403 -16290
rect 175349 -16293 175350 -16285
rect 175449 -16293 175450 -16285
rect 168772 -16410 168807 -16376
rect 165428 -16494 165463 -16460
rect 162438 -16620 162473 -16586
rect 163717 -16589 163718 -16578
rect 160967 -16689 160968 -16681
rect 160978 -16723 161013 -16689
rect 161198 -16734 161233 -16700
rect 159645 -16793 159680 -16759
rect 159848 -16838 159883 -16804
rect 159971 -16809 159972 -16767
rect 160293 -16796 160328 -16762
rect 159615 -16861 159616 -16853
rect 159626 -16895 159661 -16861
rect 159848 -16906 159883 -16872
rect 159615 -16961 159616 -16950
rect 159626 -16995 159661 -16961
rect 158563 -17045 158598 -17011
rect 158659 -17045 158694 -17011
rect 158755 -17045 158790 -17011
rect 159264 -17035 159299 -17001
rect 159336 -17035 159371 -17001
rect 159408 -17035 159443 -17001
rect 159480 -17029 159516 -17001
rect 159826 -17025 159861 -16991
rect 159871 -17025 159872 -16980
rect 159480 -17035 159515 -17029
rect 158917 -17088 158952 -17054
rect 159013 -17088 159048 -17054
rect 159109 -17088 159144 -17054
rect 160013 -17076 160014 -16809
rect 160642 -16819 161029 -16753
rect 160029 -16860 160064 -16826
rect 160378 -16832 160389 -16819
rect 160312 -16874 160389 -16832
rect 160440 -16874 161029 -16819
rect 161176 -16853 161211 -16819
rect 161221 -16853 161222 -16808
rect 160312 -16877 161029 -16874
rect 160029 -16928 160064 -16894
rect 160232 -16942 160267 -16908
rect 160277 -16942 160278 -16900
rect 160113 -16991 160114 -16980
rect 160124 -17025 160159 -16991
rect 160232 -17042 160267 -17008
rect 160277 -17042 160278 -16997
rect 160125 -17078 160160 -17044
rect 160197 -17078 160232 -17044
rect 160269 -17078 160304 -17044
rect 159271 -17131 159306 -17097
rect 159367 -17131 159402 -17097
rect 159463 -17131 159498 -17097
rect 159559 -17131 159594 -17097
rect 159655 -17131 159690 -17097
rect 160312 -17114 160457 -16877
rect 160642 -16899 161029 -16877
rect 160566 -16925 161029 -16899
rect 161363 -16904 161364 -16637
rect 161379 -16688 161414 -16654
rect 161993 -16691 162028 -16657
rect 162672 -16663 162707 -16629
rect 162717 -16663 162718 -16618
rect 162817 -16629 162818 -16618
rect 162828 -16663 162863 -16629
rect 162873 -16663 162874 -16618
rect 162973 -16629 162974 -16618
rect 163551 -16623 163586 -16589
rect 163728 -16623 163763 -16589
rect 164089 -16605 164124 -16571
rect 162984 -16663 163019 -16629
rect 162817 -16697 162818 -16671
rect 163216 -16689 163251 -16655
rect 163261 -16689 163262 -16644
rect 163361 -16655 163362 -16644
rect 163372 -16689 163407 -16655
rect 163417 -16689 163418 -16644
rect 163717 -16672 163718 -16661
rect 161379 -16756 161414 -16722
rect 161582 -16770 161617 -16736
rect 161627 -16770 161628 -16728
rect 161727 -16740 161728 -16729
rect 162347 -16734 162382 -16700
rect 161738 -16774 161773 -16740
rect 161463 -16819 161464 -16808
rect 161932 -16813 161967 -16779
rect 161977 -16813 161978 -16771
rect 162077 -16779 162078 -16771
rect 162737 -16777 162772 -16743
rect 162088 -16813 162123 -16779
rect 161474 -16853 161509 -16819
rect 161582 -16870 161617 -16836
rect 161627 -16870 161628 -16825
rect 161727 -16832 161728 -16821
rect 161738 -16866 161773 -16832
rect 162286 -16856 162321 -16822
rect 162331 -16856 162332 -16814
rect 162431 -16822 162432 -16814
rect 162442 -16856 162477 -16822
rect 161475 -16906 161510 -16872
rect 161547 -16906 161582 -16872
rect 161619 -16906 161654 -16872
rect 161932 -16913 161967 -16879
rect 161977 -16913 161978 -16868
rect 162077 -16879 162078 -16868
rect 162088 -16913 162123 -16879
rect 162672 -16895 162707 -16861
rect 162717 -16895 162718 -16853
rect 160566 -16959 161042 -16925
rect 161900 -16949 161935 -16915
rect 161972 -16949 162007 -16915
rect 162286 -16956 162321 -16922
rect 162331 -16956 162332 -16911
rect 162431 -16922 162432 -16911
rect 162442 -16956 162477 -16922
rect 160566 -16985 161029 -16959
rect 160570 -16993 160771 -16985
rect 160586 -17003 160755 -16993
rect 160312 -17140 160487 -17114
rect 159819 -17174 159854 -17140
rect 159915 -17174 159950 -17140
rect 160011 -17174 160046 -17140
rect 160107 -17174 160142 -17140
rect 160203 -17174 160238 -17140
rect 160299 -17174 160487 -17140
rect 160312 -17200 160487 -17174
rect 160512 -17174 160613 -17050
rect 160390 -17870 160425 -17200
rect 160512 -17228 160515 -17174
rect 160197 -17936 160342 -17924
rect 159865 -17970 160342 -17936
rect 160197 -17971 160342 -17970
rect 160378 -17971 160425 -17870
rect 160524 -17971 160559 -17174
rect 160782 -17971 160817 -17062
rect 160916 -17971 160951 -16985
rect 161169 -17002 161204 -16968
rect 161265 -17002 161300 -16968
rect 161361 -17002 161396 -16968
rect 161457 -17002 161492 -16968
rect 161553 -17002 161588 -16968
rect 161649 -17002 161684 -16968
rect 161745 -17002 161780 -16968
rect 162254 -16992 162289 -16958
rect 162326 -16992 162361 -16958
rect 162672 -16995 162707 -16961
rect 162717 -16995 162718 -16950
rect 162859 -17001 162860 -16697
rect 163551 -16706 163586 -16672
rect 163728 -16706 163763 -16672
rect 164024 -16723 164059 -16689
rect 164069 -16723 164070 -16681
rect 164211 -16753 164212 -16525
rect 164901 -16534 164936 -16500
rect 165078 -16534 165113 -16500
rect 165272 -16577 165307 -16543
rect 165317 -16577 165318 -16532
rect 165417 -16543 165418 -16532
rect 165626 -16537 165661 -16503
rect 165671 -16537 165672 -16492
rect 165771 -16503 165772 -16492
rect 166016 -16496 166051 -16462
rect 166061 -16496 166062 -16451
rect 166161 -16462 166162 -16451
rect 166172 -16496 166207 -16462
rect 166217 -16496 166218 -16451
rect 166317 -16462 166318 -16451
rect 166498 -16456 166533 -16422
rect 166570 -16456 166605 -16422
rect 166642 -16456 166677 -16422
rect 166786 -16456 166821 -16422
rect 166858 -16456 166893 -16422
rect 166895 -16456 166965 -16422
rect 167002 -16456 167037 -16422
rect 167072 -16456 167107 -16422
rect 166328 -16496 166363 -16462
rect 167368 -16491 167403 -16457
rect 167413 -16491 167414 -16446
rect 167513 -16457 167514 -16446
rect 167524 -16491 167559 -16457
rect 167569 -16491 167570 -16446
rect 167669 -16457 167670 -16446
rect 168245 -16451 168280 -16417
rect 168422 -16451 168457 -16417
rect 167680 -16491 167715 -16457
rect 165782 -16537 165817 -16503
rect 167061 -16505 167062 -16494
rect 165428 -16577 165463 -16543
rect 164341 -16621 164376 -16587
rect 164542 -16666 164577 -16632
rect 164665 -16637 164666 -16595
rect 164987 -16624 165022 -16590
rect 165626 -16620 165661 -16586
rect 165671 -16620 165672 -16575
rect 165771 -16586 165772 -16575
rect 166016 -16580 166051 -16546
rect 166061 -16580 166062 -16535
rect 166161 -16546 166162 -16535
rect 166172 -16580 166207 -16546
rect 166217 -16580 166218 -16535
rect 166317 -16546 166318 -16535
rect 166895 -16539 166930 -16505
rect 167072 -16539 167107 -16505
rect 166328 -16580 166363 -16546
rect 167215 -16565 167330 -16499
rect 167513 -16525 167514 -16499
rect 167910 -16517 167945 -16483
rect 167955 -16517 167956 -16472
rect 168055 -16483 168056 -16472
rect 168066 -16517 168101 -16483
rect 168111 -16517 168112 -16472
rect 168411 -16500 168412 -16489
rect 168616 -16494 168651 -16460
rect 168661 -16494 168662 -16449
rect 168761 -16460 168762 -16449
rect 168970 -16453 169005 -16419
rect 169015 -16453 169016 -16408
rect 169115 -16419 169116 -16408
rect 169296 -16413 169331 -16379
rect 169360 -16413 169403 -16379
rect 169405 -16413 169406 -16371
rect 169505 -16379 169506 -16371
rect 169440 -16413 169475 -16379
rect 169516 -16413 169551 -16379
rect 169561 -16413 169562 -16371
rect 169661 -16379 169662 -16371
rect 169610 -16413 169645 -16379
rect 169672 -16413 169717 -16379
rect 170712 -16408 170747 -16374
rect 170757 -16408 170758 -16363
rect 170857 -16374 170858 -16363
rect 170868 -16408 170903 -16374
rect 170913 -16408 170914 -16363
rect 171013 -16374 171014 -16363
rect 171589 -16367 171624 -16333
rect 171766 -16367 171801 -16333
rect 172359 -16336 172360 -16328
rect 172459 -16336 172460 -16328
rect 171024 -16408 171059 -16374
rect 169126 -16453 169161 -16419
rect 170405 -16422 170406 -16414
rect 171755 -16417 171756 -16406
rect 171960 -16410 171995 -16376
rect 172005 -16410 172006 -16365
rect 172105 -16376 172106 -16365
rect 172286 -16370 172349 -16336
rect 172358 -16370 172393 -16336
rect 172470 -16370 172505 -16336
rect 173195 -16360 173230 -16326
rect 173291 -16360 173326 -16326
rect 173387 -16360 173422 -16326
rect 173483 -16360 173518 -16326
rect 173579 -16360 173614 -16326
rect 173675 -16360 173710 -16326
rect 173771 -16360 173806 -16326
rect 175099 -16333 175100 -16322
rect 175276 -16327 175339 -16293
rect 175348 -16327 175383 -16293
rect 175460 -16327 175495 -16293
rect 175991 -16317 176026 -16283
rect 176087 -16317 176122 -16283
rect 176183 -16317 176218 -16283
rect 176279 -16317 176314 -16283
rect 176375 -16317 176410 -16283
rect 177400 -16324 177435 -16290
rect 177445 -16324 177446 -16279
rect 177545 -16290 177546 -16279
rect 177556 -16324 177591 -16290
rect 177601 -16324 177602 -16279
rect 177701 -16290 177702 -16279
rect 177880 -16284 177915 -16250
rect 177952 -16284 177987 -16250
rect 178024 -16284 178059 -16250
rect 178168 -16284 178203 -16250
rect 178240 -16284 178275 -16250
rect 178277 -16284 178347 -16250
rect 178384 -16284 178419 -16250
rect 178454 -16284 178489 -16250
rect 178981 -16274 179016 -16240
rect 179077 -16274 179112 -16240
rect 179173 -16274 179208 -16240
rect 180680 -16241 180715 -16207
rect 180744 -16241 180787 -16207
rect 180789 -16241 180790 -16199
rect 180889 -16207 180890 -16199
rect 180824 -16241 180859 -16207
rect 180900 -16241 180935 -16207
rect 180945 -16241 180946 -16199
rect 181045 -16207 181046 -16199
rect 180994 -16241 181029 -16207
rect 181056 -16241 181101 -16207
rect 181971 -16231 182006 -16197
rect 182067 -16231 182102 -16197
rect 182163 -16231 182198 -16197
rect 181787 -16250 181788 -16242
rect 177712 -16324 177747 -16290
rect 178693 -16293 178694 -16285
rect 178793 -16293 178794 -16285
rect 172116 -16410 172151 -16376
rect 168772 -16494 168807 -16460
rect 165782 -16620 165817 -16586
rect 167061 -16589 167062 -16578
rect 164311 -16689 164312 -16681
rect 164322 -16723 164357 -16689
rect 164542 -16734 164577 -16700
rect 162989 -16793 163024 -16759
rect 163192 -16838 163227 -16804
rect 163315 -16809 163316 -16767
rect 163637 -16796 163672 -16762
rect 162959 -16861 162960 -16853
rect 162970 -16895 163005 -16861
rect 163192 -16906 163227 -16872
rect 162959 -16961 162960 -16950
rect 162970 -16995 163005 -16961
rect 161907 -17045 161942 -17011
rect 162003 -17045 162038 -17011
rect 162099 -17045 162134 -17011
rect 162608 -17035 162643 -17001
rect 162680 -17035 162715 -17001
rect 162752 -17035 162787 -17001
rect 162824 -17029 162860 -17001
rect 163170 -17025 163205 -16991
rect 163215 -17025 163216 -16980
rect 162824 -17035 162859 -17029
rect 162261 -17088 162296 -17054
rect 162357 -17088 162392 -17054
rect 162453 -17088 162488 -17054
rect 163357 -17076 163358 -16809
rect 163986 -16819 164373 -16753
rect 163373 -16860 163408 -16826
rect 163722 -16832 163733 -16819
rect 163656 -16874 163733 -16832
rect 163784 -16874 164373 -16819
rect 164520 -16853 164555 -16819
rect 164565 -16853 164566 -16808
rect 163656 -16877 164373 -16874
rect 163373 -16928 163408 -16894
rect 163576 -16942 163611 -16908
rect 163621 -16942 163622 -16900
rect 163457 -16991 163458 -16980
rect 163468 -17025 163503 -16991
rect 163576 -17042 163611 -17008
rect 163621 -17042 163622 -16997
rect 163469 -17078 163504 -17044
rect 163541 -17078 163576 -17044
rect 163613 -17078 163648 -17044
rect 162615 -17131 162650 -17097
rect 162711 -17131 162746 -17097
rect 162807 -17131 162842 -17097
rect 162903 -17131 162938 -17097
rect 162999 -17131 163034 -17097
rect 163656 -17114 163801 -16877
rect 163986 -16899 164373 -16877
rect 163910 -16925 164373 -16899
rect 164707 -16904 164708 -16637
rect 164723 -16688 164758 -16654
rect 165337 -16691 165372 -16657
rect 166016 -16663 166051 -16629
rect 166061 -16663 166062 -16618
rect 166161 -16629 166162 -16618
rect 166172 -16663 166207 -16629
rect 166217 -16663 166218 -16618
rect 166317 -16629 166318 -16618
rect 166895 -16623 166930 -16589
rect 167072 -16623 167107 -16589
rect 167433 -16605 167468 -16571
rect 166328 -16663 166363 -16629
rect 166161 -16697 166162 -16671
rect 166560 -16689 166595 -16655
rect 166605 -16689 166606 -16644
rect 166705 -16655 166706 -16644
rect 166716 -16689 166751 -16655
rect 166761 -16689 166762 -16644
rect 167061 -16672 167062 -16661
rect 164723 -16756 164758 -16722
rect 164926 -16770 164961 -16736
rect 164971 -16770 164972 -16728
rect 165071 -16740 165072 -16729
rect 165691 -16734 165726 -16700
rect 165082 -16774 165117 -16740
rect 164807 -16819 164808 -16808
rect 165276 -16813 165311 -16779
rect 165321 -16813 165322 -16771
rect 165421 -16779 165422 -16771
rect 166081 -16777 166116 -16743
rect 165432 -16813 165467 -16779
rect 164818 -16853 164853 -16819
rect 164926 -16870 164961 -16836
rect 164971 -16870 164972 -16825
rect 165071 -16832 165072 -16821
rect 165082 -16866 165117 -16832
rect 165630 -16856 165665 -16822
rect 165675 -16856 165676 -16814
rect 165775 -16822 165776 -16814
rect 165786 -16856 165821 -16822
rect 164819 -16906 164854 -16872
rect 164891 -16906 164926 -16872
rect 164963 -16906 164998 -16872
rect 165276 -16913 165311 -16879
rect 165321 -16913 165322 -16868
rect 165421 -16879 165422 -16868
rect 165432 -16913 165467 -16879
rect 166016 -16895 166051 -16861
rect 166061 -16895 166062 -16853
rect 163910 -16959 164386 -16925
rect 165244 -16949 165279 -16915
rect 165316 -16949 165351 -16915
rect 165630 -16956 165665 -16922
rect 165675 -16956 165676 -16911
rect 165775 -16922 165776 -16911
rect 165786 -16956 165821 -16922
rect 163910 -16985 164373 -16959
rect 163914 -16993 164115 -16985
rect 163930 -17003 164099 -16993
rect 163656 -17140 163831 -17114
rect 163163 -17174 163198 -17140
rect 163259 -17174 163294 -17140
rect 163355 -17174 163390 -17140
rect 163451 -17174 163486 -17140
rect 163547 -17174 163582 -17140
rect 163643 -17174 163831 -17140
rect 163656 -17200 163831 -17174
rect 163856 -17174 163957 -17050
rect 163734 -17870 163769 -17200
rect 163856 -17228 163859 -17174
rect 163541 -17936 163686 -17924
rect 163209 -17970 163686 -17936
rect 163541 -17971 163686 -17970
rect 163722 -17971 163769 -17870
rect 163868 -17971 163903 -17174
rect 164126 -17971 164161 -17062
rect 164260 -17971 164295 -16985
rect 164513 -17002 164548 -16968
rect 164609 -17002 164644 -16968
rect 164705 -17002 164740 -16968
rect 164801 -17002 164836 -16968
rect 164897 -17002 164932 -16968
rect 164993 -17002 165028 -16968
rect 165089 -17002 165124 -16968
rect 165598 -16992 165633 -16958
rect 165670 -16992 165705 -16958
rect 166016 -16995 166051 -16961
rect 166061 -16995 166062 -16950
rect 166203 -17001 166204 -16697
rect 166895 -16706 166930 -16672
rect 167072 -16706 167107 -16672
rect 167368 -16723 167403 -16689
rect 167413 -16723 167414 -16681
rect 167555 -16753 167556 -16525
rect 168245 -16534 168280 -16500
rect 168422 -16534 168457 -16500
rect 168616 -16577 168651 -16543
rect 168661 -16577 168662 -16532
rect 168761 -16543 168762 -16532
rect 168970 -16537 169005 -16503
rect 169015 -16537 169016 -16492
rect 169115 -16503 169116 -16492
rect 169360 -16496 169395 -16462
rect 169405 -16496 169406 -16451
rect 169505 -16462 169506 -16451
rect 169516 -16496 169551 -16462
rect 169561 -16496 169562 -16451
rect 169661 -16462 169662 -16451
rect 169842 -16456 169877 -16422
rect 169914 -16456 169949 -16422
rect 169986 -16456 170021 -16422
rect 170130 -16456 170165 -16422
rect 170202 -16456 170237 -16422
rect 170239 -16456 170309 -16422
rect 170346 -16456 170381 -16422
rect 170416 -16456 170451 -16422
rect 169672 -16496 169707 -16462
rect 170712 -16491 170747 -16457
rect 170757 -16491 170758 -16446
rect 170857 -16457 170858 -16446
rect 170868 -16491 170903 -16457
rect 170913 -16491 170914 -16446
rect 171013 -16457 171014 -16446
rect 171589 -16451 171624 -16417
rect 171766 -16451 171801 -16417
rect 171024 -16491 171059 -16457
rect 169126 -16537 169161 -16503
rect 170405 -16505 170406 -16494
rect 168772 -16577 168807 -16543
rect 167685 -16621 167720 -16587
rect 167886 -16666 167921 -16632
rect 168009 -16637 168010 -16595
rect 168331 -16624 168366 -16590
rect 168970 -16620 169005 -16586
rect 169015 -16620 169016 -16575
rect 169115 -16586 169116 -16575
rect 169360 -16580 169395 -16546
rect 169405 -16580 169406 -16535
rect 169505 -16546 169506 -16535
rect 169516 -16580 169551 -16546
rect 169561 -16580 169562 -16535
rect 169661 -16546 169662 -16535
rect 170239 -16539 170274 -16505
rect 170416 -16539 170451 -16505
rect 169672 -16580 169707 -16546
rect 170559 -16565 170674 -16499
rect 170857 -16525 170858 -16499
rect 171254 -16517 171289 -16483
rect 171299 -16517 171300 -16472
rect 171399 -16483 171400 -16472
rect 171410 -16517 171445 -16483
rect 171455 -16517 171456 -16472
rect 171755 -16500 171756 -16489
rect 171960 -16494 171995 -16460
rect 172005 -16494 172006 -16449
rect 172105 -16460 172106 -16449
rect 172314 -16453 172349 -16419
rect 172359 -16453 172360 -16408
rect 172459 -16419 172460 -16408
rect 172640 -16413 172675 -16379
rect 172704 -16413 172747 -16379
rect 172749 -16413 172750 -16371
rect 172849 -16379 172850 -16371
rect 172784 -16413 172819 -16379
rect 172860 -16413 172895 -16379
rect 172905 -16413 172906 -16371
rect 173005 -16379 173006 -16371
rect 172954 -16413 172989 -16379
rect 173016 -16413 173061 -16379
rect 174056 -16408 174091 -16374
rect 174101 -16408 174102 -16363
rect 174201 -16374 174202 -16363
rect 174212 -16408 174247 -16374
rect 174257 -16408 174258 -16363
rect 174357 -16374 174358 -16363
rect 174933 -16367 174968 -16333
rect 175110 -16367 175145 -16333
rect 175703 -16336 175704 -16328
rect 175803 -16336 175804 -16328
rect 174368 -16408 174403 -16374
rect 172470 -16453 172505 -16419
rect 173749 -16422 173750 -16414
rect 175099 -16417 175100 -16406
rect 175304 -16410 175339 -16376
rect 175349 -16410 175350 -16365
rect 175449 -16376 175450 -16365
rect 175630 -16370 175693 -16336
rect 175702 -16370 175737 -16336
rect 175814 -16370 175849 -16336
rect 176539 -16360 176574 -16326
rect 176635 -16360 176670 -16326
rect 176731 -16360 176766 -16326
rect 176827 -16360 176862 -16326
rect 176923 -16360 176958 -16326
rect 177019 -16360 177054 -16326
rect 177115 -16360 177150 -16326
rect 178443 -16333 178444 -16322
rect 178620 -16327 178683 -16293
rect 178692 -16327 178727 -16293
rect 178804 -16327 178839 -16293
rect 179335 -16317 179370 -16283
rect 179431 -16317 179466 -16283
rect 179527 -16317 179562 -16283
rect 179623 -16317 179658 -16283
rect 179719 -16317 179754 -16283
rect 180744 -16324 180779 -16290
rect 180789 -16324 180790 -16279
rect 180889 -16290 180890 -16279
rect 180900 -16324 180935 -16290
rect 180945 -16324 180946 -16279
rect 181045 -16290 181046 -16279
rect 181224 -16284 181259 -16250
rect 181296 -16284 181331 -16250
rect 181368 -16284 181403 -16250
rect 181512 -16284 181547 -16250
rect 181584 -16284 181619 -16250
rect 181621 -16284 181691 -16250
rect 181728 -16284 181763 -16250
rect 181798 -16284 181833 -16250
rect 182325 -16274 182360 -16240
rect 182421 -16274 182456 -16240
rect 182517 -16274 182552 -16240
rect 184024 -16241 184059 -16207
rect 184088 -16241 184131 -16207
rect 184133 -16241 184134 -16199
rect 184233 -16207 184234 -16199
rect 184168 -16241 184203 -16207
rect 184244 -16241 184279 -16207
rect 184289 -16241 184290 -16199
rect 184389 -16207 184390 -16199
rect 184338 -16241 184373 -16207
rect 184400 -16241 184445 -16207
rect 185315 -16231 185350 -16197
rect 185411 -16231 185446 -16197
rect 185507 -16231 185542 -16197
rect 185131 -16250 185132 -16242
rect 181056 -16324 181091 -16290
rect 182037 -16293 182038 -16285
rect 182137 -16293 182138 -16285
rect 175460 -16410 175495 -16376
rect 172116 -16494 172151 -16460
rect 169126 -16620 169161 -16586
rect 170405 -16589 170406 -16578
rect 167655 -16689 167656 -16681
rect 167666 -16723 167701 -16689
rect 167886 -16734 167921 -16700
rect 166333 -16793 166368 -16759
rect 166536 -16838 166571 -16804
rect 166659 -16809 166660 -16767
rect 166981 -16796 167016 -16762
rect 166303 -16861 166304 -16853
rect 166314 -16895 166349 -16861
rect 166536 -16906 166571 -16872
rect 166303 -16961 166304 -16950
rect 166314 -16995 166349 -16961
rect 165251 -17045 165286 -17011
rect 165347 -17045 165382 -17011
rect 165443 -17045 165478 -17011
rect 165952 -17035 165987 -17001
rect 166024 -17035 166059 -17001
rect 166096 -17035 166131 -17001
rect 166168 -17029 166204 -17001
rect 166514 -17025 166549 -16991
rect 166559 -17025 166560 -16980
rect 166168 -17035 166203 -17029
rect 165605 -17088 165640 -17054
rect 165701 -17088 165736 -17054
rect 165797 -17088 165832 -17054
rect 166701 -17076 166702 -16809
rect 167330 -16819 167717 -16753
rect 166717 -16860 166752 -16826
rect 167066 -16832 167077 -16819
rect 167000 -16874 167077 -16832
rect 167128 -16874 167717 -16819
rect 167864 -16853 167899 -16819
rect 167909 -16853 167910 -16808
rect 167000 -16877 167717 -16874
rect 166717 -16928 166752 -16894
rect 166920 -16942 166955 -16908
rect 166965 -16942 166966 -16900
rect 166801 -16991 166802 -16980
rect 166812 -17025 166847 -16991
rect 166920 -17042 166955 -17008
rect 166965 -17042 166966 -16997
rect 166813 -17078 166848 -17044
rect 166885 -17078 166920 -17044
rect 166957 -17078 166992 -17044
rect 165959 -17131 165994 -17097
rect 166055 -17131 166090 -17097
rect 166151 -17131 166186 -17097
rect 166247 -17131 166282 -17097
rect 166343 -17131 166378 -17097
rect 167000 -17114 167145 -16877
rect 167330 -16899 167717 -16877
rect 167254 -16925 167717 -16899
rect 168051 -16904 168052 -16637
rect 168067 -16688 168102 -16654
rect 168681 -16691 168716 -16657
rect 169360 -16663 169395 -16629
rect 169405 -16663 169406 -16618
rect 169505 -16629 169506 -16618
rect 169516 -16663 169551 -16629
rect 169561 -16663 169562 -16618
rect 169661 -16629 169662 -16618
rect 170239 -16623 170274 -16589
rect 170416 -16623 170451 -16589
rect 170777 -16605 170812 -16571
rect 169672 -16663 169707 -16629
rect 169505 -16697 169506 -16671
rect 169904 -16689 169939 -16655
rect 169949 -16689 169950 -16644
rect 170049 -16655 170050 -16644
rect 170060 -16689 170095 -16655
rect 170105 -16689 170106 -16644
rect 170405 -16672 170406 -16661
rect 168067 -16756 168102 -16722
rect 168270 -16770 168305 -16736
rect 168315 -16770 168316 -16728
rect 168415 -16740 168416 -16729
rect 169035 -16734 169070 -16700
rect 168426 -16774 168461 -16740
rect 168151 -16819 168152 -16808
rect 168620 -16813 168655 -16779
rect 168665 -16813 168666 -16771
rect 168765 -16779 168766 -16771
rect 169425 -16777 169460 -16743
rect 168776 -16813 168811 -16779
rect 168162 -16853 168197 -16819
rect 168270 -16870 168305 -16836
rect 168315 -16870 168316 -16825
rect 168415 -16832 168416 -16821
rect 168426 -16866 168461 -16832
rect 168974 -16856 169009 -16822
rect 169019 -16856 169020 -16814
rect 169119 -16822 169120 -16814
rect 169130 -16856 169165 -16822
rect 168163 -16906 168198 -16872
rect 168235 -16906 168270 -16872
rect 168307 -16906 168342 -16872
rect 168620 -16913 168655 -16879
rect 168665 -16913 168666 -16868
rect 168765 -16879 168766 -16868
rect 168776 -16913 168811 -16879
rect 169360 -16895 169395 -16861
rect 169405 -16895 169406 -16853
rect 167254 -16959 167730 -16925
rect 168588 -16949 168623 -16915
rect 168660 -16949 168695 -16915
rect 168974 -16956 169009 -16922
rect 169019 -16956 169020 -16911
rect 169119 -16922 169120 -16911
rect 169130 -16956 169165 -16922
rect 167254 -16985 167717 -16959
rect 167258 -16993 167459 -16985
rect 167274 -17003 167443 -16993
rect 167000 -17140 167175 -17114
rect 166507 -17174 166542 -17140
rect 166603 -17174 166638 -17140
rect 166699 -17174 166734 -17140
rect 166795 -17174 166830 -17140
rect 166891 -17174 166926 -17140
rect 166987 -17174 167175 -17140
rect 167000 -17200 167175 -17174
rect 167200 -17174 167301 -17050
rect 167078 -17870 167113 -17200
rect 167200 -17228 167203 -17174
rect 166885 -17936 167030 -17924
rect 166553 -17970 167030 -17936
rect 166885 -17971 167030 -17970
rect 167066 -17971 167113 -17870
rect 167212 -17971 167247 -17174
rect 167470 -17971 167505 -17062
rect 167604 -17971 167639 -16985
rect 167857 -17002 167892 -16968
rect 167953 -17002 167988 -16968
rect 168049 -17002 168084 -16968
rect 168145 -17002 168180 -16968
rect 168241 -17002 168276 -16968
rect 168337 -17002 168372 -16968
rect 168433 -17002 168468 -16968
rect 168942 -16992 168977 -16958
rect 169014 -16992 169049 -16958
rect 169360 -16995 169395 -16961
rect 169405 -16995 169406 -16950
rect 169547 -17001 169548 -16697
rect 170239 -16706 170274 -16672
rect 170416 -16706 170451 -16672
rect 170712 -16723 170747 -16689
rect 170757 -16723 170758 -16681
rect 170899 -16753 170900 -16525
rect 171589 -16534 171624 -16500
rect 171766 -16534 171801 -16500
rect 171960 -16577 171995 -16543
rect 172005 -16577 172006 -16532
rect 172105 -16543 172106 -16532
rect 172314 -16537 172349 -16503
rect 172359 -16537 172360 -16492
rect 172459 -16503 172460 -16492
rect 172704 -16496 172739 -16462
rect 172749 -16496 172750 -16451
rect 172849 -16462 172850 -16451
rect 172860 -16496 172895 -16462
rect 172905 -16496 172906 -16451
rect 173005 -16462 173006 -16451
rect 173186 -16456 173221 -16422
rect 173258 -16456 173293 -16422
rect 173330 -16456 173365 -16422
rect 173474 -16456 173509 -16422
rect 173546 -16456 173581 -16422
rect 173583 -16456 173653 -16422
rect 173690 -16456 173725 -16422
rect 173760 -16456 173795 -16422
rect 173016 -16496 173051 -16462
rect 174056 -16491 174091 -16457
rect 174101 -16491 174102 -16446
rect 174201 -16457 174202 -16446
rect 174212 -16491 174247 -16457
rect 174257 -16491 174258 -16446
rect 174357 -16457 174358 -16446
rect 174933 -16451 174968 -16417
rect 175110 -16451 175145 -16417
rect 174368 -16491 174403 -16457
rect 172470 -16537 172505 -16503
rect 173749 -16505 173750 -16494
rect 172116 -16577 172151 -16543
rect 171029 -16621 171064 -16587
rect 171230 -16666 171265 -16632
rect 171353 -16637 171354 -16595
rect 171675 -16624 171710 -16590
rect 172314 -16620 172349 -16586
rect 172359 -16620 172360 -16575
rect 172459 -16586 172460 -16575
rect 172704 -16580 172739 -16546
rect 172749 -16580 172750 -16535
rect 172849 -16546 172850 -16535
rect 172860 -16580 172895 -16546
rect 172905 -16580 172906 -16535
rect 173005 -16546 173006 -16535
rect 173583 -16539 173618 -16505
rect 173760 -16539 173795 -16505
rect 173016 -16580 173051 -16546
rect 173903 -16565 174018 -16499
rect 174201 -16525 174202 -16499
rect 174598 -16517 174633 -16483
rect 174643 -16517 174644 -16472
rect 174743 -16483 174744 -16472
rect 174754 -16517 174789 -16483
rect 174799 -16517 174800 -16472
rect 175099 -16500 175100 -16489
rect 175304 -16494 175339 -16460
rect 175349 -16494 175350 -16449
rect 175449 -16460 175450 -16449
rect 175658 -16453 175693 -16419
rect 175703 -16453 175704 -16408
rect 175803 -16419 175804 -16408
rect 175984 -16413 176019 -16379
rect 176048 -16413 176091 -16379
rect 176093 -16413 176094 -16371
rect 176193 -16379 176194 -16371
rect 176128 -16413 176163 -16379
rect 176204 -16413 176239 -16379
rect 176249 -16413 176250 -16371
rect 176349 -16379 176350 -16371
rect 176298 -16413 176333 -16379
rect 176360 -16413 176405 -16379
rect 177400 -16408 177435 -16374
rect 177445 -16408 177446 -16363
rect 177545 -16374 177546 -16363
rect 177556 -16408 177591 -16374
rect 177601 -16408 177602 -16363
rect 177701 -16374 177702 -16363
rect 178277 -16367 178312 -16333
rect 178454 -16367 178489 -16333
rect 179047 -16336 179048 -16328
rect 179147 -16336 179148 -16328
rect 177712 -16408 177747 -16374
rect 175814 -16453 175849 -16419
rect 177093 -16422 177094 -16414
rect 178443 -16417 178444 -16406
rect 178648 -16410 178683 -16376
rect 178693 -16410 178694 -16365
rect 178793 -16376 178794 -16365
rect 178974 -16370 179037 -16336
rect 179046 -16370 179081 -16336
rect 179158 -16370 179193 -16336
rect 179883 -16360 179918 -16326
rect 179979 -16360 180014 -16326
rect 180075 -16360 180110 -16326
rect 180171 -16360 180206 -16326
rect 180267 -16360 180302 -16326
rect 180363 -16360 180398 -16326
rect 180459 -16360 180494 -16326
rect 181787 -16333 181788 -16322
rect 181964 -16327 182027 -16293
rect 182036 -16327 182071 -16293
rect 182148 -16327 182183 -16293
rect 182679 -16317 182714 -16283
rect 182775 -16317 182810 -16283
rect 182871 -16317 182906 -16283
rect 182967 -16317 183002 -16283
rect 183063 -16317 183098 -16283
rect 184088 -16324 184123 -16290
rect 184133 -16324 184134 -16279
rect 184233 -16290 184234 -16279
rect 184244 -16324 184279 -16290
rect 184289 -16324 184290 -16279
rect 184389 -16290 184390 -16279
rect 184568 -16284 184603 -16250
rect 184640 -16284 184675 -16250
rect 184712 -16284 184747 -16250
rect 184856 -16284 184891 -16250
rect 184928 -16284 184963 -16250
rect 184965 -16284 185035 -16250
rect 185072 -16284 185107 -16250
rect 185142 -16284 185177 -16250
rect 185669 -16274 185704 -16240
rect 185765 -16274 185800 -16240
rect 185861 -16274 185896 -16240
rect 187368 -16241 187403 -16207
rect 187432 -16241 187475 -16207
rect 187477 -16241 187478 -16199
rect 187577 -16207 187578 -16199
rect 187512 -16241 187547 -16207
rect 187588 -16241 187623 -16207
rect 187633 -16241 187634 -16199
rect 187733 -16207 187734 -16199
rect 187682 -16241 187717 -16207
rect 187744 -16241 187789 -16207
rect 188659 -16231 188694 -16197
rect 188755 -16231 188790 -16197
rect 188851 -16231 188886 -16197
rect 188475 -16250 188476 -16242
rect 184400 -16324 184435 -16290
rect 185381 -16293 185382 -16285
rect 185481 -16293 185482 -16285
rect 178804 -16410 178839 -16376
rect 175460 -16494 175495 -16460
rect 172470 -16620 172505 -16586
rect 173749 -16589 173750 -16578
rect 170999 -16689 171000 -16681
rect 171010 -16723 171045 -16689
rect 171230 -16734 171265 -16700
rect 169677 -16793 169712 -16759
rect 169880 -16838 169915 -16804
rect 170003 -16809 170004 -16767
rect 170325 -16796 170360 -16762
rect 169647 -16861 169648 -16853
rect 169658 -16895 169693 -16861
rect 169880 -16906 169915 -16872
rect 169647 -16961 169648 -16950
rect 169658 -16995 169693 -16961
rect 168595 -17045 168630 -17011
rect 168691 -17045 168726 -17011
rect 168787 -17045 168822 -17011
rect 169296 -17035 169331 -17001
rect 169368 -17035 169403 -17001
rect 169440 -17035 169475 -17001
rect 169512 -17029 169548 -17001
rect 169858 -17025 169893 -16991
rect 169903 -17025 169904 -16980
rect 169512 -17035 169547 -17029
rect 168949 -17088 168984 -17054
rect 169045 -17088 169080 -17054
rect 169141 -17088 169176 -17054
rect 170045 -17076 170046 -16809
rect 170674 -16819 171061 -16753
rect 170061 -16860 170096 -16826
rect 170410 -16832 170421 -16819
rect 170344 -16874 170421 -16832
rect 170472 -16874 171061 -16819
rect 171208 -16853 171243 -16819
rect 171253 -16853 171254 -16808
rect 170344 -16877 171061 -16874
rect 170061 -16928 170096 -16894
rect 170264 -16942 170299 -16908
rect 170309 -16942 170310 -16900
rect 170145 -16991 170146 -16980
rect 170156 -17025 170191 -16991
rect 170264 -17042 170299 -17008
rect 170309 -17042 170310 -16997
rect 170157 -17078 170192 -17044
rect 170229 -17078 170264 -17044
rect 170301 -17078 170336 -17044
rect 169303 -17131 169338 -17097
rect 169399 -17131 169434 -17097
rect 169495 -17131 169530 -17097
rect 169591 -17131 169626 -17097
rect 169687 -17131 169722 -17097
rect 170344 -17114 170489 -16877
rect 170674 -16899 171061 -16877
rect 170598 -16925 171061 -16899
rect 171395 -16904 171396 -16637
rect 171411 -16688 171446 -16654
rect 172025 -16691 172060 -16657
rect 172704 -16663 172739 -16629
rect 172749 -16663 172750 -16618
rect 172849 -16629 172850 -16618
rect 172860 -16663 172895 -16629
rect 172905 -16663 172906 -16618
rect 173005 -16629 173006 -16618
rect 173583 -16623 173618 -16589
rect 173760 -16623 173795 -16589
rect 174121 -16605 174156 -16571
rect 173016 -16663 173051 -16629
rect 172849 -16697 172850 -16671
rect 173248 -16689 173283 -16655
rect 173293 -16689 173294 -16644
rect 173393 -16655 173394 -16644
rect 173404 -16689 173439 -16655
rect 173449 -16689 173450 -16644
rect 173749 -16672 173750 -16661
rect 171411 -16756 171446 -16722
rect 171614 -16770 171649 -16736
rect 171659 -16770 171660 -16728
rect 171759 -16740 171760 -16729
rect 172379 -16734 172414 -16700
rect 171770 -16774 171805 -16740
rect 171495 -16819 171496 -16808
rect 171964 -16813 171999 -16779
rect 172009 -16813 172010 -16771
rect 172109 -16779 172110 -16771
rect 172769 -16777 172804 -16743
rect 172120 -16813 172155 -16779
rect 171506 -16853 171541 -16819
rect 171614 -16870 171649 -16836
rect 171659 -16870 171660 -16825
rect 171759 -16832 171760 -16821
rect 171770 -16866 171805 -16832
rect 172318 -16856 172353 -16822
rect 172363 -16856 172364 -16814
rect 172463 -16822 172464 -16814
rect 172474 -16856 172509 -16822
rect 171507 -16906 171542 -16872
rect 171579 -16906 171614 -16872
rect 171651 -16906 171686 -16872
rect 171964 -16913 171999 -16879
rect 172009 -16913 172010 -16868
rect 172109 -16879 172110 -16868
rect 172120 -16913 172155 -16879
rect 172704 -16895 172739 -16861
rect 172749 -16895 172750 -16853
rect 170598 -16959 171074 -16925
rect 171932 -16949 171967 -16915
rect 172004 -16949 172039 -16915
rect 172318 -16956 172353 -16922
rect 172363 -16956 172364 -16911
rect 172463 -16922 172464 -16911
rect 172474 -16956 172509 -16922
rect 170598 -16985 171061 -16959
rect 170602 -16993 170803 -16985
rect 170618 -17003 170787 -16993
rect 170344 -17140 170519 -17114
rect 169851 -17174 169886 -17140
rect 169947 -17174 169982 -17140
rect 170043 -17174 170078 -17140
rect 170139 -17174 170174 -17140
rect 170235 -17174 170270 -17140
rect 170331 -17174 170519 -17140
rect 170344 -17200 170519 -17174
rect 170544 -17174 170645 -17050
rect 170422 -17870 170457 -17200
rect 170544 -17228 170547 -17174
rect 170229 -17936 170374 -17924
rect 169897 -17970 170374 -17936
rect 170229 -17971 170374 -17970
rect 170410 -17971 170457 -17870
rect 170556 -17971 170591 -17174
rect 170814 -17971 170849 -17062
rect 170948 -17971 170983 -16985
rect 171201 -17002 171236 -16968
rect 171297 -17002 171332 -16968
rect 171393 -17002 171428 -16968
rect 171489 -17002 171524 -16968
rect 171585 -17002 171620 -16968
rect 171681 -17002 171716 -16968
rect 171777 -17002 171812 -16968
rect 172286 -16992 172321 -16958
rect 172358 -16992 172393 -16958
rect 172704 -16995 172739 -16961
rect 172749 -16995 172750 -16950
rect 172891 -17001 172892 -16697
rect 173583 -16706 173618 -16672
rect 173760 -16706 173795 -16672
rect 174056 -16723 174091 -16689
rect 174101 -16723 174102 -16681
rect 174243 -16753 174244 -16525
rect 174933 -16534 174968 -16500
rect 175110 -16534 175145 -16500
rect 175304 -16577 175339 -16543
rect 175349 -16577 175350 -16532
rect 175449 -16543 175450 -16532
rect 175658 -16537 175693 -16503
rect 175703 -16537 175704 -16492
rect 175803 -16503 175804 -16492
rect 176048 -16496 176083 -16462
rect 176093 -16496 176094 -16451
rect 176193 -16462 176194 -16451
rect 176204 -16496 176239 -16462
rect 176249 -16496 176250 -16451
rect 176349 -16462 176350 -16451
rect 176530 -16456 176565 -16422
rect 176602 -16456 176637 -16422
rect 176674 -16456 176709 -16422
rect 176818 -16456 176853 -16422
rect 176890 -16456 176925 -16422
rect 176927 -16456 176997 -16422
rect 177034 -16456 177069 -16422
rect 177104 -16456 177139 -16422
rect 176360 -16496 176395 -16462
rect 177400 -16491 177435 -16457
rect 177445 -16491 177446 -16446
rect 177545 -16457 177546 -16446
rect 177556 -16491 177591 -16457
rect 177601 -16491 177602 -16446
rect 177701 -16457 177702 -16446
rect 178277 -16451 178312 -16417
rect 178454 -16451 178489 -16417
rect 177712 -16491 177747 -16457
rect 175814 -16537 175849 -16503
rect 177093 -16505 177094 -16494
rect 175460 -16577 175495 -16543
rect 174373 -16621 174408 -16587
rect 174574 -16666 174609 -16632
rect 174697 -16637 174698 -16595
rect 175019 -16624 175054 -16590
rect 175658 -16620 175693 -16586
rect 175703 -16620 175704 -16575
rect 175803 -16586 175804 -16575
rect 176048 -16580 176083 -16546
rect 176093 -16580 176094 -16535
rect 176193 -16546 176194 -16535
rect 176204 -16580 176239 -16546
rect 176249 -16580 176250 -16535
rect 176349 -16546 176350 -16535
rect 176927 -16539 176962 -16505
rect 177104 -16539 177139 -16505
rect 176360 -16580 176395 -16546
rect 177247 -16565 177362 -16499
rect 177545 -16525 177546 -16499
rect 177942 -16517 177977 -16483
rect 177987 -16517 177988 -16472
rect 178087 -16483 178088 -16472
rect 178098 -16517 178133 -16483
rect 178143 -16517 178144 -16472
rect 178443 -16500 178444 -16489
rect 178648 -16494 178683 -16460
rect 178693 -16494 178694 -16449
rect 178793 -16460 178794 -16449
rect 179002 -16453 179037 -16419
rect 179047 -16453 179048 -16408
rect 179147 -16419 179148 -16408
rect 179328 -16413 179363 -16379
rect 179392 -16413 179435 -16379
rect 179437 -16413 179438 -16371
rect 179537 -16379 179538 -16371
rect 179472 -16413 179507 -16379
rect 179548 -16413 179583 -16379
rect 179593 -16413 179594 -16371
rect 179693 -16379 179694 -16371
rect 179642 -16413 179677 -16379
rect 179704 -16413 179749 -16379
rect 180744 -16408 180779 -16374
rect 180789 -16408 180790 -16363
rect 180889 -16374 180890 -16363
rect 180900 -16408 180935 -16374
rect 180945 -16408 180946 -16363
rect 181045 -16374 181046 -16363
rect 181621 -16367 181656 -16333
rect 181798 -16367 181833 -16333
rect 182391 -16336 182392 -16328
rect 182491 -16336 182492 -16328
rect 181056 -16408 181091 -16374
rect 179158 -16453 179193 -16419
rect 180437 -16422 180438 -16414
rect 181787 -16417 181788 -16406
rect 181992 -16410 182027 -16376
rect 182037 -16410 182038 -16365
rect 182137 -16376 182138 -16365
rect 182318 -16370 182381 -16336
rect 182390 -16370 182425 -16336
rect 182502 -16370 182537 -16336
rect 183227 -16360 183262 -16326
rect 183323 -16360 183358 -16326
rect 183419 -16360 183454 -16326
rect 183515 -16360 183550 -16326
rect 183611 -16360 183646 -16326
rect 183707 -16360 183742 -16326
rect 183803 -16360 183838 -16326
rect 185131 -16333 185132 -16322
rect 185308 -16327 185371 -16293
rect 185380 -16327 185415 -16293
rect 185492 -16327 185527 -16293
rect 186023 -16317 186058 -16283
rect 186119 -16317 186154 -16283
rect 186215 -16317 186250 -16283
rect 186311 -16317 186346 -16283
rect 186407 -16317 186442 -16283
rect 187432 -16324 187467 -16290
rect 187477 -16324 187478 -16279
rect 187577 -16290 187578 -16279
rect 187588 -16324 187623 -16290
rect 187633 -16324 187634 -16279
rect 187733 -16290 187734 -16279
rect 187912 -16284 187947 -16250
rect 187984 -16284 188019 -16250
rect 188056 -16284 188091 -16250
rect 188200 -16284 188235 -16250
rect 188272 -16284 188307 -16250
rect 188309 -16284 188379 -16250
rect 188416 -16284 188451 -16250
rect 188486 -16284 188521 -16250
rect 189013 -16274 189048 -16240
rect 189109 -16274 189144 -16240
rect 189205 -16274 189240 -16240
rect 190712 -16241 190747 -16207
rect 190776 -16241 190819 -16207
rect 190821 -16241 190822 -16199
rect 190921 -16207 190922 -16199
rect 190856 -16241 190891 -16207
rect 190932 -16241 190967 -16207
rect 190977 -16241 190978 -16199
rect 191077 -16207 191078 -16199
rect 191026 -16241 191061 -16207
rect 191088 -16241 191133 -16207
rect 192003 -16231 192038 -16197
rect 192099 -16231 192134 -16197
rect 192195 -16231 192230 -16197
rect 191819 -16250 191820 -16242
rect 187744 -16324 187779 -16290
rect 188725 -16293 188726 -16285
rect 188825 -16293 188826 -16285
rect 182148 -16410 182183 -16376
rect 178804 -16494 178839 -16460
rect 175814 -16620 175849 -16586
rect 177093 -16589 177094 -16578
rect 174343 -16689 174344 -16681
rect 174354 -16723 174389 -16689
rect 174574 -16734 174609 -16700
rect 173021 -16793 173056 -16759
rect 173224 -16838 173259 -16804
rect 173347 -16809 173348 -16767
rect 173669 -16796 173704 -16762
rect 172991 -16861 172992 -16853
rect 173002 -16895 173037 -16861
rect 173224 -16906 173259 -16872
rect 172991 -16961 172992 -16950
rect 173002 -16995 173037 -16961
rect 171939 -17045 171974 -17011
rect 172035 -17045 172070 -17011
rect 172131 -17045 172166 -17011
rect 172640 -17035 172675 -17001
rect 172712 -17035 172747 -17001
rect 172784 -17035 172819 -17001
rect 172856 -17029 172892 -17001
rect 173202 -17025 173237 -16991
rect 173247 -17025 173248 -16980
rect 172856 -17035 172891 -17029
rect 172293 -17088 172328 -17054
rect 172389 -17088 172424 -17054
rect 172485 -17088 172520 -17054
rect 173389 -17076 173390 -16809
rect 174018 -16819 174405 -16753
rect 173405 -16860 173440 -16826
rect 173754 -16832 173765 -16819
rect 173688 -16874 173765 -16832
rect 173816 -16874 174405 -16819
rect 174552 -16853 174587 -16819
rect 174597 -16853 174598 -16808
rect 173688 -16877 174405 -16874
rect 173405 -16928 173440 -16894
rect 173608 -16942 173643 -16908
rect 173653 -16942 173654 -16900
rect 173489 -16991 173490 -16980
rect 173500 -17025 173535 -16991
rect 173608 -17042 173643 -17008
rect 173653 -17042 173654 -16997
rect 173501 -17078 173536 -17044
rect 173573 -17078 173608 -17044
rect 173645 -17078 173680 -17044
rect 172647 -17131 172682 -17097
rect 172743 -17131 172778 -17097
rect 172839 -17131 172874 -17097
rect 172935 -17131 172970 -17097
rect 173031 -17131 173066 -17097
rect 173688 -17114 173833 -16877
rect 174018 -16899 174405 -16877
rect 173942 -16925 174405 -16899
rect 174739 -16904 174740 -16637
rect 174755 -16688 174790 -16654
rect 175369 -16691 175404 -16657
rect 176048 -16663 176083 -16629
rect 176093 -16663 176094 -16618
rect 176193 -16629 176194 -16618
rect 176204 -16663 176239 -16629
rect 176249 -16663 176250 -16618
rect 176349 -16629 176350 -16618
rect 176927 -16623 176962 -16589
rect 177104 -16623 177139 -16589
rect 177465 -16605 177500 -16571
rect 176360 -16663 176395 -16629
rect 176193 -16697 176194 -16671
rect 176592 -16689 176627 -16655
rect 176637 -16689 176638 -16644
rect 176737 -16655 176738 -16644
rect 176748 -16689 176783 -16655
rect 176793 -16689 176794 -16644
rect 177093 -16672 177094 -16661
rect 174755 -16756 174790 -16722
rect 174958 -16770 174993 -16736
rect 175003 -16770 175004 -16728
rect 175103 -16740 175104 -16729
rect 175723 -16734 175758 -16700
rect 175114 -16774 175149 -16740
rect 174839 -16819 174840 -16808
rect 175308 -16813 175343 -16779
rect 175353 -16813 175354 -16771
rect 175453 -16779 175454 -16771
rect 176113 -16777 176148 -16743
rect 175464 -16813 175499 -16779
rect 174850 -16853 174885 -16819
rect 174958 -16870 174993 -16836
rect 175003 -16870 175004 -16825
rect 175103 -16832 175104 -16821
rect 175114 -16866 175149 -16832
rect 175662 -16856 175697 -16822
rect 175707 -16856 175708 -16814
rect 175807 -16822 175808 -16814
rect 175818 -16856 175853 -16822
rect 174851 -16906 174886 -16872
rect 174923 -16906 174958 -16872
rect 174995 -16906 175030 -16872
rect 175308 -16913 175343 -16879
rect 175353 -16913 175354 -16868
rect 175453 -16879 175454 -16868
rect 175464 -16913 175499 -16879
rect 176048 -16895 176083 -16861
rect 176093 -16895 176094 -16853
rect 173942 -16959 174418 -16925
rect 175276 -16949 175311 -16915
rect 175348 -16949 175383 -16915
rect 175662 -16956 175697 -16922
rect 175707 -16956 175708 -16911
rect 175807 -16922 175808 -16911
rect 175818 -16956 175853 -16922
rect 173942 -16985 174405 -16959
rect 173946 -16993 174147 -16985
rect 173962 -17003 174131 -16993
rect 173688 -17140 173863 -17114
rect 173195 -17174 173230 -17140
rect 173291 -17174 173326 -17140
rect 173387 -17174 173422 -17140
rect 173483 -17174 173518 -17140
rect 173579 -17174 173614 -17140
rect 173675 -17174 173863 -17140
rect 173688 -17200 173863 -17174
rect 173888 -17174 173989 -17050
rect 173766 -17870 173801 -17200
rect 173888 -17228 173891 -17174
rect 173573 -17936 173718 -17924
rect 173241 -17970 173718 -17936
rect 173573 -17971 173718 -17970
rect 173754 -17971 173801 -17870
rect 173900 -17971 173935 -17174
rect 174158 -17971 174193 -17062
rect 174292 -17971 174327 -16985
rect 174545 -17002 174580 -16968
rect 174641 -17002 174676 -16968
rect 174737 -17002 174772 -16968
rect 174833 -17002 174868 -16968
rect 174929 -17002 174964 -16968
rect 175025 -17002 175060 -16968
rect 175121 -17002 175156 -16968
rect 175630 -16992 175665 -16958
rect 175702 -16992 175737 -16958
rect 176048 -16995 176083 -16961
rect 176093 -16995 176094 -16950
rect 176235 -17001 176236 -16697
rect 176927 -16706 176962 -16672
rect 177104 -16706 177139 -16672
rect 177400 -16723 177435 -16689
rect 177445 -16723 177446 -16681
rect 177587 -16753 177588 -16525
rect 178277 -16534 178312 -16500
rect 178454 -16534 178489 -16500
rect 178648 -16577 178683 -16543
rect 178693 -16577 178694 -16532
rect 178793 -16543 178794 -16532
rect 179002 -16537 179037 -16503
rect 179047 -16537 179048 -16492
rect 179147 -16503 179148 -16492
rect 179392 -16496 179427 -16462
rect 179437 -16496 179438 -16451
rect 179537 -16462 179538 -16451
rect 179548 -16496 179583 -16462
rect 179593 -16496 179594 -16451
rect 179693 -16462 179694 -16451
rect 179874 -16456 179909 -16422
rect 179946 -16456 179981 -16422
rect 180018 -16456 180053 -16422
rect 180162 -16456 180197 -16422
rect 180234 -16456 180269 -16422
rect 180271 -16456 180341 -16422
rect 180378 -16456 180413 -16422
rect 180448 -16456 180483 -16422
rect 179704 -16496 179739 -16462
rect 180744 -16491 180779 -16457
rect 180789 -16491 180790 -16446
rect 180889 -16457 180890 -16446
rect 180900 -16491 180935 -16457
rect 180945 -16491 180946 -16446
rect 181045 -16457 181046 -16446
rect 181621 -16451 181656 -16417
rect 181798 -16451 181833 -16417
rect 181056 -16491 181091 -16457
rect 179158 -16537 179193 -16503
rect 180437 -16505 180438 -16494
rect 178804 -16577 178839 -16543
rect 177717 -16621 177752 -16587
rect 177918 -16666 177953 -16632
rect 178041 -16637 178042 -16595
rect 178363 -16624 178398 -16590
rect 179002 -16620 179037 -16586
rect 179047 -16620 179048 -16575
rect 179147 -16586 179148 -16575
rect 179392 -16580 179427 -16546
rect 179437 -16580 179438 -16535
rect 179537 -16546 179538 -16535
rect 179548 -16580 179583 -16546
rect 179593 -16580 179594 -16535
rect 179693 -16546 179694 -16535
rect 180271 -16539 180306 -16505
rect 180448 -16539 180483 -16505
rect 179704 -16580 179739 -16546
rect 180591 -16565 180706 -16499
rect 180889 -16525 180890 -16499
rect 181286 -16517 181321 -16483
rect 181331 -16517 181332 -16472
rect 181431 -16483 181432 -16472
rect 181442 -16517 181477 -16483
rect 181487 -16517 181488 -16472
rect 181787 -16500 181788 -16489
rect 181992 -16494 182027 -16460
rect 182037 -16494 182038 -16449
rect 182137 -16460 182138 -16449
rect 182346 -16453 182381 -16419
rect 182391 -16453 182392 -16408
rect 182491 -16419 182492 -16408
rect 182672 -16413 182707 -16379
rect 182736 -16413 182779 -16379
rect 182781 -16413 182782 -16371
rect 182881 -16379 182882 -16371
rect 182816 -16413 182851 -16379
rect 182892 -16413 182927 -16379
rect 182937 -16413 182938 -16371
rect 183037 -16379 183038 -16371
rect 182986 -16413 183021 -16379
rect 183048 -16413 183093 -16379
rect 184088 -16408 184123 -16374
rect 184133 -16408 184134 -16363
rect 184233 -16374 184234 -16363
rect 184244 -16408 184279 -16374
rect 184289 -16408 184290 -16363
rect 184389 -16374 184390 -16363
rect 184965 -16367 185000 -16333
rect 185142 -16367 185177 -16333
rect 185735 -16336 185736 -16328
rect 185835 -16336 185836 -16328
rect 184400 -16408 184435 -16374
rect 182502 -16453 182537 -16419
rect 183781 -16422 183782 -16414
rect 185131 -16417 185132 -16406
rect 185336 -16410 185371 -16376
rect 185381 -16410 185382 -16365
rect 185481 -16376 185482 -16365
rect 185662 -16370 185725 -16336
rect 185734 -16370 185769 -16336
rect 185846 -16370 185881 -16336
rect 186571 -16360 186606 -16326
rect 186667 -16360 186702 -16326
rect 186763 -16360 186798 -16326
rect 186859 -16360 186894 -16326
rect 186955 -16360 186990 -16326
rect 187051 -16360 187086 -16326
rect 187147 -16360 187182 -16326
rect 188475 -16333 188476 -16322
rect 188652 -16327 188715 -16293
rect 188724 -16327 188759 -16293
rect 188836 -16327 188871 -16293
rect 189367 -16317 189402 -16283
rect 189463 -16317 189498 -16283
rect 189559 -16317 189594 -16283
rect 189655 -16317 189690 -16283
rect 189751 -16317 189786 -16283
rect 190776 -16324 190811 -16290
rect 190821 -16324 190822 -16279
rect 190921 -16290 190922 -16279
rect 190932 -16324 190967 -16290
rect 190977 -16324 190978 -16279
rect 191077 -16290 191078 -16279
rect 191256 -16284 191291 -16250
rect 191328 -16284 191363 -16250
rect 191400 -16284 191435 -16250
rect 191544 -16284 191579 -16250
rect 191616 -16284 191651 -16250
rect 191653 -16284 191723 -16250
rect 191760 -16284 191795 -16250
rect 191830 -16284 191865 -16250
rect 192357 -16274 192392 -16240
rect 192453 -16274 192488 -16240
rect 192549 -16274 192584 -16240
rect 194056 -16241 194091 -16207
rect 194120 -16241 194163 -16207
rect 194165 -16241 194166 -16199
rect 194265 -16207 194266 -16199
rect 194200 -16241 194235 -16207
rect 194276 -16241 194311 -16207
rect 194321 -16241 194322 -16199
rect 194421 -16207 194422 -16199
rect 194370 -16241 194405 -16207
rect 194432 -16241 194477 -16207
rect 195347 -16231 195382 -16197
rect 195443 -16231 195478 -16197
rect 195539 -16231 195574 -16197
rect 195163 -16250 195164 -16242
rect 191088 -16324 191123 -16290
rect 192069 -16293 192070 -16285
rect 192169 -16293 192170 -16285
rect 185492 -16410 185527 -16376
rect 182148 -16494 182183 -16460
rect 179158 -16620 179193 -16586
rect 180437 -16589 180438 -16578
rect 177687 -16689 177688 -16681
rect 177698 -16723 177733 -16689
rect 177918 -16734 177953 -16700
rect 176365 -16793 176400 -16759
rect 176568 -16838 176603 -16804
rect 176691 -16809 176692 -16767
rect 177013 -16796 177048 -16762
rect 176335 -16861 176336 -16853
rect 176346 -16895 176381 -16861
rect 176568 -16906 176603 -16872
rect 176335 -16961 176336 -16950
rect 176346 -16995 176381 -16961
rect 175283 -17045 175318 -17011
rect 175379 -17045 175414 -17011
rect 175475 -17045 175510 -17011
rect 175984 -17035 176019 -17001
rect 176056 -17035 176091 -17001
rect 176128 -17035 176163 -17001
rect 176200 -17029 176236 -17001
rect 176546 -17025 176581 -16991
rect 176591 -17025 176592 -16980
rect 176200 -17035 176235 -17029
rect 175637 -17088 175672 -17054
rect 175733 -17088 175768 -17054
rect 175829 -17088 175864 -17054
rect 176733 -17076 176734 -16809
rect 177362 -16819 177749 -16753
rect 176749 -16860 176784 -16826
rect 177098 -16832 177109 -16819
rect 177032 -16874 177109 -16832
rect 177160 -16874 177749 -16819
rect 177896 -16853 177931 -16819
rect 177941 -16853 177942 -16808
rect 177032 -16877 177749 -16874
rect 176749 -16928 176784 -16894
rect 176952 -16942 176987 -16908
rect 176997 -16942 176998 -16900
rect 176833 -16991 176834 -16980
rect 176844 -17025 176879 -16991
rect 176952 -17042 176987 -17008
rect 176997 -17042 176998 -16997
rect 176845 -17078 176880 -17044
rect 176917 -17078 176952 -17044
rect 176989 -17078 177024 -17044
rect 175991 -17131 176026 -17097
rect 176087 -17131 176122 -17097
rect 176183 -17131 176218 -17097
rect 176279 -17131 176314 -17097
rect 176375 -17131 176410 -17097
rect 177032 -17114 177177 -16877
rect 177362 -16899 177749 -16877
rect 177286 -16925 177749 -16899
rect 178083 -16904 178084 -16637
rect 178099 -16688 178134 -16654
rect 178713 -16691 178748 -16657
rect 179392 -16663 179427 -16629
rect 179437 -16663 179438 -16618
rect 179537 -16629 179538 -16618
rect 179548 -16663 179583 -16629
rect 179593 -16663 179594 -16618
rect 179693 -16629 179694 -16618
rect 180271 -16623 180306 -16589
rect 180448 -16623 180483 -16589
rect 180809 -16605 180844 -16571
rect 179704 -16663 179739 -16629
rect 179537 -16697 179538 -16671
rect 179936 -16689 179971 -16655
rect 179981 -16689 179982 -16644
rect 180081 -16655 180082 -16644
rect 180092 -16689 180127 -16655
rect 180137 -16689 180138 -16644
rect 180437 -16672 180438 -16661
rect 178099 -16756 178134 -16722
rect 178302 -16770 178337 -16736
rect 178347 -16770 178348 -16728
rect 178447 -16740 178448 -16729
rect 179067 -16734 179102 -16700
rect 178458 -16774 178493 -16740
rect 178183 -16819 178184 -16808
rect 178652 -16813 178687 -16779
rect 178697 -16813 178698 -16771
rect 178797 -16779 178798 -16771
rect 179457 -16777 179492 -16743
rect 178808 -16813 178843 -16779
rect 178194 -16853 178229 -16819
rect 178302 -16870 178337 -16836
rect 178347 -16870 178348 -16825
rect 178447 -16832 178448 -16821
rect 178458 -16866 178493 -16832
rect 179006 -16856 179041 -16822
rect 179051 -16856 179052 -16814
rect 179151 -16822 179152 -16814
rect 179162 -16856 179197 -16822
rect 178195 -16906 178230 -16872
rect 178267 -16906 178302 -16872
rect 178339 -16906 178374 -16872
rect 178652 -16913 178687 -16879
rect 178697 -16913 178698 -16868
rect 178797 -16879 178798 -16868
rect 178808 -16913 178843 -16879
rect 179392 -16895 179427 -16861
rect 179437 -16895 179438 -16853
rect 177286 -16959 177762 -16925
rect 178620 -16949 178655 -16915
rect 178692 -16949 178727 -16915
rect 179006 -16956 179041 -16922
rect 179051 -16956 179052 -16911
rect 179151 -16922 179152 -16911
rect 179162 -16956 179197 -16922
rect 177286 -16985 177749 -16959
rect 177290 -16993 177491 -16985
rect 177306 -17003 177475 -16993
rect 177032 -17140 177207 -17114
rect 176539 -17174 176574 -17140
rect 176635 -17174 176670 -17140
rect 176731 -17174 176766 -17140
rect 176827 -17174 176862 -17140
rect 176923 -17174 176958 -17140
rect 177019 -17174 177207 -17140
rect 177032 -17200 177207 -17174
rect 177232 -17174 177333 -17050
rect 177110 -17870 177145 -17200
rect 177232 -17228 177235 -17174
rect 176917 -17936 177062 -17924
rect 176585 -17970 177062 -17936
rect 176917 -17971 177062 -17970
rect 177098 -17971 177145 -17870
rect 177244 -17971 177279 -17174
rect 177502 -17971 177537 -17062
rect 177636 -17971 177671 -16985
rect 177889 -17002 177924 -16968
rect 177985 -17002 178020 -16968
rect 178081 -17002 178116 -16968
rect 178177 -17002 178212 -16968
rect 178273 -17002 178308 -16968
rect 178369 -17002 178404 -16968
rect 178465 -17002 178500 -16968
rect 178974 -16992 179009 -16958
rect 179046 -16992 179081 -16958
rect 179392 -16995 179427 -16961
rect 179437 -16995 179438 -16950
rect 179579 -17001 179580 -16697
rect 180271 -16706 180306 -16672
rect 180448 -16706 180483 -16672
rect 180744 -16723 180779 -16689
rect 180789 -16723 180790 -16681
rect 180931 -16753 180932 -16525
rect 181621 -16534 181656 -16500
rect 181798 -16534 181833 -16500
rect 181992 -16577 182027 -16543
rect 182037 -16577 182038 -16532
rect 182137 -16543 182138 -16532
rect 182346 -16537 182381 -16503
rect 182391 -16537 182392 -16492
rect 182491 -16503 182492 -16492
rect 182736 -16496 182771 -16462
rect 182781 -16496 182782 -16451
rect 182881 -16462 182882 -16451
rect 182892 -16496 182927 -16462
rect 182937 -16496 182938 -16451
rect 183037 -16462 183038 -16451
rect 183218 -16456 183253 -16422
rect 183290 -16456 183325 -16422
rect 183362 -16456 183397 -16422
rect 183506 -16456 183541 -16422
rect 183578 -16456 183613 -16422
rect 183615 -16456 183685 -16422
rect 183722 -16456 183757 -16422
rect 183792 -16456 183827 -16422
rect 183048 -16496 183083 -16462
rect 184088 -16491 184123 -16457
rect 184133 -16491 184134 -16446
rect 184233 -16457 184234 -16446
rect 184244 -16491 184279 -16457
rect 184289 -16491 184290 -16446
rect 184389 -16457 184390 -16446
rect 184965 -16451 185000 -16417
rect 185142 -16451 185177 -16417
rect 184400 -16491 184435 -16457
rect 182502 -16537 182537 -16503
rect 183781 -16505 183782 -16494
rect 182148 -16577 182183 -16543
rect 181061 -16621 181096 -16587
rect 181262 -16666 181297 -16632
rect 181385 -16637 181386 -16595
rect 181707 -16624 181742 -16590
rect 182346 -16620 182381 -16586
rect 182391 -16620 182392 -16575
rect 182491 -16586 182492 -16575
rect 182736 -16580 182771 -16546
rect 182781 -16580 182782 -16535
rect 182881 -16546 182882 -16535
rect 182892 -16580 182927 -16546
rect 182937 -16580 182938 -16535
rect 183037 -16546 183038 -16535
rect 183615 -16539 183650 -16505
rect 183792 -16539 183827 -16505
rect 183048 -16580 183083 -16546
rect 183935 -16565 184050 -16499
rect 184233 -16525 184234 -16499
rect 184630 -16517 184665 -16483
rect 184675 -16517 184676 -16472
rect 184775 -16483 184776 -16472
rect 184786 -16517 184821 -16483
rect 184831 -16517 184832 -16472
rect 185131 -16500 185132 -16489
rect 185336 -16494 185371 -16460
rect 185381 -16494 185382 -16449
rect 185481 -16460 185482 -16449
rect 185690 -16453 185725 -16419
rect 185735 -16453 185736 -16408
rect 185835 -16419 185836 -16408
rect 186016 -16413 186051 -16379
rect 186080 -16413 186123 -16379
rect 186125 -16413 186126 -16371
rect 186225 -16379 186226 -16371
rect 186160 -16413 186195 -16379
rect 186236 -16413 186271 -16379
rect 186281 -16413 186282 -16371
rect 186381 -16379 186382 -16371
rect 186330 -16413 186365 -16379
rect 186392 -16413 186437 -16379
rect 187432 -16408 187467 -16374
rect 187477 -16408 187478 -16363
rect 187577 -16374 187578 -16363
rect 187588 -16408 187623 -16374
rect 187633 -16408 187634 -16363
rect 187733 -16374 187734 -16363
rect 188309 -16367 188344 -16333
rect 188486 -16367 188521 -16333
rect 189079 -16336 189080 -16328
rect 189179 -16336 189180 -16328
rect 187744 -16408 187779 -16374
rect 185846 -16453 185881 -16419
rect 187125 -16422 187126 -16414
rect 188475 -16417 188476 -16406
rect 188680 -16410 188715 -16376
rect 188725 -16410 188726 -16365
rect 188825 -16376 188826 -16365
rect 189006 -16370 189069 -16336
rect 189078 -16370 189113 -16336
rect 189190 -16370 189225 -16336
rect 189915 -16360 189950 -16326
rect 190011 -16360 190046 -16326
rect 190107 -16360 190142 -16326
rect 190203 -16360 190238 -16326
rect 190299 -16360 190334 -16326
rect 190395 -16360 190430 -16326
rect 190491 -16360 190526 -16326
rect 191819 -16333 191820 -16322
rect 191996 -16327 192059 -16293
rect 192068 -16327 192103 -16293
rect 192180 -16327 192215 -16293
rect 192711 -16317 192746 -16283
rect 192807 -16317 192842 -16283
rect 192903 -16317 192938 -16283
rect 192999 -16317 193034 -16283
rect 193095 -16317 193130 -16283
rect 194120 -16324 194155 -16290
rect 194165 -16324 194166 -16279
rect 194265 -16290 194266 -16279
rect 194276 -16324 194311 -16290
rect 194321 -16324 194322 -16279
rect 194421 -16290 194422 -16279
rect 194600 -16284 194635 -16250
rect 194672 -16284 194707 -16250
rect 194744 -16284 194779 -16250
rect 194888 -16284 194923 -16250
rect 194960 -16284 194995 -16250
rect 194997 -16284 195067 -16250
rect 195104 -16284 195139 -16250
rect 195174 -16284 195209 -16250
rect 195701 -16274 195736 -16240
rect 195797 -16274 195832 -16240
rect 195893 -16274 195928 -16240
rect 197400 -16241 197435 -16207
rect 197464 -16241 197507 -16207
rect 197509 -16241 197510 -16199
rect 197609 -16207 197610 -16199
rect 197544 -16241 197579 -16207
rect 197620 -16241 197655 -16207
rect 197665 -16241 197666 -16199
rect 197765 -16207 197766 -16199
rect 197714 -16241 197749 -16207
rect 197776 -16241 197821 -16207
rect 198691 -16231 198726 -16197
rect 198787 -16231 198822 -16197
rect 198883 -16231 198918 -16197
rect 198507 -16250 198508 -16242
rect 194432 -16324 194467 -16290
rect 195413 -16293 195414 -16285
rect 195513 -16293 195514 -16285
rect 188836 -16410 188871 -16376
rect 185492 -16494 185527 -16460
rect 182502 -16620 182537 -16586
rect 183781 -16589 183782 -16578
rect 181031 -16689 181032 -16681
rect 181042 -16723 181077 -16689
rect 181262 -16734 181297 -16700
rect 179709 -16793 179744 -16759
rect 179912 -16838 179947 -16804
rect 180035 -16809 180036 -16767
rect 180357 -16796 180392 -16762
rect 179679 -16861 179680 -16853
rect 179690 -16895 179725 -16861
rect 179912 -16906 179947 -16872
rect 179679 -16961 179680 -16950
rect 179690 -16995 179725 -16961
rect 178627 -17045 178662 -17011
rect 178723 -17045 178758 -17011
rect 178819 -17045 178854 -17011
rect 179328 -17035 179363 -17001
rect 179400 -17035 179435 -17001
rect 179472 -17035 179507 -17001
rect 179544 -17029 179580 -17001
rect 179890 -17025 179925 -16991
rect 179935 -17025 179936 -16980
rect 179544 -17035 179579 -17029
rect 178981 -17088 179016 -17054
rect 179077 -17088 179112 -17054
rect 179173 -17088 179208 -17054
rect 180077 -17076 180078 -16809
rect 180706 -16819 181093 -16753
rect 180093 -16860 180128 -16826
rect 180442 -16832 180453 -16819
rect 180376 -16874 180453 -16832
rect 180504 -16874 181093 -16819
rect 181240 -16853 181275 -16819
rect 181285 -16853 181286 -16808
rect 180376 -16877 181093 -16874
rect 180093 -16928 180128 -16894
rect 180296 -16942 180331 -16908
rect 180341 -16942 180342 -16900
rect 180177 -16991 180178 -16980
rect 180188 -17025 180223 -16991
rect 180296 -17042 180331 -17008
rect 180341 -17042 180342 -16997
rect 180189 -17078 180224 -17044
rect 180261 -17078 180296 -17044
rect 180333 -17078 180368 -17044
rect 179335 -17131 179370 -17097
rect 179431 -17131 179466 -17097
rect 179527 -17131 179562 -17097
rect 179623 -17131 179658 -17097
rect 179719 -17131 179754 -17097
rect 180376 -17114 180521 -16877
rect 180706 -16899 181093 -16877
rect 180630 -16925 181093 -16899
rect 181427 -16904 181428 -16637
rect 181443 -16688 181478 -16654
rect 182057 -16691 182092 -16657
rect 182736 -16663 182771 -16629
rect 182781 -16663 182782 -16618
rect 182881 -16629 182882 -16618
rect 182892 -16663 182927 -16629
rect 182937 -16663 182938 -16618
rect 183037 -16629 183038 -16618
rect 183615 -16623 183650 -16589
rect 183792 -16623 183827 -16589
rect 184153 -16605 184188 -16571
rect 183048 -16663 183083 -16629
rect 182881 -16697 182882 -16671
rect 183280 -16689 183315 -16655
rect 183325 -16689 183326 -16644
rect 183425 -16655 183426 -16644
rect 183436 -16689 183471 -16655
rect 183481 -16689 183482 -16644
rect 183781 -16672 183782 -16661
rect 181443 -16756 181478 -16722
rect 181646 -16770 181681 -16736
rect 181691 -16770 181692 -16728
rect 181791 -16740 181792 -16729
rect 182411 -16734 182446 -16700
rect 181802 -16774 181837 -16740
rect 181527 -16819 181528 -16808
rect 181996 -16813 182031 -16779
rect 182041 -16813 182042 -16771
rect 182141 -16779 182142 -16771
rect 182801 -16777 182836 -16743
rect 182152 -16813 182187 -16779
rect 181538 -16853 181573 -16819
rect 181646 -16870 181681 -16836
rect 181691 -16870 181692 -16825
rect 181791 -16832 181792 -16821
rect 181802 -16866 181837 -16832
rect 182350 -16856 182385 -16822
rect 182395 -16856 182396 -16814
rect 182495 -16822 182496 -16814
rect 182506 -16856 182541 -16822
rect 181539 -16906 181574 -16872
rect 181611 -16906 181646 -16872
rect 181683 -16906 181718 -16872
rect 181996 -16913 182031 -16879
rect 182041 -16913 182042 -16868
rect 182141 -16879 182142 -16868
rect 182152 -16913 182187 -16879
rect 182736 -16895 182771 -16861
rect 182781 -16895 182782 -16853
rect 180630 -16959 181106 -16925
rect 181964 -16949 181999 -16915
rect 182036 -16949 182071 -16915
rect 182350 -16956 182385 -16922
rect 182395 -16956 182396 -16911
rect 182495 -16922 182496 -16911
rect 182506 -16956 182541 -16922
rect 180630 -16985 181093 -16959
rect 180634 -16993 180835 -16985
rect 180650 -17003 180819 -16993
rect 180376 -17140 180551 -17114
rect 179883 -17174 179918 -17140
rect 179979 -17174 180014 -17140
rect 180075 -17174 180110 -17140
rect 180171 -17174 180206 -17140
rect 180267 -17174 180302 -17140
rect 180363 -17174 180551 -17140
rect 180376 -17200 180551 -17174
rect 180576 -17174 180677 -17050
rect 180454 -17870 180489 -17200
rect 180576 -17228 180579 -17174
rect 180261 -17936 180406 -17924
rect 179929 -17970 180406 -17936
rect 180261 -17971 180406 -17970
rect 180442 -17971 180489 -17870
rect 180588 -17971 180623 -17174
rect 180846 -17971 180881 -17062
rect 180980 -17971 181015 -16985
rect 181233 -17002 181268 -16968
rect 181329 -17002 181364 -16968
rect 181425 -17002 181460 -16968
rect 181521 -17002 181556 -16968
rect 181617 -17002 181652 -16968
rect 181713 -17002 181748 -16968
rect 181809 -17002 181844 -16968
rect 182318 -16992 182353 -16958
rect 182390 -16992 182425 -16958
rect 182736 -16995 182771 -16961
rect 182781 -16995 182782 -16950
rect 182923 -17001 182924 -16697
rect 183615 -16706 183650 -16672
rect 183792 -16706 183827 -16672
rect 184088 -16723 184123 -16689
rect 184133 -16723 184134 -16681
rect 184275 -16753 184276 -16525
rect 184965 -16534 185000 -16500
rect 185142 -16534 185177 -16500
rect 185336 -16577 185371 -16543
rect 185381 -16577 185382 -16532
rect 185481 -16543 185482 -16532
rect 185690 -16537 185725 -16503
rect 185735 -16537 185736 -16492
rect 185835 -16503 185836 -16492
rect 186080 -16496 186115 -16462
rect 186125 -16496 186126 -16451
rect 186225 -16462 186226 -16451
rect 186236 -16496 186271 -16462
rect 186281 -16496 186282 -16451
rect 186381 -16462 186382 -16451
rect 186562 -16456 186597 -16422
rect 186634 -16456 186669 -16422
rect 186706 -16456 186741 -16422
rect 186850 -16456 186885 -16422
rect 186922 -16456 186957 -16422
rect 186959 -16456 187029 -16422
rect 187066 -16456 187101 -16422
rect 187136 -16456 187171 -16422
rect 186392 -16496 186427 -16462
rect 187432 -16491 187467 -16457
rect 187477 -16491 187478 -16446
rect 187577 -16457 187578 -16446
rect 187588 -16491 187623 -16457
rect 187633 -16491 187634 -16446
rect 187733 -16457 187734 -16446
rect 188309 -16451 188344 -16417
rect 188486 -16451 188521 -16417
rect 187744 -16491 187779 -16457
rect 185846 -16537 185881 -16503
rect 187125 -16505 187126 -16494
rect 185492 -16577 185527 -16543
rect 184405 -16621 184440 -16587
rect 184606 -16666 184641 -16632
rect 184729 -16637 184730 -16595
rect 185051 -16624 185086 -16590
rect 185690 -16620 185725 -16586
rect 185735 -16620 185736 -16575
rect 185835 -16586 185836 -16575
rect 186080 -16580 186115 -16546
rect 186125 -16580 186126 -16535
rect 186225 -16546 186226 -16535
rect 186236 -16580 186271 -16546
rect 186281 -16580 186282 -16535
rect 186381 -16546 186382 -16535
rect 186959 -16539 186994 -16505
rect 187136 -16539 187171 -16505
rect 186392 -16580 186427 -16546
rect 187279 -16565 187394 -16499
rect 187577 -16525 187578 -16499
rect 187974 -16517 188009 -16483
rect 188019 -16517 188020 -16472
rect 188119 -16483 188120 -16472
rect 188130 -16517 188165 -16483
rect 188175 -16517 188176 -16472
rect 188475 -16500 188476 -16489
rect 188680 -16494 188715 -16460
rect 188725 -16494 188726 -16449
rect 188825 -16460 188826 -16449
rect 189034 -16453 189069 -16419
rect 189079 -16453 189080 -16408
rect 189179 -16419 189180 -16408
rect 189360 -16413 189395 -16379
rect 189424 -16413 189467 -16379
rect 189469 -16413 189470 -16371
rect 189569 -16379 189570 -16371
rect 189504 -16413 189539 -16379
rect 189580 -16413 189615 -16379
rect 189625 -16413 189626 -16371
rect 189725 -16379 189726 -16371
rect 189674 -16413 189709 -16379
rect 189736 -16413 189781 -16379
rect 190776 -16408 190811 -16374
rect 190821 -16408 190822 -16363
rect 190921 -16374 190922 -16363
rect 190932 -16408 190967 -16374
rect 190977 -16408 190978 -16363
rect 191077 -16374 191078 -16363
rect 191653 -16367 191688 -16333
rect 191830 -16367 191865 -16333
rect 192423 -16336 192424 -16328
rect 192523 -16336 192524 -16328
rect 191088 -16408 191123 -16374
rect 189190 -16453 189225 -16419
rect 190469 -16422 190470 -16414
rect 191819 -16417 191820 -16406
rect 192024 -16410 192059 -16376
rect 192069 -16410 192070 -16365
rect 192169 -16376 192170 -16365
rect 192350 -16370 192413 -16336
rect 192422 -16370 192457 -16336
rect 192534 -16370 192569 -16336
rect 193259 -16360 193294 -16326
rect 193355 -16360 193390 -16326
rect 193451 -16360 193486 -16326
rect 193547 -16360 193582 -16326
rect 193643 -16360 193678 -16326
rect 193739 -16360 193774 -16326
rect 193835 -16360 193870 -16326
rect 195163 -16333 195164 -16322
rect 195340 -16327 195403 -16293
rect 195412 -16327 195447 -16293
rect 195524 -16327 195559 -16293
rect 196055 -16317 196090 -16283
rect 196151 -16317 196186 -16283
rect 196247 -16317 196282 -16283
rect 196343 -16317 196378 -16283
rect 196439 -16317 196474 -16283
rect 197464 -16324 197499 -16290
rect 197509 -16324 197510 -16279
rect 197609 -16290 197610 -16279
rect 197620 -16324 197655 -16290
rect 197665 -16324 197666 -16279
rect 197765 -16290 197766 -16279
rect 197944 -16284 197979 -16250
rect 198016 -16284 198051 -16250
rect 198088 -16284 198123 -16250
rect 198232 -16284 198267 -16250
rect 198304 -16284 198339 -16250
rect 198341 -16284 198411 -16250
rect 198448 -16284 198483 -16250
rect 198518 -16284 198553 -16250
rect 199045 -16274 199080 -16240
rect 199141 -16274 199176 -16240
rect 199237 -16274 199272 -16240
rect 200744 -16241 200779 -16207
rect 200808 -16241 200851 -16207
rect 200853 -16241 200854 -16199
rect 200953 -16207 200954 -16199
rect 200888 -16241 200923 -16207
rect 200964 -16241 200999 -16207
rect 201009 -16241 201010 -16199
rect 201109 -16207 201110 -16199
rect 201058 -16241 201093 -16207
rect 201120 -16241 201165 -16207
rect 202035 -16231 202070 -16197
rect 202131 -16231 202166 -16197
rect 202227 -16231 202262 -16197
rect 201851 -16250 201852 -16242
rect 197776 -16324 197811 -16290
rect 198757 -16293 198758 -16285
rect 198857 -16293 198858 -16285
rect 192180 -16410 192215 -16376
rect 188836 -16494 188871 -16460
rect 185846 -16620 185881 -16586
rect 187125 -16589 187126 -16578
rect 184375 -16689 184376 -16681
rect 184386 -16723 184421 -16689
rect 184606 -16734 184641 -16700
rect 183053 -16793 183088 -16759
rect 183256 -16838 183291 -16804
rect 183379 -16809 183380 -16767
rect 183701 -16796 183736 -16762
rect 183023 -16861 183024 -16853
rect 183034 -16895 183069 -16861
rect 183256 -16906 183291 -16872
rect 183023 -16961 183024 -16950
rect 183034 -16995 183069 -16961
rect 181971 -17045 182006 -17011
rect 182067 -17045 182102 -17011
rect 182163 -17045 182198 -17011
rect 182672 -17035 182707 -17001
rect 182744 -17035 182779 -17001
rect 182816 -17035 182851 -17001
rect 182888 -17029 182924 -17001
rect 183234 -17025 183269 -16991
rect 183279 -17025 183280 -16980
rect 182888 -17035 182923 -17029
rect 182325 -17088 182360 -17054
rect 182421 -17088 182456 -17054
rect 182517 -17088 182552 -17054
rect 183421 -17076 183422 -16809
rect 184050 -16819 184437 -16753
rect 183437 -16860 183472 -16826
rect 183786 -16832 183797 -16819
rect 183720 -16874 183797 -16832
rect 183848 -16874 184437 -16819
rect 184584 -16853 184619 -16819
rect 184629 -16853 184630 -16808
rect 183720 -16877 184437 -16874
rect 183437 -16928 183472 -16894
rect 183640 -16942 183675 -16908
rect 183685 -16942 183686 -16900
rect 183521 -16991 183522 -16980
rect 183532 -17025 183567 -16991
rect 183640 -17042 183675 -17008
rect 183685 -17042 183686 -16997
rect 183533 -17078 183568 -17044
rect 183605 -17078 183640 -17044
rect 183677 -17078 183712 -17044
rect 182679 -17131 182714 -17097
rect 182775 -17131 182810 -17097
rect 182871 -17131 182906 -17097
rect 182967 -17131 183002 -17097
rect 183063 -17131 183098 -17097
rect 183720 -17114 183865 -16877
rect 184050 -16899 184437 -16877
rect 183974 -16925 184437 -16899
rect 184771 -16904 184772 -16637
rect 184787 -16688 184822 -16654
rect 185401 -16691 185436 -16657
rect 186080 -16663 186115 -16629
rect 186125 -16663 186126 -16618
rect 186225 -16629 186226 -16618
rect 186236 -16663 186271 -16629
rect 186281 -16663 186282 -16618
rect 186381 -16629 186382 -16618
rect 186959 -16623 186994 -16589
rect 187136 -16623 187171 -16589
rect 187497 -16605 187532 -16571
rect 186392 -16663 186427 -16629
rect 186225 -16697 186226 -16671
rect 186624 -16689 186659 -16655
rect 186669 -16689 186670 -16644
rect 186769 -16655 186770 -16644
rect 186780 -16689 186815 -16655
rect 186825 -16689 186826 -16644
rect 187125 -16672 187126 -16661
rect 184787 -16756 184822 -16722
rect 184990 -16770 185025 -16736
rect 185035 -16770 185036 -16728
rect 185135 -16740 185136 -16729
rect 185755 -16734 185790 -16700
rect 185146 -16774 185181 -16740
rect 184871 -16819 184872 -16808
rect 185340 -16813 185375 -16779
rect 185385 -16813 185386 -16771
rect 185485 -16779 185486 -16771
rect 186145 -16777 186180 -16743
rect 185496 -16813 185531 -16779
rect 184882 -16853 184917 -16819
rect 184990 -16870 185025 -16836
rect 185035 -16870 185036 -16825
rect 185135 -16832 185136 -16821
rect 185146 -16866 185181 -16832
rect 185694 -16856 185729 -16822
rect 185739 -16856 185740 -16814
rect 185839 -16822 185840 -16814
rect 185850 -16856 185885 -16822
rect 184883 -16906 184918 -16872
rect 184955 -16906 184990 -16872
rect 185027 -16906 185062 -16872
rect 185340 -16913 185375 -16879
rect 185385 -16913 185386 -16868
rect 185485 -16879 185486 -16868
rect 185496 -16913 185531 -16879
rect 186080 -16895 186115 -16861
rect 186125 -16895 186126 -16853
rect 183974 -16959 184450 -16925
rect 185308 -16949 185343 -16915
rect 185380 -16949 185415 -16915
rect 185694 -16956 185729 -16922
rect 185739 -16956 185740 -16911
rect 185839 -16922 185840 -16911
rect 185850 -16956 185885 -16922
rect 183974 -16985 184437 -16959
rect 183978 -16993 184179 -16985
rect 183994 -17003 184163 -16993
rect 183720 -17140 183895 -17114
rect 183227 -17174 183262 -17140
rect 183323 -17174 183358 -17140
rect 183419 -17174 183454 -17140
rect 183515 -17174 183550 -17140
rect 183611 -17174 183646 -17140
rect 183707 -17174 183895 -17140
rect 183720 -17200 183895 -17174
rect 183920 -17174 184021 -17050
rect 183798 -17870 183833 -17200
rect 183920 -17228 183923 -17174
rect 183605 -17936 183750 -17924
rect 183273 -17970 183750 -17936
rect 183605 -17971 183750 -17970
rect 183786 -17971 183833 -17870
rect 183932 -17971 183967 -17174
rect 184190 -17971 184225 -17062
rect 184324 -17971 184359 -16985
rect 184577 -17002 184612 -16968
rect 184673 -17002 184708 -16968
rect 184769 -17002 184804 -16968
rect 184865 -17002 184900 -16968
rect 184961 -17002 184996 -16968
rect 185057 -17002 185092 -16968
rect 185153 -17002 185188 -16968
rect 185662 -16992 185697 -16958
rect 185734 -16992 185769 -16958
rect 186080 -16995 186115 -16961
rect 186125 -16995 186126 -16950
rect 186267 -17001 186268 -16697
rect 186959 -16706 186994 -16672
rect 187136 -16706 187171 -16672
rect 187432 -16723 187467 -16689
rect 187477 -16723 187478 -16681
rect 187619 -16753 187620 -16525
rect 188309 -16534 188344 -16500
rect 188486 -16534 188521 -16500
rect 188680 -16577 188715 -16543
rect 188725 -16577 188726 -16532
rect 188825 -16543 188826 -16532
rect 189034 -16537 189069 -16503
rect 189079 -16537 189080 -16492
rect 189179 -16503 189180 -16492
rect 189424 -16496 189459 -16462
rect 189469 -16496 189470 -16451
rect 189569 -16462 189570 -16451
rect 189580 -16496 189615 -16462
rect 189625 -16496 189626 -16451
rect 189725 -16462 189726 -16451
rect 189906 -16456 189941 -16422
rect 189978 -16456 190013 -16422
rect 190050 -16456 190085 -16422
rect 190194 -16456 190229 -16422
rect 190266 -16456 190301 -16422
rect 190303 -16456 190373 -16422
rect 190410 -16456 190445 -16422
rect 190480 -16456 190515 -16422
rect 189736 -16496 189771 -16462
rect 190776 -16491 190811 -16457
rect 190821 -16491 190822 -16446
rect 190921 -16457 190922 -16446
rect 190932 -16491 190967 -16457
rect 190977 -16491 190978 -16446
rect 191077 -16457 191078 -16446
rect 191653 -16451 191688 -16417
rect 191830 -16451 191865 -16417
rect 191088 -16491 191123 -16457
rect 189190 -16537 189225 -16503
rect 190469 -16505 190470 -16494
rect 188836 -16577 188871 -16543
rect 187749 -16621 187784 -16587
rect 187950 -16666 187985 -16632
rect 188073 -16637 188074 -16595
rect 188395 -16624 188430 -16590
rect 189034 -16620 189069 -16586
rect 189079 -16620 189080 -16575
rect 189179 -16586 189180 -16575
rect 189424 -16580 189459 -16546
rect 189469 -16580 189470 -16535
rect 189569 -16546 189570 -16535
rect 189580 -16580 189615 -16546
rect 189625 -16580 189626 -16535
rect 189725 -16546 189726 -16535
rect 190303 -16539 190338 -16505
rect 190480 -16539 190515 -16505
rect 189736 -16580 189771 -16546
rect 190623 -16565 190738 -16499
rect 190921 -16525 190922 -16499
rect 191318 -16517 191353 -16483
rect 191363 -16517 191364 -16472
rect 191463 -16483 191464 -16472
rect 191474 -16517 191509 -16483
rect 191519 -16517 191520 -16472
rect 191819 -16500 191820 -16489
rect 192024 -16494 192059 -16460
rect 192069 -16494 192070 -16449
rect 192169 -16460 192170 -16449
rect 192378 -16453 192413 -16419
rect 192423 -16453 192424 -16408
rect 192523 -16419 192524 -16408
rect 192704 -16413 192739 -16379
rect 192768 -16413 192811 -16379
rect 192813 -16413 192814 -16371
rect 192913 -16379 192914 -16371
rect 192848 -16413 192883 -16379
rect 192924 -16413 192959 -16379
rect 192969 -16413 192970 -16371
rect 193069 -16379 193070 -16371
rect 193018 -16413 193053 -16379
rect 193080 -16413 193125 -16379
rect 194120 -16408 194155 -16374
rect 194165 -16408 194166 -16363
rect 194265 -16374 194266 -16363
rect 194276 -16408 194311 -16374
rect 194321 -16408 194322 -16363
rect 194421 -16374 194422 -16363
rect 194997 -16367 195032 -16333
rect 195174 -16367 195209 -16333
rect 195767 -16336 195768 -16328
rect 195867 -16336 195868 -16328
rect 194432 -16408 194467 -16374
rect 192534 -16453 192569 -16419
rect 193813 -16422 193814 -16414
rect 195163 -16417 195164 -16406
rect 195368 -16410 195403 -16376
rect 195413 -16410 195414 -16365
rect 195513 -16376 195514 -16365
rect 195694 -16370 195757 -16336
rect 195766 -16370 195801 -16336
rect 195878 -16370 195913 -16336
rect 196603 -16360 196638 -16326
rect 196699 -16360 196734 -16326
rect 196795 -16360 196830 -16326
rect 196891 -16360 196926 -16326
rect 196987 -16360 197022 -16326
rect 197083 -16360 197118 -16326
rect 197179 -16360 197214 -16326
rect 198507 -16333 198508 -16322
rect 198684 -16327 198747 -16293
rect 198756 -16327 198791 -16293
rect 198868 -16327 198903 -16293
rect 199399 -16317 199434 -16283
rect 199495 -16317 199530 -16283
rect 199591 -16317 199626 -16283
rect 199687 -16317 199722 -16283
rect 199783 -16317 199818 -16283
rect 200808 -16324 200843 -16290
rect 200853 -16324 200854 -16279
rect 200953 -16290 200954 -16279
rect 200964 -16324 200999 -16290
rect 201009 -16324 201010 -16279
rect 201109 -16290 201110 -16279
rect 201288 -16284 201323 -16250
rect 201360 -16284 201395 -16250
rect 201432 -16284 201467 -16250
rect 201576 -16284 201611 -16250
rect 201648 -16284 201683 -16250
rect 201685 -16284 201755 -16250
rect 201792 -16284 201827 -16250
rect 201862 -16284 201897 -16250
rect 202389 -16274 202424 -16240
rect 202485 -16274 202520 -16240
rect 202581 -16274 202616 -16240
rect 204088 -16241 204123 -16207
rect 204152 -16241 204195 -16207
rect 204197 -16241 204198 -16199
rect 204297 -16207 204298 -16199
rect 204232 -16241 204267 -16207
rect 204308 -16241 204343 -16207
rect 204353 -16241 204354 -16199
rect 204453 -16207 204454 -16199
rect 204402 -16241 204437 -16207
rect 204464 -16241 204509 -16207
rect 205379 -16231 205414 -16197
rect 205475 -16231 205510 -16197
rect 205571 -16231 205606 -16197
rect 205195 -16250 205196 -16242
rect 201120 -16324 201155 -16290
rect 202101 -16293 202102 -16285
rect 202201 -16293 202202 -16285
rect 195524 -16410 195559 -16376
rect 192180 -16494 192215 -16460
rect 189190 -16620 189225 -16586
rect 190469 -16589 190470 -16578
rect 187719 -16689 187720 -16681
rect 187730 -16723 187765 -16689
rect 187950 -16734 187985 -16700
rect 186397 -16793 186432 -16759
rect 186600 -16838 186635 -16804
rect 186723 -16809 186724 -16767
rect 187045 -16796 187080 -16762
rect 186367 -16861 186368 -16853
rect 186378 -16895 186413 -16861
rect 186600 -16906 186635 -16872
rect 186367 -16961 186368 -16950
rect 186378 -16995 186413 -16961
rect 185315 -17045 185350 -17011
rect 185411 -17045 185446 -17011
rect 185507 -17045 185542 -17011
rect 186016 -17035 186051 -17001
rect 186088 -17035 186123 -17001
rect 186160 -17035 186195 -17001
rect 186232 -17029 186268 -17001
rect 186578 -17025 186613 -16991
rect 186623 -17025 186624 -16980
rect 186232 -17035 186267 -17029
rect 185669 -17088 185704 -17054
rect 185765 -17088 185800 -17054
rect 185861 -17088 185896 -17054
rect 186765 -17076 186766 -16809
rect 187394 -16819 187781 -16753
rect 186781 -16860 186816 -16826
rect 187130 -16832 187141 -16819
rect 187064 -16874 187141 -16832
rect 187192 -16874 187781 -16819
rect 187928 -16853 187963 -16819
rect 187973 -16853 187974 -16808
rect 187064 -16877 187781 -16874
rect 186781 -16928 186816 -16894
rect 186984 -16942 187019 -16908
rect 187029 -16942 187030 -16900
rect 186865 -16991 186866 -16980
rect 186876 -17025 186911 -16991
rect 186984 -17042 187019 -17008
rect 187029 -17042 187030 -16997
rect 186877 -17078 186912 -17044
rect 186949 -17078 186984 -17044
rect 187021 -17078 187056 -17044
rect 186023 -17131 186058 -17097
rect 186119 -17131 186154 -17097
rect 186215 -17131 186250 -17097
rect 186311 -17131 186346 -17097
rect 186407 -17131 186442 -17097
rect 187064 -17114 187209 -16877
rect 187394 -16899 187781 -16877
rect 187318 -16925 187781 -16899
rect 188115 -16904 188116 -16637
rect 188131 -16688 188166 -16654
rect 188745 -16691 188780 -16657
rect 189424 -16663 189459 -16629
rect 189469 -16663 189470 -16618
rect 189569 -16629 189570 -16618
rect 189580 -16663 189615 -16629
rect 189625 -16663 189626 -16618
rect 189725 -16629 189726 -16618
rect 190303 -16623 190338 -16589
rect 190480 -16623 190515 -16589
rect 190841 -16605 190876 -16571
rect 189736 -16663 189771 -16629
rect 189569 -16697 189570 -16671
rect 189968 -16689 190003 -16655
rect 190013 -16689 190014 -16644
rect 190113 -16655 190114 -16644
rect 190124 -16689 190159 -16655
rect 190169 -16689 190170 -16644
rect 190469 -16672 190470 -16661
rect 188131 -16756 188166 -16722
rect 188334 -16770 188369 -16736
rect 188379 -16770 188380 -16728
rect 188479 -16740 188480 -16729
rect 189099 -16734 189134 -16700
rect 188490 -16774 188525 -16740
rect 188215 -16819 188216 -16808
rect 188684 -16813 188719 -16779
rect 188729 -16813 188730 -16771
rect 188829 -16779 188830 -16771
rect 189489 -16777 189524 -16743
rect 188840 -16813 188875 -16779
rect 188226 -16853 188261 -16819
rect 188334 -16870 188369 -16836
rect 188379 -16870 188380 -16825
rect 188479 -16832 188480 -16821
rect 188490 -16866 188525 -16832
rect 189038 -16856 189073 -16822
rect 189083 -16856 189084 -16814
rect 189183 -16822 189184 -16814
rect 189194 -16856 189229 -16822
rect 188227 -16906 188262 -16872
rect 188299 -16906 188334 -16872
rect 188371 -16906 188406 -16872
rect 188684 -16913 188719 -16879
rect 188729 -16913 188730 -16868
rect 188829 -16879 188830 -16868
rect 188840 -16913 188875 -16879
rect 189424 -16895 189459 -16861
rect 189469 -16895 189470 -16853
rect 187318 -16959 187794 -16925
rect 188652 -16949 188687 -16915
rect 188724 -16949 188759 -16915
rect 189038 -16956 189073 -16922
rect 189083 -16956 189084 -16911
rect 189183 -16922 189184 -16911
rect 189194 -16956 189229 -16922
rect 187318 -16985 187781 -16959
rect 187322 -16993 187523 -16985
rect 187338 -17003 187507 -16993
rect 187064 -17140 187239 -17114
rect 186571 -17174 186606 -17140
rect 186667 -17174 186702 -17140
rect 186763 -17174 186798 -17140
rect 186859 -17174 186894 -17140
rect 186955 -17174 186990 -17140
rect 187051 -17174 187239 -17140
rect 187064 -17200 187239 -17174
rect 187264 -17174 187365 -17050
rect 187142 -17870 187177 -17200
rect 187264 -17228 187267 -17174
rect 186949 -17936 187094 -17924
rect 186617 -17970 187094 -17936
rect 186949 -17971 187094 -17970
rect 187130 -17971 187177 -17870
rect 187276 -17971 187311 -17174
rect 187534 -17971 187569 -17062
rect 187668 -17971 187703 -16985
rect 187921 -17002 187956 -16968
rect 188017 -17002 188052 -16968
rect 188113 -17002 188148 -16968
rect 188209 -17002 188244 -16968
rect 188305 -17002 188340 -16968
rect 188401 -17002 188436 -16968
rect 188497 -17002 188532 -16968
rect 189006 -16992 189041 -16958
rect 189078 -16992 189113 -16958
rect 189424 -16995 189459 -16961
rect 189469 -16995 189470 -16950
rect 189611 -17001 189612 -16697
rect 190303 -16706 190338 -16672
rect 190480 -16706 190515 -16672
rect 190776 -16723 190811 -16689
rect 190821 -16723 190822 -16681
rect 190963 -16753 190964 -16525
rect 191653 -16534 191688 -16500
rect 191830 -16534 191865 -16500
rect 192024 -16577 192059 -16543
rect 192069 -16577 192070 -16532
rect 192169 -16543 192170 -16532
rect 192378 -16537 192413 -16503
rect 192423 -16537 192424 -16492
rect 192523 -16503 192524 -16492
rect 192768 -16496 192803 -16462
rect 192813 -16496 192814 -16451
rect 192913 -16462 192914 -16451
rect 192924 -16496 192959 -16462
rect 192969 -16496 192970 -16451
rect 193069 -16462 193070 -16451
rect 193250 -16456 193285 -16422
rect 193322 -16456 193357 -16422
rect 193394 -16456 193429 -16422
rect 193538 -16456 193573 -16422
rect 193610 -16456 193645 -16422
rect 193647 -16456 193717 -16422
rect 193754 -16456 193789 -16422
rect 193824 -16456 193859 -16422
rect 193080 -16496 193115 -16462
rect 194120 -16491 194155 -16457
rect 194165 -16491 194166 -16446
rect 194265 -16457 194266 -16446
rect 194276 -16491 194311 -16457
rect 194321 -16491 194322 -16446
rect 194421 -16457 194422 -16446
rect 194997 -16451 195032 -16417
rect 195174 -16451 195209 -16417
rect 194432 -16491 194467 -16457
rect 192534 -16537 192569 -16503
rect 193813 -16505 193814 -16494
rect 192180 -16577 192215 -16543
rect 191093 -16621 191128 -16587
rect 191294 -16666 191329 -16632
rect 191417 -16637 191418 -16595
rect 191739 -16624 191774 -16590
rect 192378 -16620 192413 -16586
rect 192423 -16620 192424 -16575
rect 192523 -16586 192524 -16575
rect 192768 -16580 192803 -16546
rect 192813 -16580 192814 -16535
rect 192913 -16546 192914 -16535
rect 192924 -16580 192959 -16546
rect 192969 -16580 192970 -16535
rect 193069 -16546 193070 -16535
rect 193647 -16539 193682 -16505
rect 193824 -16539 193859 -16505
rect 193080 -16580 193115 -16546
rect 193967 -16565 194082 -16499
rect 194265 -16525 194266 -16499
rect 194662 -16517 194697 -16483
rect 194707 -16517 194708 -16472
rect 194807 -16483 194808 -16472
rect 194818 -16517 194853 -16483
rect 194863 -16517 194864 -16472
rect 195163 -16500 195164 -16489
rect 195368 -16494 195403 -16460
rect 195413 -16494 195414 -16449
rect 195513 -16460 195514 -16449
rect 195722 -16453 195757 -16419
rect 195767 -16453 195768 -16408
rect 195867 -16419 195868 -16408
rect 196048 -16413 196083 -16379
rect 196112 -16413 196155 -16379
rect 196157 -16413 196158 -16371
rect 196257 -16379 196258 -16371
rect 196192 -16413 196227 -16379
rect 196268 -16413 196303 -16379
rect 196313 -16413 196314 -16371
rect 196413 -16379 196414 -16371
rect 196362 -16413 196397 -16379
rect 196424 -16413 196469 -16379
rect 197464 -16408 197499 -16374
rect 197509 -16408 197510 -16363
rect 197609 -16374 197610 -16363
rect 197620 -16408 197655 -16374
rect 197665 -16408 197666 -16363
rect 197765 -16374 197766 -16363
rect 198341 -16367 198376 -16333
rect 198518 -16367 198553 -16333
rect 199111 -16336 199112 -16328
rect 199211 -16336 199212 -16328
rect 197776 -16408 197811 -16374
rect 195878 -16453 195913 -16419
rect 197157 -16422 197158 -16414
rect 198507 -16417 198508 -16406
rect 198712 -16410 198747 -16376
rect 198757 -16410 198758 -16365
rect 198857 -16376 198858 -16365
rect 199038 -16370 199101 -16336
rect 199110 -16370 199145 -16336
rect 199222 -16370 199257 -16336
rect 199947 -16360 199982 -16326
rect 200043 -16360 200078 -16326
rect 200139 -16360 200174 -16326
rect 200235 -16360 200270 -16326
rect 200331 -16360 200366 -16326
rect 200427 -16360 200462 -16326
rect 200523 -16360 200558 -16326
rect 201851 -16333 201852 -16322
rect 202028 -16327 202091 -16293
rect 202100 -16327 202135 -16293
rect 202212 -16327 202247 -16293
rect 202743 -16317 202778 -16283
rect 202839 -16317 202874 -16283
rect 202935 -16317 202970 -16283
rect 203031 -16317 203066 -16283
rect 203127 -16317 203162 -16283
rect 204152 -16324 204187 -16290
rect 204197 -16324 204198 -16279
rect 204297 -16290 204298 -16279
rect 204308 -16324 204343 -16290
rect 204353 -16324 204354 -16279
rect 204453 -16290 204454 -16279
rect 204632 -16284 204667 -16250
rect 204704 -16284 204739 -16250
rect 204776 -16284 204811 -16250
rect 204920 -16284 204955 -16250
rect 204992 -16284 205027 -16250
rect 205029 -16284 205099 -16250
rect 205136 -16284 205171 -16250
rect 205206 -16284 205241 -16250
rect 205733 -16274 205768 -16240
rect 205829 -16274 205864 -16240
rect 205925 -16274 205960 -16240
rect 207432 -16241 207467 -16207
rect 207496 -16241 207539 -16207
rect 207541 -16241 207542 -16199
rect 207641 -16207 207642 -16199
rect 207576 -16241 207611 -16207
rect 207652 -16241 207687 -16207
rect 207697 -16241 207698 -16199
rect 207797 -16207 207798 -16199
rect 207746 -16241 207781 -16207
rect 207808 -16241 207853 -16207
rect 208723 -16231 208758 -16197
rect 208819 -16231 208854 -16197
rect 208915 -16231 208950 -16197
rect 208539 -16250 208540 -16242
rect 204464 -16324 204499 -16290
rect 205445 -16293 205446 -16285
rect 205545 -16293 205546 -16285
rect 198868 -16410 198903 -16376
rect 195524 -16494 195559 -16460
rect 192534 -16620 192569 -16586
rect 193813 -16589 193814 -16578
rect 191063 -16689 191064 -16681
rect 191074 -16723 191109 -16689
rect 191294 -16734 191329 -16700
rect 189741 -16793 189776 -16759
rect 189944 -16838 189979 -16804
rect 190067 -16809 190068 -16767
rect 190389 -16796 190424 -16762
rect 189711 -16861 189712 -16853
rect 189722 -16895 189757 -16861
rect 189944 -16906 189979 -16872
rect 189711 -16961 189712 -16950
rect 189722 -16995 189757 -16961
rect 188659 -17045 188694 -17011
rect 188755 -17045 188790 -17011
rect 188851 -17045 188886 -17011
rect 189360 -17035 189395 -17001
rect 189432 -17035 189467 -17001
rect 189504 -17035 189539 -17001
rect 189576 -17029 189612 -17001
rect 189922 -17025 189957 -16991
rect 189967 -17025 189968 -16980
rect 189576 -17035 189611 -17029
rect 189013 -17088 189048 -17054
rect 189109 -17088 189144 -17054
rect 189205 -17088 189240 -17054
rect 190109 -17076 190110 -16809
rect 190738 -16819 191125 -16753
rect 190125 -16860 190160 -16826
rect 190474 -16832 190485 -16819
rect 190408 -16874 190485 -16832
rect 190536 -16874 191125 -16819
rect 191272 -16853 191307 -16819
rect 191317 -16853 191318 -16808
rect 190408 -16877 191125 -16874
rect 190125 -16928 190160 -16894
rect 190328 -16942 190363 -16908
rect 190373 -16942 190374 -16900
rect 190209 -16991 190210 -16980
rect 190220 -17025 190255 -16991
rect 190328 -17042 190363 -17008
rect 190373 -17042 190374 -16997
rect 190221 -17078 190256 -17044
rect 190293 -17078 190328 -17044
rect 190365 -17078 190400 -17044
rect 189367 -17131 189402 -17097
rect 189463 -17131 189498 -17097
rect 189559 -17131 189594 -17097
rect 189655 -17131 189690 -17097
rect 189751 -17131 189786 -17097
rect 190408 -17114 190553 -16877
rect 190738 -16899 191125 -16877
rect 190662 -16925 191125 -16899
rect 191459 -16904 191460 -16637
rect 191475 -16688 191510 -16654
rect 192089 -16691 192124 -16657
rect 192768 -16663 192803 -16629
rect 192813 -16663 192814 -16618
rect 192913 -16629 192914 -16618
rect 192924 -16663 192959 -16629
rect 192969 -16663 192970 -16618
rect 193069 -16629 193070 -16618
rect 193647 -16623 193682 -16589
rect 193824 -16623 193859 -16589
rect 194185 -16605 194220 -16571
rect 193080 -16663 193115 -16629
rect 192913 -16697 192914 -16671
rect 193312 -16689 193347 -16655
rect 193357 -16689 193358 -16644
rect 193457 -16655 193458 -16644
rect 193468 -16689 193503 -16655
rect 193513 -16689 193514 -16644
rect 193813 -16672 193814 -16661
rect 191475 -16756 191510 -16722
rect 191678 -16770 191713 -16736
rect 191723 -16770 191724 -16728
rect 191823 -16740 191824 -16729
rect 192443 -16734 192478 -16700
rect 191834 -16774 191869 -16740
rect 191559 -16819 191560 -16808
rect 192028 -16813 192063 -16779
rect 192073 -16813 192074 -16771
rect 192173 -16779 192174 -16771
rect 192833 -16777 192868 -16743
rect 192184 -16813 192219 -16779
rect 191570 -16853 191605 -16819
rect 191678 -16870 191713 -16836
rect 191723 -16870 191724 -16825
rect 191823 -16832 191824 -16821
rect 191834 -16866 191869 -16832
rect 192382 -16856 192417 -16822
rect 192427 -16856 192428 -16814
rect 192527 -16822 192528 -16814
rect 192538 -16856 192573 -16822
rect 191571 -16906 191606 -16872
rect 191643 -16906 191678 -16872
rect 191715 -16906 191750 -16872
rect 192028 -16913 192063 -16879
rect 192073 -16913 192074 -16868
rect 192173 -16879 192174 -16868
rect 192184 -16913 192219 -16879
rect 192768 -16895 192803 -16861
rect 192813 -16895 192814 -16853
rect 190662 -16959 191138 -16925
rect 191996 -16949 192031 -16915
rect 192068 -16949 192103 -16915
rect 192382 -16956 192417 -16922
rect 192427 -16956 192428 -16911
rect 192527 -16922 192528 -16911
rect 192538 -16956 192573 -16922
rect 190662 -16985 191125 -16959
rect 190666 -16993 190867 -16985
rect 190682 -17003 190851 -16993
rect 190408 -17140 190583 -17114
rect 189915 -17174 189950 -17140
rect 190011 -17174 190046 -17140
rect 190107 -17174 190142 -17140
rect 190203 -17174 190238 -17140
rect 190299 -17174 190334 -17140
rect 190395 -17174 190583 -17140
rect 190408 -17200 190583 -17174
rect 190608 -17174 190709 -17050
rect 190486 -17870 190521 -17200
rect 190608 -17228 190611 -17174
rect 190293 -17936 190438 -17924
rect 189961 -17970 190438 -17936
rect 190293 -17971 190438 -17970
rect 190474 -17971 190521 -17870
rect 190620 -17971 190655 -17174
rect 190878 -17971 190913 -17062
rect 191012 -17971 191047 -16985
rect 191265 -17002 191300 -16968
rect 191361 -17002 191396 -16968
rect 191457 -17002 191492 -16968
rect 191553 -17002 191588 -16968
rect 191649 -17002 191684 -16968
rect 191745 -17002 191780 -16968
rect 191841 -17002 191876 -16968
rect 192350 -16992 192385 -16958
rect 192422 -16992 192457 -16958
rect 192768 -16995 192803 -16961
rect 192813 -16995 192814 -16950
rect 192955 -17001 192956 -16697
rect 193647 -16706 193682 -16672
rect 193824 -16706 193859 -16672
rect 194120 -16723 194155 -16689
rect 194165 -16723 194166 -16681
rect 194307 -16753 194308 -16525
rect 194997 -16534 195032 -16500
rect 195174 -16534 195209 -16500
rect 195368 -16577 195403 -16543
rect 195413 -16577 195414 -16532
rect 195513 -16543 195514 -16532
rect 195722 -16537 195757 -16503
rect 195767 -16537 195768 -16492
rect 195867 -16503 195868 -16492
rect 196112 -16496 196147 -16462
rect 196157 -16496 196158 -16451
rect 196257 -16462 196258 -16451
rect 196268 -16496 196303 -16462
rect 196313 -16496 196314 -16451
rect 196413 -16462 196414 -16451
rect 196594 -16456 196629 -16422
rect 196666 -16456 196701 -16422
rect 196738 -16456 196773 -16422
rect 196882 -16456 196917 -16422
rect 196954 -16456 196989 -16422
rect 196991 -16456 197061 -16422
rect 197098 -16456 197133 -16422
rect 197168 -16456 197203 -16422
rect 196424 -16496 196459 -16462
rect 197464 -16491 197499 -16457
rect 197509 -16491 197510 -16446
rect 197609 -16457 197610 -16446
rect 197620 -16491 197655 -16457
rect 197665 -16491 197666 -16446
rect 197765 -16457 197766 -16446
rect 198341 -16451 198376 -16417
rect 198518 -16451 198553 -16417
rect 197776 -16491 197811 -16457
rect 195878 -16537 195913 -16503
rect 197157 -16505 197158 -16494
rect 195524 -16577 195559 -16543
rect 194437 -16621 194472 -16587
rect 194638 -16666 194673 -16632
rect 194761 -16637 194762 -16595
rect 195083 -16624 195118 -16590
rect 195722 -16620 195757 -16586
rect 195767 -16620 195768 -16575
rect 195867 -16586 195868 -16575
rect 196112 -16580 196147 -16546
rect 196157 -16580 196158 -16535
rect 196257 -16546 196258 -16535
rect 196268 -16580 196303 -16546
rect 196313 -16580 196314 -16535
rect 196413 -16546 196414 -16535
rect 196991 -16539 197026 -16505
rect 197168 -16539 197203 -16505
rect 196424 -16580 196459 -16546
rect 197311 -16565 197426 -16499
rect 197609 -16525 197610 -16499
rect 198006 -16517 198041 -16483
rect 198051 -16517 198052 -16472
rect 198151 -16483 198152 -16472
rect 198162 -16517 198197 -16483
rect 198207 -16517 198208 -16472
rect 198507 -16500 198508 -16489
rect 198712 -16494 198747 -16460
rect 198757 -16494 198758 -16449
rect 198857 -16460 198858 -16449
rect 199066 -16453 199101 -16419
rect 199111 -16453 199112 -16408
rect 199211 -16419 199212 -16408
rect 199392 -16413 199427 -16379
rect 199456 -16413 199499 -16379
rect 199501 -16413 199502 -16371
rect 199601 -16379 199602 -16371
rect 199536 -16413 199571 -16379
rect 199612 -16413 199647 -16379
rect 199657 -16413 199658 -16371
rect 199757 -16379 199758 -16371
rect 199706 -16413 199741 -16379
rect 199768 -16413 199813 -16379
rect 200808 -16408 200843 -16374
rect 200853 -16408 200854 -16363
rect 200953 -16374 200954 -16363
rect 200964 -16408 200999 -16374
rect 201009 -16408 201010 -16363
rect 201109 -16374 201110 -16363
rect 201685 -16367 201720 -16333
rect 201862 -16367 201897 -16333
rect 202455 -16336 202456 -16328
rect 202555 -16336 202556 -16328
rect 201120 -16408 201155 -16374
rect 199222 -16453 199257 -16419
rect 200501 -16422 200502 -16414
rect 201851 -16417 201852 -16406
rect 202056 -16410 202091 -16376
rect 202101 -16410 202102 -16365
rect 202201 -16376 202202 -16365
rect 202382 -16370 202445 -16336
rect 202454 -16370 202489 -16336
rect 202566 -16370 202601 -16336
rect 203291 -16360 203326 -16326
rect 203387 -16360 203422 -16326
rect 203483 -16360 203518 -16326
rect 203579 -16360 203614 -16326
rect 203675 -16360 203710 -16326
rect 203771 -16360 203806 -16326
rect 203867 -16360 203902 -16326
rect 205195 -16333 205196 -16322
rect 205372 -16327 205435 -16293
rect 205444 -16327 205479 -16293
rect 205556 -16327 205591 -16293
rect 206087 -16317 206122 -16283
rect 206183 -16317 206218 -16283
rect 206279 -16317 206314 -16283
rect 206375 -16317 206410 -16283
rect 206471 -16317 206506 -16283
rect 207496 -16324 207531 -16290
rect 207541 -16324 207542 -16279
rect 207641 -16290 207642 -16279
rect 207652 -16324 207687 -16290
rect 207697 -16324 207698 -16279
rect 207797 -16290 207798 -16279
rect 207976 -16284 208011 -16250
rect 208048 -16284 208083 -16250
rect 208120 -16284 208155 -16250
rect 208264 -16284 208299 -16250
rect 208336 -16284 208371 -16250
rect 208373 -16284 208443 -16250
rect 208480 -16284 208515 -16250
rect 208550 -16284 208585 -16250
rect 209077 -16274 209112 -16240
rect 209173 -16274 209208 -16240
rect 209269 -16274 209304 -16240
rect 210776 -16241 210811 -16207
rect 210840 -16241 210883 -16207
rect 210885 -16241 210886 -16199
rect 210985 -16207 210986 -16199
rect 210920 -16241 210955 -16207
rect 210996 -16241 211031 -16207
rect 211041 -16241 211042 -16199
rect 211141 -16207 211142 -16199
rect 211090 -16241 211125 -16207
rect 211152 -16241 211197 -16207
rect 212067 -16231 212102 -16197
rect 212163 -16231 212198 -16197
rect 212259 -16231 212294 -16197
rect 211883 -16250 211884 -16242
rect 207808 -16324 207843 -16290
rect 208789 -16293 208790 -16285
rect 208889 -16293 208890 -16285
rect 202212 -16410 202247 -16376
rect 198868 -16494 198903 -16460
rect 195878 -16620 195913 -16586
rect 197157 -16589 197158 -16578
rect 194407 -16689 194408 -16681
rect 194418 -16723 194453 -16689
rect 194638 -16734 194673 -16700
rect 193085 -16793 193120 -16759
rect 193288 -16838 193323 -16804
rect 193411 -16809 193412 -16767
rect 193733 -16796 193768 -16762
rect 193055 -16861 193056 -16853
rect 193066 -16895 193101 -16861
rect 193288 -16906 193323 -16872
rect 193055 -16961 193056 -16950
rect 193066 -16995 193101 -16961
rect 192003 -17045 192038 -17011
rect 192099 -17045 192134 -17011
rect 192195 -17045 192230 -17011
rect 192704 -17035 192739 -17001
rect 192776 -17035 192811 -17001
rect 192848 -17035 192883 -17001
rect 192920 -17029 192956 -17001
rect 193266 -17025 193301 -16991
rect 193311 -17025 193312 -16980
rect 192920 -17035 192955 -17029
rect 192357 -17088 192392 -17054
rect 192453 -17088 192488 -17054
rect 192549 -17088 192584 -17054
rect 193453 -17076 193454 -16809
rect 194082 -16819 194469 -16753
rect 193469 -16860 193504 -16826
rect 193818 -16832 193829 -16819
rect 193752 -16874 193829 -16832
rect 193880 -16874 194469 -16819
rect 194616 -16853 194651 -16819
rect 194661 -16853 194662 -16808
rect 193752 -16877 194469 -16874
rect 193469 -16928 193504 -16894
rect 193672 -16942 193707 -16908
rect 193717 -16942 193718 -16900
rect 193553 -16991 193554 -16980
rect 193564 -17025 193599 -16991
rect 193672 -17042 193707 -17008
rect 193717 -17042 193718 -16997
rect 193565 -17078 193600 -17044
rect 193637 -17078 193672 -17044
rect 193709 -17078 193744 -17044
rect 192711 -17131 192746 -17097
rect 192807 -17131 192842 -17097
rect 192903 -17131 192938 -17097
rect 192999 -17131 193034 -17097
rect 193095 -17131 193130 -17097
rect 193752 -17114 193897 -16877
rect 194082 -16899 194469 -16877
rect 194006 -16925 194469 -16899
rect 194803 -16904 194804 -16637
rect 194819 -16688 194854 -16654
rect 195433 -16691 195468 -16657
rect 196112 -16663 196147 -16629
rect 196157 -16663 196158 -16618
rect 196257 -16629 196258 -16618
rect 196268 -16663 196303 -16629
rect 196313 -16663 196314 -16618
rect 196413 -16629 196414 -16618
rect 196991 -16623 197026 -16589
rect 197168 -16623 197203 -16589
rect 197529 -16605 197564 -16571
rect 196424 -16663 196459 -16629
rect 196257 -16697 196258 -16671
rect 196656 -16689 196691 -16655
rect 196701 -16689 196702 -16644
rect 196801 -16655 196802 -16644
rect 196812 -16689 196847 -16655
rect 196857 -16689 196858 -16644
rect 197157 -16672 197158 -16661
rect 194819 -16756 194854 -16722
rect 195022 -16770 195057 -16736
rect 195067 -16770 195068 -16728
rect 195167 -16740 195168 -16729
rect 195787 -16734 195822 -16700
rect 195178 -16774 195213 -16740
rect 194903 -16819 194904 -16808
rect 195372 -16813 195407 -16779
rect 195417 -16813 195418 -16771
rect 195517 -16779 195518 -16771
rect 196177 -16777 196212 -16743
rect 195528 -16813 195563 -16779
rect 194914 -16853 194949 -16819
rect 195022 -16870 195057 -16836
rect 195067 -16870 195068 -16825
rect 195167 -16832 195168 -16821
rect 195178 -16866 195213 -16832
rect 195726 -16856 195761 -16822
rect 195771 -16856 195772 -16814
rect 195871 -16822 195872 -16814
rect 195882 -16856 195917 -16822
rect 194915 -16906 194950 -16872
rect 194987 -16906 195022 -16872
rect 195059 -16906 195094 -16872
rect 195372 -16913 195407 -16879
rect 195417 -16913 195418 -16868
rect 195517 -16879 195518 -16868
rect 195528 -16913 195563 -16879
rect 196112 -16895 196147 -16861
rect 196157 -16895 196158 -16853
rect 194006 -16959 194482 -16925
rect 195340 -16949 195375 -16915
rect 195412 -16949 195447 -16915
rect 195726 -16956 195761 -16922
rect 195771 -16956 195772 -16911
rect 195871 -16922 195872 -16911
rect 195882 -16956 195917 -16922
rect 194006 -16985 194469 -16959
rect 194010 -16993 194211 -16985
rect 194026 -17003 194195 -16993
rect 193752 -17140 193927 -17114
rect 193259 -17174 193294 -17140
rect 193355 -17174 193390 -17140
rect 193451 -17174 193486 -17140
rect 193547 -17174 193582 -17140
rect 193643 -17174 193678 -17140
rect 193739 -17174 193927 -17140
rect 193752 -17200 193927 -17174
rect 193952 -17174 194053 -17050
rect 193830 -17870 193865 -17200
rect 193952 -17228 193955 -17174
rect 193637 -17936 193782 -17924
rect 193305 -17970 193782 -17936
rect 193637 -17971 193782 -17970
rect 193818 -17971 193865 -17870
rect 193964 -17971 193999 -17174
rect 194222 -17971 194257 -17062
rect 194356 -17971 194391 -16985
rect 194609 -17002 194644 -16968
rect 194705 -17002 194740 -16968
rect 194801 -17002 194836 -16968
rect 194897 -17002 194932 -16968
rect 194993 -17002 195028 -16968
rect 195089 -17002 195124 -16968
rect 195185 -17002 195220 -16968
rect 195694 -16992 195729 -16958
rect 195766 -16992 195801 -16958
rect 196112 -16995 196147 -16961
rect 196157 -16995 196158 -16950
rect 196299 -17001 196300 -16697
rect 196991 -16706 197026 -16672
rect 197168 -16706 197203 -16672
rect 197464 -16723 197499 -16689
rect 197509 -16723 197510 -16681
rect 197651 -16753 197652 -16525
rect 198341 -16534 198376 -16500
rect 198518 -16534 198553 -16500
rect 198712 -16577 198747 -16543
rect 198757 -16577 198758 -16532
rect 198857 -16543 198858 -16532
rect 199066 -16537 199101 -16503
rect 199111 -16537 199112 -16492
rect 199211 -16503 199212 -16492
rect 199456 -16496 199491 -16462
rect 199501 -16496 199502 -16451
rect 199601 -16462 199602 -16451
rect 199612 -16496 199647 -16462
rect 199657 -16496 199658 -16451
rect 199757 -16462 199758 -16451
rect 199938 -16456 199973 -16422
rect 200010 -16456 200045 -16422
rect 200082 -16456 200117 -16422
rect 200226 -16456 200261 -16422
rect 200298 -16456 200333 -16422
rect 200335 -16456 200405 -16422
rect 200442 -16456 200477 -16422
rect 200512 -16456 200547 -16422
rect 199768 -16496 199803 -16462
rect 200808 -16491 200843 -16457
rect 200853 -16491 200854 -16446
rect 200953 -16457 200954 -16446
rect 200964 -16491 200999 -16457
rect 201009 -16491 201010 -16446
rect 201109 -16457 201110 -16446
rect 201685 -16451 201720 -16417
rect 201862 -16451 201897 -16417
rect 201120 -16491 201155 -16457
rect 199222 -16537 199257 -16503
rect 200501 -16505 200502 -16494
rect 198868 -16577 198903 -16543
rect 197781 -16621 197816 -16587
rect 197982 -16666 198017 -16632
rect 198105 -16637 198106 -16595
rect 198427 -16624 198462 -16590
rect 199066 -16620 199101 -16586
rect 199111 -16620 199112 -16575
rect 199211 -16586 199212 -16575
rect 199456 -16580 199491 -16546
rect 199501 -16580 199502 -16535
rect 199601 -16546 199602 -16535
rect 199612 -16580 199647 -16546
rect 199657 -16580 199658 -16535
rect 199757 -16546 199758 -16535
rect 200335 -16539 200370 -16505
rect 200512 -16539 200547 -16505
rect 199768 -16580 199803 -16546
rect 200655 -16565 200770 -16499
rect 200953 -16525 200954 -16499
rect 201350 -16517 201385 -16483
rect 201395 -16517 201396 -16472
rect 201495 -16483 201496 -16472
rect 201506 -16517 201541 -16483
rect 201551 -16517 201552 -16472
rect 201851 -16500 201852 -16489
rect 202056 -16494 202091 -16460
rect 202101 -16494 202102 -16449
rect 202201 -16460 202202 -16449
rect 202410 -16453 202445 -16419
rect 202455 -16453 202456 -16408
rect 202555 -16419 202556 -16408
rect 202736 -16413 202771 -16379
rect 202800 -16413 202843 -16379
rect 202845 -16413 202846 -16371
rect 202945 -16379 202946 -16371
rect 202880 -16413 202915 -16379
rect 202956 -16413 202991 -16379
rect 203001 -16413 203002 -16371
rect 203101 -16379 203102 -16371
rect 203050 -16413 203085 -16379
rect 203112 -16413 203157 -16379
rect 204152 -16408 204187 -16374
rect 204197 -16408 204198 -16363
rect 204297 -16374 204298 -16363
rect 204308 -16408 204343 -16374
rect 204353 -16408 204354 -16363
rect 204453 -16374 204454 -16363
rect 205029 -16367 205064 -16333
rect 205206 -16367 205241 -16333
rect 205799 -16336 205800 -16328
rect 205899 -16336 205900 -16328
rect 204464 -16408 204499 -16374
rect 202566 -16453 202601 -16419
rect 203845 -16422 203846 -16414
rect 205195 -16417 205196 -16406
rect 205400 -16410 205435 -16376
rect 205445 -16410 205446 -16365
rect 205545 -16376 205546 -16365
rect 205726 -16370 205789 -16336
rect 205798 -16370 205833 -16336
rect 205910 -16370 205945 -16336
rect 206635 -16360 206670 -16326
rect 206731 -16360 206766 -16326
rect 206827 -16360 206862 -16326
rect 206923 -16360 206958 -16326
rect 207019 -16360 207054 -16326
rect 207115 -16360 207150 -16326
rect 207211 -16360 207246 -16326
rect 208539 -16333 208540 -16322
rect 208716 -16327 208779 -16293
rect 208788 -16327 208823 -16293
rect 208900 -16327 208935 -16293
rect 209431 -16317 209466 -16283
rect 209527 -16317 209562 -16283
rect 209623 -16317 209658 -16283
rect 209719 -16317 209754 -16283
rect 209815 -16317 209850 -16283
rect 210840 -16324 210875 -16290
rect 210885 -16324 210886 -16279
rect 210985 -16290 210986 -16279
rect 210996 -16324 211031 -16290
rect 211041 -16324 211042 -16279
rect 211141 -16290 211142 -16279
rect 211320 -16284 211355 -16250
rect 211392 -16284 211427 -16250
rect 211464 -16284 211499 -16250
rect 211608 -16284 211643 -16250
rect 211680 -16284 211715 -16250
rect 211717 -16284 211787 -16250
rect 211824 -16284 211859 -16250
rect 211894 -16284 211929 -16250
rect 212421 -16274 212456 -16240
rect 212517 -16274 212552 -16240
rect 212613 -16274 212648 -16240
rect 211152 -16324 211187 -16290
rect 212133 -16293 212134 -16285
rect 212233 -16293 212234 -16285
rect 205556 -16410 205591 -16376
rect 202212 -16494 202247 -16460
rect 199222 -16620 199257 -16586
rect 200501 -16589 200502 -16578
rect 197751 -16689 197752 -16681
rect 197762 -16723 197797 -16689
rect 197982 -16734 198017 -16700
rect 196429 -16793 196464 -16759
rect 196632 -16838 196667 -16804
rect 196755 -16809 196756 -16767
rect 197077 -16796 197112 -16762
rect 196399 -16861 196400 -16853
rect 196410 -16895 196445 -16861
rect 196632 -16906 196667 -16872
rect 196399 -16961 196400 -16950
rect 196410 -16995 196445 -16961
rect 195347 -17045 195382 -17011
rect 195443 -17045 195478 -17011
rect 195539 -17045 195574 -17011
rect 196048 -17035 196083 -17001
rect 196120 -17035 196155 -17001
rect 196192 -17035 196227 -17001
rect 196264 -17029 196300 -17001
rect 196610 -17025 196645 -16991
rect 196655 -17025 196656 -16980
rect 196264 -17035 196299 -17029
rect 195701 -17088 195736 -17054
rect 195797 -17088 195832 -17054
rect 195893 -17088 195928 -17054
rect 196797 -17076 196798 -16809
rect 197426 -16819 197813 -16753
rect 196813 -16860 196848 -16826
rect 197162 -16832 197173 -16819
rect 197096 -16874 197173 -16832
rect 197224 -16874 197813 -16819
rect 197960 -16853 197995 -16819
rect 198005 -16853 198006 -16808
rect 197096 -16877 197813 -16874
rect 196813 -16928 196848 -16894
rect 197016 -16942 197051 -16908
rect 197061 -16942 197062 -16900
rect 196897 -16991 196898 -16980
rect 196908 -17025 196943 -16991
rect 197016 -17042 197051 -17008
rect 197061 -17042 197062 -16997
rect 196909 -17078 196944 -17044
rect 196981 -17078 197016 -17044
rect 197053 -17078 197088 -17044
rect 196055 -17131 196090 -17097
rect 196151 -17131 196186 -17097
rect 196247 -17131 196282 -17097
rect 196343 -17131 196378 -17097
rect 196439 -17131 196474 -17097
rect 197096 -17114 197241 -16877
rect 197426 -16899 197813 -16877
rect 197350 -16925 197813 -16899
rect 198147 -16904 198148 -16637
rect 198163 -16688 198198 -16654
rect 198777 -16691 198812 -16657
rect 199456 -16663 199491 -16629
rect 199501 -16663 199502 -16618
rect 199601 -16629 199602 -16618
rect 199612 -16663 199647 -16629
rect 199657 -16663 199658 -16618
rect 199757 -16629 199758 -16618
rect 200335 -16623 200370 -16589
rect 200512 -16623 200547 -16589
rect 200873 -16605 200908 -16571
rect 199768 -16663 199803 -16629
rect 199601 -16697 199602 -16671
rect 200000 -16689 200035 -16655
rect 200045 -16689 200046 -16644
rect 200145 -16655 200146 -16644
rect 200156 -16689 200191 -16655
rect 200201 -16689 200202 -16644
rect 200501 -16672 200502 -16661
rect 198163 -16756 198198 -16722
rect 198366 -16770 198401 -16736
rect 198411 -16770 198412 -16728
rect 198511 -16740 198512 -16729
rect 199131 -16734 199166 -16700
rect 198522 -16774 198557 -16740
rect 198247 -16819 198248 -16808
rect 198716 -16813 198751 -16779
rect 198761 -16813 198762 -16771
rect 198861 -16779 198862 -16771
rect 199521 -16777 199556 -16743
rect 198872 -16813 198907 -16779
rect 198258 -16853 198293 -16819
rect 198366 -16870 198401 -16836
rect 198411 -16870 198412 -16825
rect 198511 -16832 198512 -16821
rect 198522 -16866 198557 -16832
rect 199070 -16856 199105 -16822
rect 199115 -16856 199116 -16814
rect 199215 -16822 199216 -16814
rect 199226 -16856 199261 -16822
rect 198259 -16906 198294 -16872
rect 198331 -16906 198366 -16872
rect 198403 -16906 198438 -16872
rect 198716 -16913 198751 -16879
rect 198761 -16913 198762 -16868
rect 198861 -16879 198862 -16868
rect 198872 -16913 198907 -16879
rect 199456 -16895 199491 -16861
rect 199501 -16895 199502 -16853
rect 197350 -16959 197826 -16925
rect 198684 -16949 198719 -16915
rect 198756 -16949 198791 -16915
rect 199070 -16956 199105 -16922
rect 199115 -16956 199116 -16911
rect 199215 -16922 199216 -16911
rect 199226 -16956 199261 -16922
rect 197350 -16985 197813 -16959
rect 197354 -16993 197555 -16985
rect 197370 -17003 197539 -16993
rect 197096 -17140 197271 -17114
rect 196603 -17174 196638 -17140
rect 196699 -17174 196734 -17140
rect 196795 -17174 196830 -17140
rect 196891 -17174 196926 -17140
rect 196987 -17174 197022 -17140
rect 197083 -17174 197271 -17140
rect 197096 -17200 197271 -17174
rect 197296 -17174 197397 -17050
rect 197174 -17870 197209 -17200
rect 197296 -17228 197299 -17174
rect 196981 -17936 197126 -17924
rect 196649 -17970 197126 -17936
rect 196981 -17971 197126 -17970
rect 197162 -17971 197209 -17870
rect 197308 -17971 197343 -17174
rect 197566 -17971 197601 -17062
rect 197700 -17971 197735 -16985
rect 197953 -17002 197988 -16968
rect 198049 -17002 198084 -16968
rect 198145 -17002 198180 -16968
rect 198241 -17002 198276 -16968
rect 198337 -17002 198372 -16968
rect 198433 -17002 198468 -16968
rect 198529 -17002 198564 -16968
rect 199038 -16992 199073 -16958
rect 199110 -16992 199145 -16958
rect 199456 -16995 199491 -16961
rect 199501 -16995 199502 -16950
rect 199643 -17001 199644 -16697
rect 200335 -16706 200370 -16672
rect 200512 -16706 200547 -16672
rect 200808 -16723 200843 -16689
rect 200853 -16723 200854 -16681
rect 200995 -16753 200996 -16525
rect 201685 -16534 201720 -16500
rect 201862 -16534 201897 -16500
rect 202056 -16577 202091 -16543
rect 202101 -16577 202102 -16532
rect 202201 -16543 202202 -16532
rect 202410 -16537 202445 -16503
rect 202455 -16537 202456 -16492
rect 202555 -16503 202556 -16492
rect 202800 -16496 202835 -16462
rect 202845 -16496 202846 -16451
rect 202945 -16462 202946 -16451
rect 202956 -16496 202991 -16462
rect 203001 -16496 203002 -16451
rect 203101 -16462 203102 -16451
rect 203282 -16456 203317 -16422
rect 203354 -16456 203389 -16422
rect 203426 -16456 203461 -16422
rect 203570 -16456 203605 -16422
rect 203642 -16456 203677 -16422
rect 203679 -16456 203749 -16422
rect 203786 -16456 203821 -16422
rect 203856 -16456 203891 -16422
rect 203112 -16496 203147 -16462
rect 204152 -16491 204187 -16457
rect 204197 -16491 204198 -16446
rect 204297 -16457 204298 -16446
rect 204308 -16491 204343 -16457
rect 204353 -16491 204354 -16446
rect 204453 -16457 204454 -16446
rect 205029 -16451 205064 -16417
rect 205206 -16451 205241 -16417
rect 204464 -16491 204499 -16457
rect 202566 -16537 202601 -16503
rect 203845 -16505 203846 -16494
rect 202212 -16577 202247 -16543
rect 201125 -16621 201160 -16587
rect 201326 -16666 201361 -16632
rect 201449 -16637 201450 -16595
rect 201771 -16624 201806 -16590
rect 202410 -16620 202445 -16586
rect 202455 -16620 202456 -16575
rect 202555 -16586 202556 -16575
rect 202800 -16580 202835 -16546
rect 202845 -16580 202846 -16535
rect 202945 -16546 202946 -16535
rect 202956 -16580 202991 -16546
rect 203001 -16580 203002 -16535
rect 203101 -16546 203102 -16535
rect 203679 -16539 203714 -16505
rect 203856 -16539 203891 -16505
rect 203112 -16580 203147 -16546
rect 203999 -16565 204114 -16499
rect 204297 -16525 204298 -16499
rect 204694 -16517 204729 -16483
rect 204739 -16517 204740 -16472
rect 204839 -16483 204840 -16472
rect 204850 -16517 204885 -16483
rect 204895 -16517 204896 -16472
rect 205195 -16500 205196 -16489
rect 205400 -16494 205435 -16460
rect 205445 -16494 205446 -16449
rect 205545 -16460 205546 -16449
rect 205754 -16453 205789 -16419
rect 205799 -16453 205800 -16408
rect 205899 -16419 205900 -16408
rect 206080 -16413 206115 -16379
rect 206144 -16413 206187 -16379
rect 206189 -16413 206190 -16371
rect 206289 -16379 206290 -16371
rect 206224 -16413 206259 -16379
rect 206300 -16413 206335 -16379
rect 206345 -16413 206346 -16371
rect 206445 -16379 206446 -16371
rect 206394 -16413 206429 -16379
rect 206456 -16413 206501 -16379
rect 207496 -16408 207531 -16374
rect 207541 -16408 207542 -16363
rect 207641 -16374 207642 -16363
rect 207652 -16408 207687 -16374
rect 207697 -16408 207698 -16363
rect 207797 -16374 207798 -16363
rect 208373 -16367 208408 -16333
rect 208550 -16367 208585 -16333
rect 209143 -16336 209144 -16328
rect 209243 -16336 209244 -16328
rect 207808 -16408 207843 -16374
rect 205910 -16453 205945 -16419
rect 207189 -16422 207190 -16414
rect 208539 -16417 208540 -16406
rect 208744 -16410 208779 -16376
rect 208789 -16410 208790 -16365
rect 208889 -16376 208890 -16365
rect 209070 -16370 209133 -16336
rect 209142 -16370 209177 -16336
rect 209254 -16370 209289 -16336
rect 209979 -16360 210014 -16326
rect 210075 -16360 210110 -16326
rect 210171 -16360 210206 -16326
rect 210267 -16360 210302 -16326
rect 210363 -16360 210398 -16326
rect 210459 -16360 210494 -16326
rect 210555 -16360 210590 -16326
rect 211883 -16333 211884 -16322
rect 212060 -16327 212123 -16293
rect 212132 -16327 212167 -16293
rect 212244 -16327 212279 -16293
rect 212775 -16317 212810 -16283
rect 212871 -16317 212906 -16283
rect 212967 -16317 213002 -16283
rect 213063 -16317 213098 -16283
rect 213159 -16317 213194 -16283
rect 208900 -16410 208935 -16376
rect 205556 -16494 205591 -16460
rect 202566 -16620 202601 -16586
rect 203845 -16589 203846 -16578
rect 201095 -16689 201096 -16681
rect 201106 -16723 201141 -16689
rect 201326 -16734 201361 -16700
rect 199773 -16793 199808 -16759
rect 199976 -16838 200011 -16804
rect 200099 -16809 200100 -16767
rect 200421 -16796 200456 -16762
rect 199743 -16861 199744 -16853
rect 199754 -16895 199789 -16861
rect 199976 -16906 200011 -16872
rect 199743 -16961 199744 -16950
rect 199754 -16995 199789 -16961
rect 198691 -17045 198726 -17011
rect 198787 -17045 198822 -17011
rect 198883 -17045 198918 -17011
rect 199392 -17035 199427 -17001
rect 199464 -17035 199499 -17001
rect 199536 -17035 199571 -17001
rect 199608 -17029 199644 -17001
rect 199954 -17025 199989 -16991
rect 199999 -17025 200000 -16980
rect 199608 -17035 199643 -17029
rect 199045 -17088 199080 -17054
rect 199141 -17088 199176 -17054
rect 199237 -17088 199272 -17054
rect 200141 -17076 200142 -16809
rect 200770 -16819 201157 -16753
rect 200157 -16860 200192 -16826
rect 200506 -16832 200517 -16819
rect 200440 -16874 200517 -16832
rect 200568 -16874 201157 -16819
rect 201304 -16853 201339 -16819
rect 201349 -16853 201350 -16808
rect 200440 -16877 201157 -16874
rect 200157 -16928 200192 -16894
rect 200360 -16942 200395 -16908
rect 200405 -16942 200406 -16900
rect 200241 -16991 200242 -16980
rect 200252 -17025 200287 -16991
rect 200360 -17042 200395 -17008
rect 200405 -17042 200406 -16997
rect 200253 -17078 200288 -17044
rect 200325 -17078 200360 -17044
rect 200397 -17078 200432 -17044
rect 199399 -17131 199434 -17097
rect 199495 -17131 199530 -17097
rect 199591 -17131 199626 -17097
rect 199687 -17131 199722 -17097
rect 199783 -17131 199818 -17097
rect 200440 -17114 200585 -16877
rect 200770 -16899 201157 -16877
rect 200694 -16925 201157 -16899
rect 201491 -16904 201492 -16637
rect 201507 -16688 201542 -16654
rect 202121 -16691 202156 -16657
rect 202800 -16663 202835 -16629
rect 202845 -16663 202846 -16618
rect 202945 -16629 202946 -16618
rect 202956 -16663 202991 -16629
rect 203001 -16663 203002 -16618
rect 203101 -16629 203102 -16618
rect 203679 -16623 203714 -16589
rect 203856 -16623 203891 -16589
rect 204217 -16605 204252 -16571
rect 203112 -16663 203147 -16629
rect 202945 -16697 202946 -16671
rect 203344 -16689 203379 -16655
rect 203389 -16689 203390 -16644
rect 203489 -16655 203490 -16644
rect 203500 -16689 203535 -16655
rect 203545 -16689 203546 -16644
rect 203845 -16672 203846 -16661
rect 201507 -16756 201542 -16722
rect 201710 -16770 201745 -16736
rect 201755 -16770 201756 -16728
rect 201855 -16740 201856 -16729
rect 202475 -16734 202510 -16700
rect 201866 -16774 201901 -16740
rect 201591 -16819 201592 -16808
rect 202060 -16813 202095 -16779
rect 202105 -16813 202106 -16771
rect 202205 -16779 202206 -16771
rect 202865 -16777 202900 -16743
rect 202216 -16813 202251 -16779
rect 201602 -16853 201637 -16819
rect 201710 -16870 201745 -16836
rect 201755 -16870 201756 -16825
rect 201855 -16832 201856 -16821
rect 201866 -16866 201901 -16832
rect 202414 -16856 202449 -16822
rect 202459 -16856 202460 -16814
rect 202559 -16822 202560 -16814
rect 202570 -16856 202605 -16822
rect 201603 -16906 201638 -16872
rect 201675 -16906 201710 -16872
rect 201747 -16906 201782 -16872
rect 202060 -16913 202095 -16879
rect 202105 -16913 202106 -16868
rect 202205 -16879 202206 -16868
rect 202216 -16913 202251 -16879
rect 202800 -16895 202835 -16861
rect 202845 -16895 202846 -16853
rect 200694 -16959 201170 -16925
rect 202028 -16949 202063 -16915
rect 202100 -16949 202135 -16915
rect 202414 -16956 202449 -16922
rect 202459 -16956 202460 -16911
rect 202559 -16922 202560 -16911
rect 202570 -16956 202605 -16922
rect 200694 -16985 201157 -16959
rect 200698 -16993 200899 -16985
rect 200714 -17003 200883 -16993
rect 200440 -17140 200615 -17114
rect 199947 -17174 199982 -17140
rect 200043 -17174 200078 -17140
rect 200139 -17174 200174 -17140
rect 200235 -17174 200270 -17140
rect 200331 -17174 200366 -17140
rect 200427 -17174 200615 -17140
rect 200440 -17200 200615 -17174
rect 200640 -17174 200741 -17050
rect 200518 -17870 200553 -17200
rect 200640 -17228 200643 -17174
rect 200325 -17936 200470 -17924
rect 199993 -17970 200470 -17936
rect 200325 -17971 200470 -17970
rect 200506 -17971 200553 -17870
rect 200652 -17971 200687 -17174
rect 200910 -17971 200945 -17062
rect 201044 -17971 201079 -16985
rect 201297 -17002 201332 -16968
rect 201393 -17002 201428 -16968
rect 201489 -17002 201524 -16968
rect 201585 -17002 201620 -16968
rect 201681 -17002 201716 -16968
rect 201777 -17002 201812 -16968
rect 201873 -17002 201908 -16968
rect 202382 -16992 202417 -16958
rect 202454 -16992 202489 -16958
rect 202800 -16995 202835 -16961
rect 202845 -16995 202846 -16950
rect 202987 -17001 202988 -16697
rect 203679 -16706 203714 -16672
rect 203856 -16706 203891 -16672
rect 204152 -16723 204187 -16689
rect 204197 -16723 204198 -16681
rect 204339 -16753 204340 -16525
rect 205029 -16534 205064 -16500
rect 205206 -16534 205241 -16500
rect 205400 -16577 205435 -16543
rect 205445 -16577 205446 -16532
rect 205545 -16543 205546 -16532
rect 205754 -16537 205789 -16503
rect 205799 -16537 205800 -16492
rect 205899 -16503 205900 -16492
rect 206144 -16496 206179 -16462
rect 206189 -16496 206190 -16451
rect 206289 -16462 206290 -16451
rect 206300 -16496 206335 -16462
rect 206345 -16496 206346 -16451
rect 206445 -16462 206446 -16451
rect 206626 -16456 206661 -16422
rect 206698 -16456 206733 -16422
rect 206770 -16456 206805 -16422
rect 206914 -16456 206949 -16422
rect 206986 -16456 207021 -16422
rect 207023 -16456 207093 -16422
rect 207130 -16456 207165 -16422
rect 207200 -16456 207235 -16422
rect 206456 -16496 206491 -16462
rect 207496 -16491 207531 -16457
rect 207541 -16491 207542 -16446
rect 207641 -16457 207642 -16446
rect 207652 -16491 207687 -16457
rect 207697 -16491 207698 -16446
rect 207797 -16457 207798 -16446
rect 208373 -16451 208408 -16417
rect 208550 -16451 208585 -16417
rect 207808 -16491 207843 -16457
rect 205910 -16537 205945 -16503
rect 207189 -16505 207190 -16494
rect 205556 -16577 205591 -16543
rect 204469 -16621 204504 -16587
rect 204670 -16666 204705 -16632
rect 204793 -16637 204794 -16595
rect 205115 -16624 205150 -16590
rect 205754 -16620 205789 -16586
rect 205799 -16620 205800 -16575
rect 205899 -16586 205900 -16575
rect 206144 -16580 206179 -16546
rect 206189 -16580 206190 -16535
rect 206289 -16546 206290 -16535
rect 206300 -16580 206335 -16546
rect 206345 -16580 206346 -16535
rect 206445 -16546 206446 -16535
rect 207023 -16539 207058 -16505
rect 207200 -16539 207235 -16505
rect 206456 -16580 206491 -16546
rect 207343 -16565 207458 -16499
rect 207641 -16525 207642 -16499
rect 208038 -16517 208073 -16483
rect 208083 -16517 208084 -16472
rect 208183 -16483 208184 -16472
rect 208194 -16517 208229 -16483
rect 208239 -16517 208240 -16472
rect 208539 -16500 208540 -16489
rect 208744 -16494 208779 -16460
rect 208789 -16494 208790 -16449
rect 208889 -16460 208890 -16449
rect 209098 -16453 209133 -16419
rect 209143 -16453 209144 -16408
rect 209243 -16419 209244 -16408
rect 209424 -16413 209459 -16379
rect 209488 -16413 209531 -16379
rect 209533 -16413 209534 -16371
rect 209633 -16379 209634 -16371
rect 209568 -16413 209603 -16379
rect 209644 -16413 209679 -16379
rect 209689 -16413 209690 -16371
rect 209789 -16379 209790 -16371
rect 209738 -16413 209773 -16379
rect 209800 -16413 209845 -16379
rect 210840 -16408 210875 -16374
rect 210885 -16408 210886 -16363
rect 210985 -16374 210986 -16363
rect 210996 -16408 211031 -16374
rect 211041 -16408 211042 -16363
rect 211141 -16374 211142 -16363
rect 211717 -16367 211752 -16333
rect 211894 -16367 211929 -16333
rect 212487 -16336 212488 -16328
rect 212587 -16336 212588 -16328
rect 211152 -16408 211187 -16374
rect 209254 -16453 209289 -16419
rect 210533 -16422 210534 -16414
rect 211883 -16417 211884 -16406
rect 212088 -16410 212123 -16376
rect 212133 -16410 212134 -16365
rect 212233 -16376 212234 -16365
rect 212414 -16370 212477 -16336
rect 212486 -16370 212521 -16336
rect 212598 -16370 212633 -16336
rect 213323 -16360 213358 -16326
rect 213419 -16360 213454 -16326
rect 213515 -16360 213550 -16326
rect 213611 -16360 213646 -16326
rect 213707 -16360 213742 -16326
rect 213803 -16360 213838 -16326
rect 213899 -16360 213934 -16326
rect 212244 -16410 212279 -16376
rect 208900 -16494 208935 -16460
rect 205910 -16620 205945 -16586
rect 207189 -16589 207190 -16578
rect 204439 -16689 204440 -16681
rect 204450 -16723 204485 -16689
rect 204670 -16734 204705 -16700
rect 203117 -16793 203152 -16759
rect 203320 -16838 203355 -16804
rect 203443 -16809 203444 -16767
rect 203765 -16796 203800 -16762
rect 203087 -16861 203088 -16853
rect 203098 -16895 203133 -16861
rect 203320 -16906 203355 -16872
rect 203087 -16961 203088 -16950
rect 203098 -16995 203133 -16961
rect 202035 -17045 202070 -17011
rect 202131 -17045 202166 -17011
rect 202227 -17045 202262 -17011
rect 202736 -17035 202771 -17001
rect 202808 -17035 202843 -17001
rect 202880 -17035 202915 -17001
rect 202952 -17029 202988 -17001
rect 203298 -17025 203333 -16991
rect 203343 -17025 203344 -16980
rect 202952 -17035 202987 -17029
rect 202389 -17088 202424 -17054
rect 202485 -17088 202520 -17054
rect 202581 -17088 202616 -17054
rect 203485 -17076 203486 -16809
rect 204114 -16819 204501 -16753
rect 203501 -16860 203536 -16826
rect 203850 -16832 203861 -16819
rect 203784 -16874 203861 -16832
rect 203912 -16874 204501 -16819
rect 204648 -16853 204683 -16819
rect 204693 -16853 204694 -16808
rect 203784 -16877 204501 -16874
rect 203501 -16928 203536 -16894
rect 203704 -16942 203739 -16908
rect 203749 -16942 203750 -16900
rect 203585 -16991 203586 -16980
rect 203596 -17025 203631 -16991
rect 203704 -17042 203739 -17008
rect 203749 -17042 203750 -16997
rect 203597 -17078 203632 -17044
rect 203669 -17078 203704 -17044
rect 203741 -17078 203776 -17044
rect 202743 -17131 202778 -17097
rect 202839 -17131 202874 -17097
rect 202935 -17131 202970 -17097
rect 203031 -17131 203066 -17097
rect 203127 -17131 203162 -17097
rect 203784 -17114 203929 -16877
rect 204114 -16899 204501 -16877
rect 204038 -16925 204501 -16899
rect 204835 -16904 204836 -16637
rect 204851 -16688 204886 -16654
rect 205465 -16691 205500 -16657
rect 206144 -16663 206179 -16629
rect 206189 -16663 206190 -16618
rect 206289 -16629 206290 -16618
rect 206300 -16663 206335 -16629
rect 206345 -16663 206346 -16618
rect 206445 -16629 206446 -16618
rect 207023 -16623 207058 -16589
rect 207200 -16623 207235 -16589
rect 207561 -16605 207596 -16571
rect 206456 -16663 206491 -16629
rect 206289 -16697 206290 -16671
rect 206688 -16689 206723 -16655
rect 206733 -16689 206734 -16644
rect 206833 -16655 206834 -16644
rect 206844 -16689 206879 -16655
rect 206889 -16689 206890 -16644
rect 207189 -16672 207190 -16661
rect 204851 -16756 204886 -16722
rect 205054 -16770 205089 -16736
rect 205099 -16770 205100 -16728
rect 205199 -16740 205200 -16729
rect 205819 -16734 205854 -16700
rect 205210 -16774 205245 -16740
rect 204935 -16819 204936 -16808
rect 205404 -16813 205439 -16779
rect 205449 -16813 205450 -16771
rect 205549 -16779 205550 -16771
rect 206209 -16777 206244 -16743
rect 205560 -16813 205595 -16779
rect 204946 -16853 204981 -16819
rect 205054 -16870 205089 -16836
rect 205099 -16870 205100 -16825
rect 205199 -16832 205200 -16821
rect 205210 -16866 205245 -16832
rect 205758 -16856 205793 -16822
rect 205803 -16856 205804 -16814
rect 205903 -16822 205904 -16814
rect 205914 -16856 205949 -16822
rect 204947 -16906 204982 -16872
rect 205019 -16906 205054 -16872
rect 205091 -16906 205126 -16872
rect 205404 -16913 205439 -16879
rect 205449 -16913 205450 -16868
rect 205549 -16879 205550 -16868
rect 205560 -16913 205595 -16879
rect 206144 -16895 206179 -16861
rect 206189 -16895 206190 -16853
rect 204038 -16959 204514 -16925
rect 205372 -16949 205407 -16915
rect 205444 -16949 205479 -16915
rect 205758 -16956 205793 -16922
rect 205803 -16956 205804 -16911
rect 205903 -16922 205904 -16911
rect 205914 -16956 205949 -16922
rect 204038 -16985 204501 -16959
rect 204042 -16993 204243 -16985
rect 204058 -17003 204227 -16993
rect 203784 -17140 203959 -17114
rect 203291 -17174 203326 -17140
rect 203387 -17174 203422 -17140
rect 203483 -17174 203518 -17140
rect 203579 -17174 203614 -17140
rect 203675 -17174 203710 -17140
rect 203771 -17174 203959 -17140
rect 203784 -17200 203959 -17174
rect 203984 -17174 204085 -17050
rect 203862 -17870 203897 -17200
rect 203984 -17228 203987 -17174
rect 203669 -17936 203814 -17924
rect 203337 -17970 203814 -17936
rect 203669 -17971 203814 -17970
rect 203850 -17971 203897 -17870
rect 203996 -17971 204031 -17174
rect 204254 -17971 204289 -17062
rect 204388 -17971 204423 -16985
rect 204641 -17002 204676 -16968
rect 204737 -17002 204772 -16968
rect 204833 -17002 204868 -16968
rect 204929 -17002 204964 -16968
rect 205025 -17002 205060 -16968
rect 205121 -17002 205156 -16968
rect 205217 -17002 205252 -16968
rect 205726 -16992 205761 -16958
rect 205798 -16992 205833 -16958
rect 206144 -16995 206179 -16961
rect 206189 -16995 206190 -16950
rect 206331 -17001 206332 -16697
rect 207023 -16706 207058 -16672
rect 207200 -16706 207235 -16672
rect 207496 -16723 207531 -16689
rect 207541 -16723 207542 -16681
rect 207683 -16753 207684 -16525
rect 208373 -16534 208408 -16500
rect 208550 -16534 208585 -16500
rect 208744 -16577 208779 -16543
rect 208789 -16577 208790 -16532
rect 208889 -16543 208890 -16532
rect 209098 -16537 209133 -16503
rect 209143 -16537 209144 -16492
rect 209243 -16503 209244 -16492
rect 209488 -16496 209523 -16462
rect 209533 -16496 209534 -16451
rect 209633 -16462 209634 -16451
rect 209644 -16496 209679 -16462
rect 209689 -16496 209690 -16451
rect 209789 -16462 209790 -16451
rect 209970 -16456 210005 -16422
rect 210042 -16456 210077 -16422
rect 210114 -16456 210149 -16422
rect 210258 -16456 210293 -16422
rect 210330 -16456 210365 -16422
rect 210367 -16456 210437 -16422
rect 210474 -16456 210509 -16422
rect 210544 -16456 210579 -16422
rect 209800 -16496 209835 -16462
rect 210840 -16491 210875 -16457
rect 210885 -16491 210886 -16446
rect 210985 -16457 210986 -16446
rect 210996 -16491 211031 -16457
rect 211041 -16491 211042 -16446
rect 211141 -16457 211142 -16446
rect 211717 -16451 211752 -16417
rect 211894 -16451 211929 -16417
rect 211152 -16491 211187 -16457
rect 209254 -16537 209289 -16503
rect 210533 -16505 210534 -16494
rect 208900 -16577 208935 -16543
rect 207813 -16621 207848 -16587
rect 208014 -16666 208049 -16632
rect 208137 -16637 208138 -16595
rect 208459 -16624 208494 -16590
rect 209098 -16620 209133 -16586
rect 209143 -16620 209144 -16575
rect 209243 -16586 209244 -16575
rect 209488 -16580 209523 -16546
rect 209533 -16580 209534 -16535
rect 209633 -16546 209634 -16535
rect 209644 -16580 209679 -16546
rect 209689 -16580 209690 -16535
rect 209789 -16546 209790 -16535
rect 210367 -16539 210402 -16505
rect 210544 -16539 210579 -16505
rect 209800 -16580 209835 -16546
rect 210687 -16565 210802 -16499
rect 210985 -16525 210986 -16499
rect 211382 -16517 211417 -16483
rect 211427 -16517 211428 -16472
rect 211527 -16483 211528 -16472
rect 211538 -16517 211573 -16483
rect 211583 -16517 211584 -16472
rect 211883 -16500 211884 -16489
rect 212088 -16494 212123 -16460
rect 212133 -16494 212134 -16449
rect 212233 -16460 212234 -16449
rect 212442 -16453 212477 -16419
rect 212487 -16453 212488 -16408
rect 212587 -16419 212588 -16408
rect 212768 -16413 212803 -16379
rect 212832 -16413 212875 -16379
rect 212877 -16413 212878 -16371
rect 212977 -16379 212978 -16371
rect 212912 -16413 212947 -16379
rect 212988 -16413 213023 -16379
rect 213033 -16413 213034 -16371
rect 213133 -16379 213134 -16371
rect 213082 -16413 213117 -16379
rect 213144 -16413 213189 -16379
rect 212598 -16453 212633 -16419
rect 213877 -16422 213878 -16414
rect 212244 -16494 212279 -16460
rect 209254 -16620 209289 -16586
rect 210533 -16589 210534 -16578
rect 207783 -16689 207784 -16681
rect 207794 -16723 207829 -16689
rect 208014 -16734 208049 -16700
rect 206461 -16793 206496 -16759
rect 206664 -16838 206699 -16804
rect 206787 -16809 206788 -16767
rect 207109 -16796 207144 -16762
rect 206431 -16861 206432 -16853
rect 206442 -16895 206477 -16861
rect 206664 -16906 206699 -16872
rect 206431 -16961 206432 -16950
rect 206442 -16995 206477 -16961
rect 205379 -17045 205414 -17011
rect 205475 -17045 205510 -17011
rect 205571 -17045 205606 -17011
rect 206080 -17035 206115 -17001
rect 206152 -17035 206187 -17001
rect 206224 -17035 206259 -17001
rect 206296 -17029 206332 -17001
rect 206642 -17025 206677 -16991
rect 206687 -17025 206688 -16980
rect 206296 -17035 206331 -17029
rect 205733 -17088 205768 -17054
rect 205829 -17088 205864 -17054
rect 205925 -17088 205960 -17054
rect 206829 -17076 206830 -16809
rect 207458 -16819 207845 -16753
rect 206845 -16860 206880 -16826
rect 207194 -16832 207205 -16819
rect 207128 -16874 207205 -16832
rect 207256 -16874 207845 -16819
rect 207992 -16853 208027 -16819
rect 208037 -16853 208038 -16808
rect 207128 -16877 207845 -16874
rect 206845 -16928 206880 -16894
rect 207048 -16942 207083 -16908
rect 207093 -16942 207094 -16900
rect 206929 -16991 206930 -16980
rect 206940 -17025 206975 -16991
rect 207048 -17042 207083 -17008
rect 207093 -17042 207094 -16997
rect 206941 -17078 206976 -17044
rect 207013 -17078 207048 -17044
rect 207085 -17078 207120 -17044
rect 206087 -17131 206122 -17097
rect 206183 -17131 206218 -17097
rect 206279 -17131 206314 -17097
rect 206375 -17131 206410 -17097
rect 206471 -17131 206506 -17097
rect 207128 -17114 207273 -16877
rect 207458 -16899 207845 -16877
rect 207382 -16925 207845 -16899
rect 208179 -16904 208180 -16637
rect 208195 -16688 208230 -16654
rect 208809 -16691 208844 -16657
rect 209488 -16663 209523 -16629
rect 209533 -16663 209534 -16618
rect 209633 -16629 209634 -16618
rect 209644 -16663 209679 -16629
rect 209689 -16663 209690 -16618
rect 209789 -16629 209790 -16618
rect 210367 -16623 210402 -16589
rect 210544 -16623 210579 -16589
rect 210905 -16605 210940 -16571
rect 209800 -16663 209835 -16629
rect 209633 -16697 209634 -16671
rect 210032 -16689 210067 -16655
rect 210077 -16689 210078 -16644
rect 210177 -16655 210178 -16644
rect 210188 -16689 210223 -16655
rect 210233 -16689 210234 -16644
rect 210533 -16672 210534 -16661
rect 208195 -16756 208230 -16722
rect 208398 -16770 208433 -16736
rect 208443 -16770 208444 -16728
rect 208543 -16740 208544 -16729
rect 209163 -16734 209198 -16700
rect 208554 -16774 208589 -16740
rect 208279 -16819 208280 -16808
rect 208748 -16813 208783 -16779
rect 208793 -16813 208794 -16771
rect 208893 -16779 208894 -16771
rect 209553 -16777 209588 -16743
rect 208904 -16813 208939 -16779
rect 208290 -16853 208325 -16819
rect 208398 -16870 208433 -16836
rect 208443 -16870 208444 -16825
rect 208543 -16832 208544 -16821
rect 208554 -16866 208589 -16832
rect 209102 -16856 209137 -16822
rect 209147 -16856 209148 -16814
rect 209247 -16822 209248 -16814
rect 209258 -16856 209293 -16822
rect 208291 -16906 208326 -16872
rect 208363 -16906 208398 -16872
rect 208435 -16906 208470 -16872
rect 208748 -16913 208783 -16879
rect 208793 -16913 208794 -16868
rect 208893 -16879 208894 -16868
rect 208904 -16913 208939 -16879
rect 209488 -16895 209523 -16861
rect 209533 -16895 209534 -16853
rect 207382 -16959 207858 -16925
rect 208716 -16949 208751 -16915
rect 208788 -16949 208823 -16915
rect 209102 -16956 209137 -16922
rect 209147 -16956 209148 -16911
rect 209247 -16922 209248 -16911
rect 209258 -16956 209293 -16922
rect 207382 -16985 207845 -16959
rect 207386 -16993 207587 -16985
rect 207402 -17003 207571 -16993
rect 207128 -17140 207303 -17114
rect 206635 -17174 206670 -17140
rect 206731 -17174 206766 -17140
rect 206827 -17174 206862 -17140
rect 206923 -17174 206958 -17140
rect 207019 -17174 207054 -17140
rect 207115 -17174 207303 -17140
rect 207128 -17200 207303 -17174
rect 207328 -17174 207429 -17050
rect 207206 -17870 207241 -17200
rect 207328 -17228 207331 -17174
rect 207013 -17936 207158 -17924
rect 206681 -17970 207158 -17936
rect 207013 -17971 207158 -17970
rect 207194 -17971 207241 -17870
rect 207340 -17971 207375 -17174
rect 207598 -17971 207633 -17062
rect 207732 -17971 207767 -16985
rect 207985 -17002 208020 -16968
rect 208081 -17002 208116 -16968
rect 208177 -17002 208212 -16968
rect 208273 -17002 208308 -16968
rect 208369 -17002 208404 -16968
rect 208465 -17002 208500 -16968
rect 208561 -17002 208596 -16968
rect 209070 -16992 209105 -16958
rect 209142 -16992 209177 -16958
rect 209488 -16995 209523 -16961
rect 209533 -16995 209534 -16950
rect 209675 -17001 209676 -16697
rect 210367 -16706 210402 -16672
rect 210544 -16706 210579 -16672
rect 210840 -16723 210875 -16689
rect 210885 -16723 210886 -16681
rect 211027 -16753 211028 -16525
rect 211717 -16534 211752 -16500
rect 211894 -16534 211929 -16500
rect 212088 -16577 212123 -16543
rect 212133 -16577 212134 -16532
rect 212233 -16543 212234 -16532
rect 212442 -16537 212477 -16503
rect 212487 -16537 212488 -16492
rect 212587 -16503 212588 -16492
rect 212832 -16496 212867 -16462
rect 212877 -16496 212878 -16451
rect 212977 -16462 212978 -16451
rect 212988 -16496 213023 -16462
rect 213033 -16496 213034 -16451
rect 213133 -16462 213134 -16451
rect 213314 -16456 213349 -16422
rect 213386 -16456 213421 -16422
rect 213458 -16456 213493 -16422
rect 213602 -16456 213637 -16422
rect 213674 -16456 213709 -16422
rect 213711 -16456 213781 -16422
rect 213818 -16456 213853 -16422
rect 213888 -16456 213923 -16422
rect 213144 -16496 213179 -16462
rect 212598 -16537 212633 -16503
rect 213877 -16505 213878 -16494
rect 212244 -16577 212279 -16543
rect 211157 -16621 211192 -16587
rect 211358 -16666 211393 -16632
rect 211481 -16637 211482 -16595
rect 211803 -16624 211838 -16590
rect 212442 -16620 212477 -16586
rect 212487 -16620 212488 -16575
rect 212587 -16586 212588 -16575
rect 212832 -16580 212867 -16546
rect 212877 -16580 212878 -16535
rect 212977 -16546 212978 -16535
rect 212988 -16580 213023 -16546
rect 213033 -16580 213034 -16535
rect 213133 -16546 213134 -16535
rect 213711 -16539 213746 -16505
rect 213888 -16539 213923 -16505
rect 213144 -16580 213179 -16546
rect 214031 -16565 214147 -16499
rect 217375 -16565 217491 -16499
rect 220719 -16565 220835 -16499
rect 224063 -16565 224179 -16499
rect 227407 -16565 227523 -16499
rect 230751 -16565 230867 -16499
rect 234095 -16565 234211 -16499
rect 237439 -16565 237555 -16499
rect 240783 -16565 240899 -16499
rect 244127 -16565 244243 -16499
rect 247471 -16565 247587 -16499
rect 250815 -16565 250931 -16499
rect 254159 -16565 254275 -16499
rect 257503 -16565 257619 -16499
rect 260847 -16565 260963 -16499
rect 264191 -16565 264307 -16499
rect 267535 -16565 267651 -16499
rect 270879 -16565 270995 -16499
rect 274223 -16565 274339 -16499
rect 277567 -16565 277683 -16499
rect 280911 -16565 281027 -16499
rect 284255 -16565 284371 -16499
rect 287599 -16565 287715 -16499
rect 290943 -16565 291059 -16499
rect 294287 -16565 294403 -16499
rect 297631 -16565 297747 -16499
rect 300975 -16565 301091 -16499
rect 304319 -16565 304435 -16499
rect 307663 -16565 307779 -16499
rect 311007 -16565 311123 -16499
rect 314351 -16565 314467 -16499
rect 317695 -16565 317811 -16499
rect 321039 -16565 321155 -16499
rect 324383 -16565 324499 -16499
rect 327727 -16565 327843 -16499
rect 331071 -16565 331187 -16499
rect 334415 -16565 334531 -16499
rect 337759 -16565 337875 -16499
rect 341103 -16565 341219 -16499
rect 344447 -16565 344563 -16499
rect 347791 -16565 347907 -16499
rect 351135 -16565 351251 -16499
rect 354479 -16565 354595 -16499
rect 357823 -16565 357939 -16499
rect 361167 -16565 361283 -16499
rect 364511 -16565 364627 -16499
rect 367855 -16565 367971 -16499
rect 371199 -16565 371315 -16499
rect 374543 -16565 374659 -16499
rect 377887 -16565 378003 -16499
rect 381231 -16565 381347 -16499
rect 384575 -16565 384691 -16499
rect 387919 -16565 388035 -16499
rect 391263 -16565 391379 -16499
rect 394607 -16565 394723 -16499
rect 397951 -16565 398067 -16499
rect 401295 -16565 401411 -16499
rect 404639 -16565 404755 -16499
rect 407983 -16565 408099 -16499
rect 411327 -16565 411443 -16499
rect 414671 -16565 414787 -16499
rect 418015 -16565 418131 -16499
rect 421359 -16565 421475 -16499
rect 424703 -16565 424819 -16499
rect 212598 -16620 212633 -16586
rect 213877 -16589 213878 -16578
rect 211127 -16689 211128 -16681
rect 211138 -16723 211173 -16689
rect 211358 -16734 211393 -16700
rect 209805 -16793 209840 -16759
rect 210008 -16838 210043 -16804
rect 210131 -16809 210132 -16767
rect 210453 -16796 210488 -16762
rect 209775 -16861 209776 -16853
rect 209786 -16895 209821 -16861
rect 210008 -16906 210043 -16872
rect 209775 -16961 209776 -16950
rect 209786 -16995 209821 -16961
rect 208723 -17045 208758 -17011
rect 208819 -17045 208854 -17011
rect 208915 -17045 208950 -17011
rect 209424 -17035 209459 -17001
rect 209496 -17035 209531 -17001
rect 209568 -17035 209603 -17001
rect 209640 -17029 209676 -17001
rect 209986 -17025 210021 -16991
rect 210031 -17025 210032 -16980
rect 209640 -17035 209675 -17029
rect 209077 -17088 209112 -17054
rect 209173 -17088 209208 -17054
rect 209269 -17088 209304 -17054
rect 210173 -17076 210174 -16809
rect 210802 -16819 211189 -16753
rect 210189 -16860 210224 -16826
rect 210538 -16832 210549 -16819
rect 210472 -16874 210549 -16832
rect 210600 -16874 211189 -16819
rect 211336 -16853 211371 -16819
rect 211381 -16853 211382 -16808
rect 210472 -16877 211189 -16874
rect 210189 -16928 210224 -16894
rect 210392 -16942 210427 -16908
rect 210437 -16942 210438 -16900
rect 210273 -16991 210274 -16980
rect 210284 -17025 210319 -16991
rect 210392 -17042 210427 -17008
rect 210437 -17042 210438 -16997
rect 210285 -17078 210320 -17044
rect 210357 -17078 210392 -17044
rect 210429 -17078 210464 -17044
rect 209431 -17131 209466 -17097
rect 209527 -17131 209562 -17097
rect 209623 -17131 209658 -17097
rect 209719 -17131 209754 -17097
rect 209815 -17131 209850 -17097
rect 210472 -17114 210617 -16877
rect 210802 -16899 211189 -16877
rect 210726 -16925 211189 -16899
rect 211523 -16904 211524 -16637
rect 211539 -16688 211574 -16654
rect 212153 -16691 212188 -16657
rect 212832 -16663 212867 -16629
rect 212877 -16663 212878 -16618
rect 212977 -16629 212978 -16618
rect 212988 -16663 213023 -16629
rect 213033 -16663 213034 -16618
rect 213133 -16629 213134 -16618
rect 213711 -16623 213746 -16589
rect 213888 -16623 213923 -16589
rect 213144 -16663 213179 -16629
rect 212977 -16697 212978 -16671
rect 213376 -16689 213411 -16655
rect 213421 -16689 213422 -16644
rect 213521 -16655 213522 -16644
rect 213532 -16689 213567 -16655
rect 213577 -16689 213578 -16644
rect 213877 -16672 213878 -16661
rect 211539 -16756 211574 -16722
rect 211742 -16770 211777 -16736
rect 211787 -16770 211788 -16728
rect 211887 -16740 211888 -16729
rect 212507 -16734 212542 -16700
rect 211898 -16774 211933 -16740
rect 211623 -16819 211624 -16808
rect 212092 -16813 212127 -16779
rect 212137 -16813 212138 -16771
rect 212237 -16779 212238 -16771
rect 212897 -16777 212932 -16743
rect 212248 -16813 212283 -16779
rect 211634 -16853 211669 -16819
rect 211742 -16870 211777 -16836
rect 211787 -16870 211788 -16825
rect 211887 -16832 211888 -16821
rect 211898 -16866 211933 -16832
rect 212446 -16856 212481 -16822
rect 212491 -16856 212492 -16814
rect 212591 -16822 212592 -16814
rect 212602 -16856 212637 -16822
rect 211635 -16906 211670 -16872
rect 211707 -16906 211742 -16872
rect 211779 -16906 211814 -16872
rect 212092 -16913 212127 -16879
rect 212137 -16913 212138 -16868
rect 212237 -16879 212238 -16868
rect 212248 -16913 212283 -16879
rect 212832 -16895 212867 -16861
rect 212877 -16895 212878 -16853
rect 210726 -16959 211202 -16925
rect 212060 -16949 212095 -16915
rect 212132 -16949 212167 -16915
rect 212446 -16956 212481 -16922
rect 212491 -16956 212492 -16911
rect 212591 -16922 212592 -16911
rect 212602 -16956 212637 -16922
rect 210726 -16985 211189 -16959
rect 210730 -16993 210931 -16985
rect 210746 -17003 210915 -16993
rect 210472 -17140 210647 -17114
rect 209979 -17174 210014 -17140
rect 210075 -17174 210110 -17140
rect 210171 -17174 210206 -17140
rect 210267 -17174 210302 -17140
rect 210363 -17174 210398 -17140
rect 210459 -17174 210647 -17140
rect 210472 -17200 210647 -17174
rect 210672 -17174 210773 -17050
rect 210550 -17870 210585 -17200
rect 210672 -17228 210675 -17174
rect 210357 -17936 210502 -17924
rect 210025 -17970 210502 -17936
rect 210357 -17971 210502 -17970
rect 210538 -17971 210585 -17870
rect 210684 -17971 210719 -17174
rect 210942 -17971 210977 -17062
rect 211076 -17971 211111 -16985
rect 211329 -17002 211364 -16968
rect 211425 -17002 211460 -16968
rect 211521 -17002 211556 -16968
rect 211617 -17002 211652 -16968
rect 211713 -17002 211748 -16968
rect 211809 -17002 211844 -16968
rect 211905 -17002 211940 -16968
rect 212414 -16992 212449 -16958
rect 212486 -16992 212521 -16958
rect 212832 -16995 212867 -16961
rect 212877 -16995 212878 -16950
rect 213019 -17001 213020 -16697
rect 213711 -16706 213746 -16672
rect 213888 -16706 213923 -16672
rect 213149 -16793 213184 -16759
rect 213352 -16838 213387 -16804
rect 213475 -16809 213476 -16767
rect 213797 -16796 213832 -16762
rect 213119 -16861 213120 -16853
rect 213130 -16895 213165 -16861
rect 213352 -16906 213387 -16872
rect 213119 -16961 213120 -16950
rect 213130 -16995 213165 -16961
rect 212067 -17045 212102 -17011
rect 212163 -17045 212198 -17011
rect 212259 -17045 212294 -17011
rect 212768 -17035 212803 -17001
rect 212840 -17035 212875 -17001
rect 212912 -17035 212947 -17001
rect 212984 -17029 213020 -17001
rect 213330 -17025 213365 -16991
rect 213375 -17025 213376 -16980
rect 212984 -17035 213019 -17029
rect 212421 -17088 212456 -17054
rect 212517 -17088 212552 -17054
rect 212613 -17088 212648 -17054
rect 213517 -17076 213518 -16809
rect 214147 -16819 214533 -16753
rect 217491 -16819 217877 -16753
rect 220835 -16819 221221 -16753
rect 224179 -16819 224565 -16753
rect 227523 -16819 227909 -16753
rect 230867 -16819 231253 -16753
rect 234211 -16819 234597 -16753
rect 237555 -16819 237941 -16753
rect 240899 -16819 241285 -16753
rect 244243 -16819 244629 -16753
rect 247587 -16819 247973 -16753
rect 250931 -16819 251317 -16753
rect 254275 -16819 254661 -16753
rect 257619 -16819 258005 -16753
rect 260963 -16819 261349 -16753
rect 264307 -16819 264693 -16753
rect 267651 -16819 268037 -16753
rect 270995 -16819 271381 -16753
rect 274339 -16819 274725 -16753
rect 277683 -16819 278069 -16753
rect 281027 -16819 281413 -16753
rect 284371 -16819 284757 -16753
rect 287715 -16819 288101 -16753
rect 291059 -16819 291445 -16753
rect 294403 -16819 294789 -16753
rect 297747 -16819 298133 -16753
rect 301091 -16819 301477 -16753
rect 304435 -16819 304821 -16753
rect 307779 -16819 308165 -16753
rect 311123 -16819 311509 -16753
rect 314467 -16819 314853 -16753
rect 317811 -16819 318197 -16753
rect 321155 -16819 321541 -16753
rect 324499 -16819 324885 -16753
rect 327843 -16819 328229 -16753
rect 331187 -16819 331573 -16753
rect 334531 -16819 334917 -16753
rect 337875 -16819 338261 -16753
rect 341219 -16819 341605 -16753
rect 344563 -16819 344949 -16753
rect 347907 -16819 348293 -16753
rect 351251 -16819 351637 -16753
rect 354595 -16819 354981 -16753
rect 357939 -16819 358325 -16753
rect 361283 -16819 361669 -16753
rect 364627 -16819 365013 -16753
rect 367971 -16819 368357 -16753
rect 371315 -16819 371701 -16753
rect 374659 -16819 375045 -16753
rect 378003 -16819 378389 -16753
rect 381347 -16819 381733 -16753
rect 384691 -16819 385077 -16753
rect 388035 -16819 388421 -16753
rect 391379 -16819 391765 -16753
rect 394723 -16819 395109 -16753
rect 398067 -16819 398453 -16753
rect 401411 -16819 401797 -16753
rect 404755 -16819 405141 -16753
rect 408099 -16819 408485 -16753
rect 411443 -16819 411829 -16753
rect 414787 -16819 415173 -16753
rect 418131 -16819 418517 -16753
rect 421475 -16819 421861 -16753
rect 424819 -16819 425205 -16753
rect 213533 -16860 213568 -16826
rect 213882 -16832 213893 -16819
rect 213816 -16874 213893 -16832
rect 213945 -16874 214533 -16819
rect 217227 -16832 217237 -16819
rect 213816 -16877 214533 -16874
rect 213533 -16928 213568 -16894
rect 213736 -16942 213771 -16908
rect 213781 -16942 213782 -16900
rect 213617 -16991 213618 -16980
rect 213628 -17025 213663 -16991
rect 213736 -17042 213771 -17008
rect 213781 -17042 213782 -16997
rect 213629 -17078 213664 -17044
rect 213701 -17078 213736 -17044
rect 213773 -17078 213808 -17044
rect 212775 -17131 212810 -17097
rect 212871 -17131 212906 -17097
rect 212967 -17131 213002 -17097
rect 213063 -17131 213098 -17097
rect 213159 -17131 213194 -17097
rect 213816 -17114 213961 -16877
rect 214147 -16899 214533 -16877
rect 214071 -16985 214533 -16899
rect 217161 -16874 217237 -16832
rect 217289 -16874 217877 -16819
rect 220571 -16832 220581 -16819
rect 217161 -16877 217877 -16874
rect 214074 -16993 214275 -16985
rect 214090 -17003 214259 -16993
rect 213816 -17140 213991 -17114
rect 213323 -17174 213358 -17140
rect 213419 -17174 213454 -17140
rect 213515 -17174 213550 -17140
rect 213611 -17174 213646 -17140
rect 213707 -17174 213742 -17140
rect 213803 -17174 213991 -17140
rect 213816 -17200 213991 -17174
rect 214016 -17174 214117 -17050
rect 213894 -17870 213929 -17200
rect 214016 -17228 214019 -17174
rect 213701 -17936 213846 -17924
rect 213369 -17970 213846 -17936
rect 213701 -17971 213846 -17970
rect 213882 -17971 213929 -17870
rect 214028 -17971 214063 -17174
rect 214286 -17971 214321 -17062
rect 214420 -17971 214455 -16985
rect 217161 -17114 217305 -16877
rect 217491 -16899 217877 -16877
rect 217415 -16985 217877 -16899
rect 220505 -16874 220581 -16832
rect 220633 -16874 221221 -16819
rect 223915 -16832 223925 -16819
rect 220505 -16877 221221 -16874
rect 217419 -16993 217619 -16985
rect 217435 -16997 217603 -16993
rect 217161 -17200 217335 -17114
rect 217361 -17174 217461 -17050
rect 220505 -17114 220649 -16877
rect 220835 -16899 221221 -16877
rect 220759 -16985 221221 -16899
rect 223849 -16874 223925 -16832
rect 223977 -16874 224565 -16819
rect 227259 -16832 227269 -16819
rect 223849 -16877 224565 -16874
rect 220763 -16993 220963 -16985
rect 220779 -16997 220947 -16993
rect 217361 -17228 217363 -17174
rect 220505 -17200 220679 -17114
rect 220705 -17174 220805 -17050
rect 223849 -17114 223993 -16877
rect 224179 -16899 224565 -16877
rect 224103 -16985 224565 -16899
rect 227193 -16874 227269 -16832
rect 227321 -16874 227909 -16819
rect 230603 -16832 230613 -16819
rect 227193 -16877 227909 -16874
rect 224107 -16993 224307 -16985
rect 224123 -16997 224291 -16993
rect 220705 -17228 220707 -17174
rect 223849 -17200 224023 -17114
rect 224049 -17174 224149 -17050
rect 227193 -17114 227337 -16877
rect 227523 -16899 227909 -16877
rect 227447 -16985 227909 -16899
rect 230537 -16874 230613 -16832
rect 230665 -16874 231253 -16819
rect 233947 -16832 233957 -16819
rect 230537 -16877 231253 -16874
rect 227451 -16993 227651 -16985
rect 227467 -16997 227635 -16993
rect 224049 -17228 224051 -17174
rect 227193 -17200 227367 -17114
rect 227393 -17174 227493 -17050
rect 230537 -17114 230681 -16877
rect 230867 -16899 231253 -16877
rect 230791 -16985 231253 -16899
rect 233881 -16874 233957 -16832
rect 234009 -16874 234597 -16819
rect 237291 -16832 237301 -16819
rect 233881 -16877 234597 -16874
rect 230795 -16993 230995 -16985
rect 230811 -16997 230979 -16993
rect 227393 -17228 227395 -17174
rect 230537 -17200 230711 -17114
rect 230737 -17174 230837 -17050
rect 233881 -17114 234025 -16877
rect 234211 -16899 234597 -16877
rect 234135 -16985 234597 -16899
rect 237225 -16874 237301 -16832
rect 237353 -16874 237941 -16819
rect 240635 -16832 240645 -16819
rect 237225 -16877 237941 -16874
rect 234139 -16993 234339 -16985
rect 234155 -16997 234323 -16993
rect 230737 -17228 230739 -17174
rect 233881 -17200 234055 -17114
rect 234081 -17174 234181 -17050
rect 237225 -17114 237369 -16877
rect 237555 -16899 237941 -16877
rect 237479 -16985 237941 -16899
rect 240569 -16874 240645 -16832
rect 240697 -16874 241285 -16819
rect 243979 -16832 243989 -16819
rect 240569 -16877 241285 -16874
rect 237483 -16993 237683 -16985
rect 237499 -16997 237667 -16993
rect 234081 -17228 234083 -17174
rect 237225 -17200 237399 -17114
rect 237425 -17174 237525 -17050
rect 240569 -17114 240713 -16877
rect 240899 -16899 241285 -16877
rect 240823 -16985 241285 -16899
rect 243913 -16874 243989 -16832
rect 244041 -16874 244629 -16819
rect 247323 -16832 247333 -16819
rect 243913 -16877 244629 -16874
rect 240827 -16993 241027 -16985
rect 240843 -16997 241011 -16993
rect 237425 -17228 237427 -17174
rect 240569 -17200 240743 -17114
rect 240769 -17174 240869 -17050
rect 243913 -17114 244057 -16877
rect 244243 -16899 244629 -16877
rect 244167 -16985 244629 -16899
rect 247257 -16874 247333 -16832
rect 247385 -16874 247973 -16819
rect 250667 -16832 250677 -16819
rect 247257 -16877 247973 -16874
rect 244171 -16993 244371 -16985
rect 244187 -16997 244355 -16993
rect 240769 -17228 240771 -17174
rect 243913 -17200 244087 -17114
rect 244113 -17174 244213 -17050
rect 247257 -17114 247401 -16877
rect 247587 -16899 247973 -16877
rect 247511 -16985 247973 -16899
rect 250601 -16874 250677 -16832
rect 250729 -16874 251317 -16819
rect 254011 -16832 254021 -16819
rect 250601 -16877 251317 -16874
rect 247515 -16993 247715 -16985
rect 247531 -16997 247699 -16993
rect 244113 -17228 244115 -17174
rect 247257 -17200 247431 -17114
rect 247457 -17174 247557 -17050
rect 250601 -17114 250745 -16877
rect 250931 -16899 251317 -16877
rect 250855 -16985 251317 -16899
rect 253945 -16874 254021 -16832
rect 254073 -16874 254661 -16819
rect 257355 -16832 257365 -16819
rect 253945 -16877 254661 -16874
rect 250859 -16993 251059 -16985
rect 250875 -16997 251043 -16993
rect 247457 -17228 247459 -17174
rect 250601 -17200 250775 -17114
rect 250801 -17174 250901 -17050
rect 253945 -17114 254089 -16877
rect 254275 -16899 254661 -16877
rect 254199 -16985 254661 -16899
rect 257289 -16874 257365 -16832
rect 257417 -16874 258005 -16819
rect 260699 -16832 260709 -16819
rect 257289 -16877 258005 -16874
rect 254203 -16993 254403 -16985
rect 254219 -16997 254387 -16993
rect 250801 -17228 250803 -17174
rect 253945 -17200 254119 -17114
rect 254145 -17174 254245 -17050
rect 257289 -17114 257433 -16877
rect 257619 -16899 258005 -16877
rect 257543 -16985 258005 -16899
rect 260633 -16874 260709 -16832
rect 260761 -16874 261349 -16819
rect 264043 -16832 264053 -16819
rect 260633 -16877 261349 -16874
rect 257547 -16993 257747 -16985
rect 257563 -16997 257731 -16993
rect 254145 -17228 254147 -17174
rect 257289 -17200 257463 -17114
rect 257489 -17174 257589 -17050
rect 260633 -17114 260777 -16877
rect 260963 -16899 261349 -16877
rect 260887 -16985 261349 -16899
rect 263977 -16874 264053 -16832
rect 264105 -16874 264693 -16819
rect 267387 -16832 267397 -16819
rect 263977 -16877 264693 -16874
rect 260891 -16993 261091 -16985
rect 260907 -16997 261075 -16993
rect 257489 -17228 257491 -17174
rect 260633 -17200 260807 -17114
rect 260833 -17174 260933 -17050
rect 263977 -17114 264121 -16877
rect 264307 -16899 264693 -16877
rect 264231 -16985 264693 -16899
rect 267321 -16874 267397 -16832
rect 267449 -16874 268037 -16819
rect 270731 -16832 270741 -16819
rect 267321 -16877 268037 -16874
rect 264235 -16993 264435 -16985
rect 264251 -16997 264419 -16993
rect 260833 -17228 260835 -17174
rect 263977 -17200 264151 -17114
rect 264177 -17174 264277 -17050
rect 267321 -17114 267465 -16877
rect 267651 -16899 268037 -16877
rect 267575 -16985 268037 -16899
rect 270665 -16874 270741 -16832
rect 270793 -16874 271381 -16819
rect 274075 -16832 274085 -16819
rect 270665 -16877 271381 -16874
rect 267579 -16993 267779 -16985
rect 267595 -16997 267763 -16993
rect 264177 -17228 264179 -17174
rect 267321 -17200 267495 -17114
rect 267521 -17174 267621 -17050
rect 270665 -17114 270809 -16877
rect 270995 -16899 271381 -16877
rect 270919 -16985 271381 -16899
rect 274009 -16874 274085 -16832
rect 274137 -16874 274725 -16819
rect 277419 -16832 277429 -16819
rect 274009 -16877 274725 -16874
rect 270923 -16993 271123 -16985
rect 270939 -16997 271107 -16993
rect 267521 -17228 267523 -17174
rect 270665 -17200 270839 -17114
rect 270865 -17174 270965 -17050
rect 274009 -17114 274153 -16877
rect 274339 -16899 274725 -16877
rect 274263 -16985 274725 -16899
rect 277353 -16874 277429 -16832
rect 277481 -16874 278069 -16819
rect 280763 -16832 280773 -16819
rect 277353 -16877 278069 -16874
rect 274267 -16993 274467 -16985
rect 274283 -16997 274451 -16993
rect 270865 -17228 270867 -17174
rect 274009 -17200 274183 -17114
rect 274209 -17174 274309 -17050
rect 277353 -17114 277497 -16877
rect 277683 -16899 278069 -16877
rect 277607 -16985 278069 -16899
rect 280697 -16874 280773 -16832
rect 280825 -16874 281413 -16819
rect 284107 -16832 284117 -16819
rect 280697 -16877 281413 -16874
rect 277611 -16993 277811 -16985
rect 277627 -16997 277795 -16993
rect 274209 -17228 274211 -17174
rect 277353 -17200 277527 -17114
rect 277553 -17174 277653 -17050
rect 280697 -17114 280841 -16877
rect 281027 -16899 281413 -16877
rect 280951 -16985 281413 -16899
rect 284041 -16874 284117 -16832
rect 284169 -16874 284757 -16819
rect 287451 -16832 287461 -16819
rect 284041 -16877 284757 -16874
rect 280955 -16993 281155 -16985
rect 280971 -16997 281139 -16993
rect 277553 -17228 277555 -17174
rect 280697 -17200 280871 -17114
rect 280897 -17174 280997 -17050
rect 284041 -17114 284185 -16877
rect 284371 -16899 284757 -16877
rect 284295 -16985 284757 -16899
rect 287385 -16874 287461 -16832
rect 287513 -16874 288101 -16819
rect 290795 -16832 290805 -16819
rect 287385 -16877 288101 -16874
rect 284299 -16993 284499 -16985
rect 284315 -16997 284483 -16993
rect 280897 -17228 280899 -17174
rect 284041 -17200 284215 -17114
rect 284241 -17174 284341 -17050
rect 287385 -17114 287529 -16877
rect 287715 -16899 288101 -16877
rect 287639 -16985 288101 -16899
rect 290729 -16874 290805 -16832
rect 290857 -16874 291445 -16819
rect 294139 -16832 294149 -16819
rect 290729 -16877 291445 -16874
rect 287643 -16993 287843 -16985
rect 287659 -16997 287827 -16993
rect 284241 -17228 284243 -17174
rect 287385 -17200 287559 -17114
rect 287585 -17174 287685 -17050
rect 290729 -17114 290873 -16877
rect 291059 -16899 291445 -16877
rect 290983 -16985 291445 -16899
rect 294073 -16874 294149 -16832
rect 294201 -16874 294789 -16819
rect 297483 -16832 297493 -16819
rect 294073 -16877 294789 -16874
rect 290987 -16993 291187 -16985
rect 291003 -16997 291171 -16993
rect 287585 -17228 287587 -17174
rect 290729 -17200 290903 -17114
rect 290929 -17174 291029 -17050
rect 294073 -17114 294217 -16877
rect 294403 -16899 294789 -16877
rect 294327 -16985 294789 -16899
rect 297417 -16874 297493 -16832
rect 297545 -16874 298133 -16819
rect 300827 -16832 300837 -16819
rect 297417 -16877 298133 -16874
rect 294331 -16993 294531 -16985
rect 294347 -16997 294515 -16993
rect 290929 -17228 290931 -17174
rect 294073 -17200 294247 -17114
rect 294273 -17174 294373 -17050
rect 297417 -17114 297561 -16877
rect 297747 -16899 298133 -16877
rect 297671 -16985 298133 -16899
rect 300761 -16874 300837 -16832
rect 300889 -16874 301477 -16819
rect 304171 -16832 304181 -16819
rect 300761 -16877 301477 -16874
rect 297675 -16993 297875 -16985
rect 297691 -16997 297859 -16993
rect 294273 -17228 294275 -17174
rect 297417 -17200 297591 -17114
rect 297617 -17174 297717 -17050
rect 300761 -17114 300905 -16877
rect 301091 -16899 301477 -16877
rect 301015 -16985 301477 -16899
rect 304105 -16874 304181 -16832
rect 304233 -16874 304821 -16819
rect 307515 -16832 307525 -16819
rect 304105 -16877 304821 -16874
rect 301019 -16993 301219 -16985
rect 301035 -16997 301203 -16993
rect 297617 -17228 297619 -17174
rect 300761 -17200 300935 -17114
rect 300961 -17174 301061 -17050
rect 304105 -17114 304249 -16877
rect 304435 -16899 304821 -16877
rect 304359 -16985 304821 -16899
rect 307449 -16874 307525 -16832
rect 307577 -16874 308165 -16819
rect 310859 -16832 310869 -16819
rect 307449 -16877 308165 -16874
rect 304363 -16993 304563 -16985
rect 304379 -16997 304547 -16993
rect 300961 -17228 300963 -17174
rect 304105 -17200 304279 -17114
rect 304305 -17174 304405 -17050
rect 307449 -17114 307593 -16877
rect 307779 -16899 308165 -16877
rect 307703 -16985 308165 -16899
rect 310793 -16874 310869 -16832
rect 310921 -16874 311509 -16819
rect 314203 -16832 314213 -16819
rect 310793 -16877 311509 -16874
rect 307707 -16993 307907 -16985
rect 307723 -16997 307891 -16993
rect 304305 -17228 304307 -17174
rect 307449 -17200 307623 -17114
rect 307649 -17174 307749 -17050
rect 310793 -17114 310937 -16877
rect 311123 -16899 311509 -16877
rect 311047 -16985 311509 -16899
rect 314137 -16874 314213 -16832
rect 314265 -16874 314853 -16819
rect 317547 -16832 317557 -16819
rect 314137 -16877 314853 -16874
rect 311051 -16993 311251 -16985
rect 311067 -16997 311235 -16993
rect 307649 -17228 307651 -17174
rect 310793 -17200 310967 -17114
rect 310993 -17174 311093 -17050
rect 314137 -17114 314281 -16877
rect 314467 -16899 314853 -16877
rect 314391 -16985 314853 -16899
rect 317481 -16874 317557 -16832
rect 317609 -16874 318197 -16819
rect 320891 -16832 320901 -16819
rect 317481 -16877 318197 -16874
rect 314395 -16993 314595 -16985
rect 314411 -16997 314579 -16993
rect 310993 -17228 310995 -17174
rect 314137 -17200 314311 -17114
rect 314337 -17174 314437 -17050
rect 317481 -17114 317625 -16877
rect 317811 -16899 318197 -16877
rect 317735 -16985 318197 -16899
rect 320825 -16874 320901 -16832
rect 320953 -16874 321541 -16819
rect 324235 -16832 324245 -16819
rect 320825 -16877 321541 -16874
rect 317739 -16993 317939 -16985
rect 317755 -16997 317923 -16993
rect 314337 -17228 314339 -17174
rect 317481 -17200 317655 -17114
rect 317681 -17174 317781 -17050
rect 320825 -17114 320969 -16877
rect 321155 -16899 321541 -16877
rect 321079 -16985 321541 -16899
rect 324169 -16874 324245 -16832
rect 324297 -16874 324885 -16819
rect 327579 -16832 327589 -16819
rect 324169 -16877 324885 -16874
rect 321083 -16993 321283 -16985
rect 321099 -16997 321267 -16993
rect 317681 -17228 317683 -17174
rect 320825 -17200 320999 -17114
rect 321025 -17174 321125 -17050
rect 324169 -17114 324313 -16877
rect 324499 -16899 324885 -16877
rect 324423 -16985 324885 -16899
rect 327513 -16874 327589 -16832
rect 327641 -16874 328229 -16819
rect 330923 -16832 330933 -16819
rect 327513 -16877 328229 -16874
rect 324427 -16993 324627 -16985
rect 324443 -16997 324611 -16993
rect 321025 -17228 321027 -17174
rect 324169 -17200 324343 -17114
rect 324369 -17174 324469 -17050
rect 327513 -17114 327657 -16877
rect 327843 -16899 328229 -16877
rect 327767 -16985 328229 -16899
rect 330857 -16874 330933 -16832
rect 330985 -16874 331573 -16819
rect 334267 -16832 334277 -16819
rect 330857 -16877 331573 -16874
rect 327771 -16993 327971 -16985
rect 327787 -16997 327955 -16993
rect 324369 -17228 324371 -17174
rect 327513 -17200 327687 -17114
rect 327713 -17174 327813 -17050
rect 330857 -17114 331001 -16877
rect 331187 -16899 331573 -16877
rect 331111 -16985 331573 -16899
rect 334201 -16874 334277 -16832
rect 334329 -16874 334917 -16819
rect 337611 -16832 337621 -16819
rect 334201 -16877 334917 -16874
rect 331115 -16993 331315 -16985
rect 331131 -16997 331299 -16993
rect 327713 -17228 327715 -17174
rect 330857 -17200 331031 -17114
rect 331057 -17174 331157 -17050
rect 334201 -17114 334345 -16877
rect 334531 -16899 334917 -16877
rect 334455 -16985 334917 -16899
rect 337545 -16874 337621 -16832
rect 337673 -16874 338261 -16819
rect 340955 -16832 340965 -16819
rect 337545 -16877 338261 -16874
rect 334459 -16993 334659 -16985
rect 334475 -16997 334643 -16993
rect 331057 -17228 331059 -17174
rect 334201 -17200 334375 -17114
rect 334401 -17174 334501 -17050
rect 337545 -17114 337689 -16877
rect 337875 -16899 338261 -16877
rect 337799 -16985 338261 -16899
rect 340889 -16874 340965 -16832
rect 341017 -16874 341605 -16819
rect 344299 -16832 344309 -16819
rect 340889 -16877 341605 -16874
rect 337803 -16993 338003 -16985
rect 337819 -16997 337987 -16993
rect 334401 -17228 334403 -17174
rect 337545 -17200 337719 -17114
rect 337745 -17174 337845 -17050
rect 340889 -17114 341033 -16877
rect 341219 -16899 341605 -16877
rect 341143 -16985 341605 -16899
rect 344233 -16874 344309 -16832
rect 344361 -16874 344949 -16819
rect 347643 -16832 347653 -16819
rect 344233 -16877 344949 -16874
rect 341147 -16993 341347 -16985
rect 341163 -16997 341331 -16993
rect 337745 -17228 337747 -17174
rect 340889 -17200 341063 -17114
rect 341089 -17174 341189 -17050
rect 344233 -17114 344377 -16877
rect 344563 -16899 344949 -16877
rect 344487 -16985 344949 -16899
rect 347577 -16874 347653 -16832
rect 347705 -16874 348293 -16819
rect 350987 -16832 350997 -16819
rect 347577 -16877 348293 -16874
rect 344491 -16993 344691 -16985
rect 344507 -16997 344675 -16993
rect 341089 -17228 341091 -17174
rect 344233 -17200 344407 -17114
rect 344433 -17174 344533 -17050
rect 347577 -17114 347721 -16877
rect 347907 -16899 348293 -16877
rect 347831 -16985 348293 -16899
rect 350921 -16874 350997 -16832
rect 351049 -16874 351637 -16819
rect 354331 -16832 354341 -16819
rect 350921 -16877 351637 -16874
rect 347835 -16993 348035 -16985
rect 347851 -16997 348019 -16993
rect 344433 -17228 344435 -17174
rect 347577 -17200 347751 -17114
rect 347777 -17174 347877 -17050
rect 350921 -17114 351065 -16877
rect 351251 -16899 351637 -16877
rect 351175 -16985 351637 -16899
rect 354265 -16874 354341 -16832
rect 354393 -16874 354981 -16819
rect 357675 -16832 357685 -16819
rect 354265 -16877 354981 -16874
rect 351179 -16993 351379 -16985
rect 351195 -16997 351363 -16993
rect 347777 -17228 347779 -17174
rect 350921 -17200 351095 -17114
rect 351121 -17174 351221 -17050
rect 354265 -17114 354409 -16877
rect 354595 -16899 354981 -16877
rect 354519 -16985 354981 -16899
rect 357609 -16874 357685 -16832
rect 357737 -16874 358325 -16819
rect 361019 -16832 361029 -16819
rect 357609 -16877 358325 -16874
rect 354523 -16993 354723 -16985
rect 354539 -16997 354707 -16993
rect 351121 -17228 351123 -17174
rect 354265 -17200 354439 -17114
rect 354465 -17174 354565 -17050
rect 357609 -17114 357753 -16877
rect 357939 -16899 358325 -16877
rect 357863 -16985 358325 -16899
rect 360953 -16874 361029 -16832
rect 361081 -16874 361669 -16819
rect 364363 -16832 364373 -16819
rect 360953 -16877 361669 -16874
rect 357867 -16993 358067 -16985
rect 357883 -16997 358051 -16993
rect 354465 -17228 354467 -17174
rect 357609 -17200 357783 -17114
rect 357809 -17174 357909 -17050
rect 360953 -17114 361097 -16877
rect 361283 -16899 361669 -16877
rect 361207 -16985 361669 -16899
rect 364297 -16874 364373 -16832
rect 364425 -16874 365013 -16819
rect 367707 -16832 367717 -16819
rect 364297 -16877 365013 -16874
rect 361211 -16993 361411 -16985
rect 361227 -16997 361395 -16993
rect 357809 -17228 357811 -17174
rect 360953 -17200 361127 -17114
rect 361153 -17174 361253 -17050
rect 364297 -17114 364441 -16877
rect 364627 -16899 365013 -16877
rect 364551 -16985 365013 -16899
rect 367641 -16874 367717 -16832
rect 367769 -16874 368357 -16819
rect 371051 -16832 371061 -16819
rect 367641 -16877 368357 -16874
rect 364555 -16993 364755 -16985
rect 364571 -16997 364739 -16993
rect 361153 -17228 361155 -17174
rect 364297 -17200 364471 -17114
rect 364497 -17174 364597 -17050
rect 367641 -17114 367785 -16877
rect 367971 -16899 368357 -16877
rect 367895 -16985 368357 -16899
rect 370985 -16874 371061 -16832
rect 371113 -16874 371701 -16819
rect 374395 -16832 374405 -16819
rect 370985 -16877 371701 -16874
rect 367899 -16993 368099 -16985
rect 367915 -16997 368083 -16993
rect 364497 -17228 364499 -17174
rect 367641 -17200 367815 -17114
rect 367841 -17174 367941 -17050
rect 370985 -17114 371129 -16877
rect 371315 -16899 371701 -16877
rect 371239 -16985 371701 -16899
rect 374329 -16874 374405 -16832
rect 374457 -16874 375045 -16819
rect 377739 -16832 377749 -16819
rect 374329 -16877 375045 -16874
rect 371243 -16993 371443 -16985
rect 371259 -16997 371427 -16993
rect 367841 -17228 367843 -17174
rect 370985 -17200 371159 -17114
rect 371185 -17174 371285 -17050
rect 374329 -17114 374473 -16877
rect 374659 -16899 375045 -16877
rect 374583 -16985 375045 -16899
rect 377673 -16874 377749 -16832
rect 377801 -16874 378389 -16819
rect 381083 -16832 381093 -16819
rect 377673 -16877 378389 -16874
rect 374587 -16993 374787 -16985
rect 374603 -16997 374771 -16993
rect 371185 -17228 371187 -17174
rect 374329 -17200 374503 -17114
rect 374529 -17174 374629 -17050
rect 377673 -17114 377817 -16877
rect 378003 -16899 378389 -16877
rect 377927 -16985 378389 -16899
rect 381017 -16874 381093 -16832
rect 381145 -16874 381733 -16819
rect 384427 -16832 384437 -16819
rect 381017 -16877 381733 -16874
rect 377931 -16993 378131 -16985
rect 377947 -16997 378115 -16993
rect 374529 -17228 374531 -17174
rect 377673 -17200 377847 -17114
rect 377873 -17174 377973 -17050
rect 381017 -17114 381161 -16877
rect 381347 -16899 381733 -16877
rect 381271 -16985 381733 -16899
rect 384361 -16874 384437 -16832
rect 384489 -16874 385077 -16819
rect 387771 -16832 387781 -16819
rect 384361 -16877 385077 -16874
rect 381275 -16993 381475 -16985
rect 381291 -16997 381459 -16993
rect 377873 -17228 377875 -17174
rect 381017 -17200 381191 -17114
rect 381217 -17174 381317 -17050
rect 384361 -17114 384505 -16877
rect 384691 -16899 385077 -16877
rect 384615 -16985 385077 -16899
rect 387705 -16874 387781 -16832
rect 387833 -16874 388421 -16819
rect 391115 -16832 391125 -16819
rect 387705 -16877 388421 -16874
rect 384619 -16993 384819 -16985
rect 384635 -16997 384803 -16993
rect 381217 -17228 381219 -17174
rect 384361 -17200 384535 -17114
rect 384561 -17174 384661 -17050
rect 387705 -17114 387849 -16877
rect 388035 -16899 388421 -16877
rect 387959 -16985 388421 -16899
rect 391049 -16874 391125 -16832
rect 391177 -16874 391765 -16819
rect 394459 -16832 394469 -16819
rect 391049 -16877 391765 -16874
rect 387963 -16993 388163 -16985
rect 387979 -16997 388147 -16993
rect 384561 -17228 384563 -17174
rect 387705 -17200 387879 -17114
rect 387905 -17174 388005 -17050
rect 391049 -17114 391193 -16877
rect 391379 -16899 391765 -16877
rect 391303 -16985 391765 -16899
rect 394393 -16874 394469 -16832
rect 394521 -16874 395109 -16819
rect 397803 -16832 397813 -16819
rect 394393 -16877 395109 -16874
rect 391307 -16993 391507 -16985
rect 391323 -16997 391491 -16993
rect 387905 -17228 387907 -17174
rect 391049 -17200 391223 -17114
rect 391249 -17174 391349 -17050
rect 394393 -17114 394537 -16877
rect 394723 -16899 395109 -16877
rect 394647 -16985 395109 -16899
rect 397737 -16874 397813 -16832
rect 397865 -16874 398453 -16819
rect 401147 -16832 401157 -16819
rect 397737 -16877 398453 -16874
rect 394651 -16993 394851 -16985
rect 394667 -16997 394835 -16993
rect 391249 -17228 391251 -17174
rect 394393 -17200 394567 -17114
rect 394593 -17174 394693 -17050
rect 397737 -17114 397881 -16877
rect 398067 -16899 398453 -16877
rect 397991 -16985 398453 -16899
rect 401081 -16874 401157 -16832
rect 401209 -16874 401797 -16819
rect 404491 -16832 404501 -16819
rect 401081 -16877 401797 -16874
rect 397995 -16993 398195 -16985
rect 398011 -16997 398179 -16993
rect 394593 -17228 394595 -17174
rect 397737 -17200 397911 -17114
rect 397937 -17174 398037 -17050
rect 401081 -17114 401225 -16877
rect 401411 -16899 401797 -16877
rect 401335 -16985 401797 -16899
rect 404425 -16874 404501 -16832
rect 404553 -16874 405141 -16819
rect 407835 -16832 407845 -16819
rect 404425 -16877 405141 -16874
rect 401339 -16993 401539 -16985
rect 401355 -16997 401523 -16993
rect 397937 -17228 397939 -17174
rect 401081 -17200 401255 -17114
rect 401281 -17174 401381 -17050
rect 404425 -17114 404569 -16877
rect 404755 -16899 405141 -16877
rect 404679 -16985 405141 -16899
rect 407769 -16874 407845 -16832
rect 407897 -16874 408485 -16819
rect 411179 -16832 411189 -16819
rect 407769 -16877 408485 -16874
rect 404683 -16993 404883 -16985
rect 404699 -16997 404867 -16993
rect 401281 -17228 401283 -17174
rect 404425 -17200 404599 -17114
rect 404625 -17174 404725 -17050
rect 407769 -17114 407913 -16877
rect 408099 -16899 408485 -16877
rect 408023 -16985 408485 -16899
rect 411113 -16874 411189 -16832
rect 411241 -16874 411829 -16819
rect 414523 -16832 414533 -16819
rect 411113 -16877 411829 -16874
rect 408027 -16993 408227 -16985
rect 408043 -16997 408211 -16993
rect 404625 -17228 404627 -17174
rect 407769 -17200 407943 -17114
rect 407969 -17174 408069 -17050
rect 411113 -17114 411257 -16877
rect 411443 -16899 411829 -16877
rect 411367 -16985 411829 -16899
rect 414457 -16874 414533 -16832
rect 414585 -16874 415173 -16819
rect 417867 -16832 417877 -16819
rect 414457 -16877 415173 -16874
rect 411371 -16993 411571 -16985
rect 411387 -16997 411555 -16993
rect 407969 -17228 407971 -17174
rect 411113 -17200 411287 -17114
rect 411313 -17174 411413 -17050
rect 414457 -17114 414601 -16877
rect 414787 -16899 415173 -16877
rect 414711 -16985 415173 -16899
rect 417801 -16874 417877 -16832
rect 417929 -16874 418517 -16819
rect 421211 -16832 421221 -16819
rect 417801 -16877 418517 -16874
rect 414715 -16993 414915 -16985
rect 414731 -16997 414899 -16993
rect 411313 -17228 411315 -17174
rect 414457 -17200 414631 -17114
rect 414657 -17174 414757 -17050
rect 417801 -17114 417945 -16877
rect 418131 -16899 418517 -16877
rect 418055 -16985 418517 -16899
rect 421145 -16874 421221 -16832
rect 421273 -16874 421861 -16819
rect 424555 -16832 424565 -16819
rect 421145 -16877 421861 -16874
rect 418059 -16993 418259 -16985
rect 418075 -16997 418243 -16993
rect 414657 -17228 414659 -17174
rect 417801 -17200 417975 -17114
rect 418001 -17174 418101 -17050
rect 421145 -17114 421289 -16877
rect 421475 -16899 421861 -16877
rect 421399 -16985 421861 -16899
rect 424489 -16874 424565 -16832
rect 424617 -16874 425205 -16819
rect 427899 -16832 427909 -16819
rect 424489 -16877 425205 -16874
rect 421403 -16993 421603 -16985
rect 421419 -16997 421587 -16993
rect 418001 -17228 418003 -17174
rect 421145 -17200 421319 -17114
rect 421345 -17174 421445 -17050
rect 424489 -17114 424633 -16877
rect 424819 -16899 425205 -16877
rect 424743 -16985 425205 -16899
rect 427833 -16874 427909 -16832
rect 424747 -16993 424947 -16985
rect 424763 -16997 424931 -16993
rect 421345 -17228 421347 -17174
rect 424489 -17200 424663 -17114
rect 424689 -17174 424789 -17050
rect 427833 -17114 427977 -16874
rect 424689 -17228 424691 -17174
rect 427833 -17200 428007 -17114
rect 428033 -17174 428133 -17050
rect 428033 -17228 428035 -17174
rect 217046 -17971 217190 -17924
rect 217227 -17971 217244 -17870
rect 220390 -17971 220534 -17924
rect 220571 -17971 220588 -17870
rect 223734 -17971 223878 -17924
rect 223915 -17971 223932 -17870
rect 227078 -17971 227222 -17924
rect 227259 -17971 227276 -17870
rect 230422 -17971 230566 -17924
rect 230603 -17971 230620 -17870
rect 233766 -17971 233910 -17924
rect 233947 -17971 233964 -17870
rect 237110 -17971 237254 -17924
rect 237291 -17971 237308 -17870
rect 240454 -17971 240598 -17924
rect 240635 -17971 240652 -17870
rect 243798 -17971 243942 -17924
rect 243979 -17971 243996 -17870
rect 247142 -17971 247286 -17924
rect 247323 -17971 247340 -17870
rect 250486 -17971 250630 -17924
rect 250667 -17971 250684 -17870
rect 253830 -17971 253974 -17924
rect 254011 -17971 254028 -17870
rect 257174 -17971 257318 -17924
rect 257355 -17971 257372 -17870
rect 260518 -17971 260662 -17924
rect 260699 -17971 260716 -17870
rect 263862 -17971 264006 -17924
rect 264043 -17971 264060 -17870
rect 267206 -17971 267350 -17924
rect 267387 -17971 267404 -17870
rect 270550 -17971 270694 -17924
rect 270731 -17971 270748 -17870
rect 273894 -17971 274038 -17924
rect 274075 -17971 274092 -17870
rect 277238 -17971 277382 -17924
rect 277419 -17971 277436 -17870
rect 280582 -17971 280726 -17924
rect 280763 -17971 280780 -17870
rect 283926 -17971 284070 -17924
rect 284107 -17971 284124 -17870
rect 287270 -17971 287414 -17924
rect 287451 -17971 287468 -17870
rect 290614 -17971 290758 -17924
rect 290795 -17971 290812 -17870
rect 293958 -17971 294102 -17924
rect 294139 -17971 294156 -17870
rect 297302 -17971 297446 -17924
rect 297483 -17971 297500 -17870
rect 300646 -17971 300790 -17924
rect 300827 -17971 300844 -17870
rect 303990 -17971 304134 -17924
rect 304171 -17971 304188 -17870
rect 307334 -17971 307478 -17924
rect 307515 -17971 307532 -17870
rect 310678 -17971 310822 -17924
rect 310859 -17971 310876 -17870
rect 314022 -17971 314166 -17924
rect 314203 -17971 314220 -17870
rect 317366 -17971 317510 -17924
rect 317547 -17971 317564 -17870
rect 320710 -17971 320854 -17924
rect 320891 -17971 320908 -17870
rect 324054 -17971 324198 -17924
rect 324235 -17971 324252 -17870
rect 327398 -17971 327542 -17924
rect 327579 -17971 327596 -17870
rect 330742 -17971 330886 -17924
rect 330923 -17971 330940 -17870
rect 334086 -17971 334230 -17924
rect 334267 -17971 334284 -17870
rect 337430 -17971 337574 -17924
rect 337611 -17971 337628 -17870
rect 340774 -17971 340918 -17924
rect 340955 -17971 340972 -17870
rect 344118 -17971 344262 -17924
rect 344299 -17971 344316 -17870
rect 347462 -17971 347606 -17924
rect 347643 -17971 347660 -17870
rect 350806 -17971 350950 -17924
rect 350987 -17971 351004 -17870
rect 354150 -17971 354294 -17924
rect 354331 -17971 354348 -17870
rect 357494 -17971 357638 -17924
rect 357675 -17971 357692 -17870
rect 360838 -17971 360982 -17924
rect 361019 -17971 361036 -17870
rect 364182 -17971 364326 -17924
rect 364363 -17971 364380 -17870
rect 367526 -17971 367670 -17924
rect 367707 -17971 367724 -17870
rect 370870 -17971 371014 -17924
rect 371051 -17971 371068 -17870
rect 374214 -17971 374358 -17924
rect 374395 -17971 374412 -17870
rect 377558 -17971 377702 -17924
rect 377739 -17971 377756 -17870
rect 380902 -17971 381046 -17924
rect 381083 -17971 381100 -17870
rect 384246 -17971 384390 -17924
rect 384427 -17971 384444 -17870
rect 387590 -17971 387734 -17924
rect 387771 -17971 387788 -17870
rect 390934 -17971 391078 -17924
rect 391115 -17971 391132 -17870
rect 394278 -17971 394422 -17924
rect 394459 -17971 394476 -17870
rect 397622 -17971 397766 -17924
rect 397803 -17971 397820 -17870
rect 400966 -17971 401110 -17924
rect 401147 -17971 401164 -17870
rect 404310 -17971 404454 -17924
rect 404491 -17971 404508 -17870
rect 407654 -17971 407798 -17924
rect 407835 -17971 407852 -17870
rect 410998 -17971 411142 -17924
rect 411179 -17971 411196 -17870
rect 414342 -17971 414486 -17924
rect 414523 -17971 414540 -17870
rect 417686 -17971 417830 -17924
rect 417867 -17971 417884 -17870
rect 421030 -17971 421174 -17924
rect 421211 -17971 421228 -17870
rect 424374 -17971 424518 -17924
rect 424555 -17971 424572 -17870
rect 427718 -17971 427862 -17924
rect 427899 -17971 427916 -17870
rect 39806 -17982 40586 -17971
rect 43150 -17982 43930 -17971
rect 46494 -17982 47274 -17971
rect 49838 -17982 50618 -17971
rect 53182 -17982 53962 -17971
rect 56527 -17982 57306 -17971
rect 59871 -17982 60650 -17971
rect 63215 -17982 63994 -17971
rect 66559 -17982 67338 -17971
rect 69903 -17982 70682 -17971
rect 73247 -17982 74026 -17971
rect 76591 -17982 77370 -17971
rect 79935 -17982 80714 -17971
rect 83279 -17982 84058 -17971
rect 86623 -17982 87402 -17971
rect 89967 -17982 90746 -17971
rect 93311 -17982 94090 -17971
rect 96655 -17982 97434 -17971
rect 99999 -17982 100778 -17971
rect 103343 -17982 104122 -17971
rect 106687 -17982 107466 -17971
rect 110037 -17982 110810 -17971
rect 113381 -17982 114154 -17971
rect 116725 -17982 117498 -17971
rect 120069 -17982 120842 -17971
rect 123413 -17982 124186 -17971
rect 126757 -17982 127530 -17971
rect 130101 -17982 130874 -17971
rect 133445 -17982 134218 -17971
rect 136789 -17982 137562 -17971
rect 140133 -17982 140906 -17971
rect 143477 -17982 144250 -17971
rect 146821 -17982 147594 -17971
rect 150165 -17982 150938 -17971
rect 153509 -17982 154282 -17971
rect 156853 -17982 157626 -17971
rect 160197 -17982 160970 -17971
rect 163541 -17982 164314 -17971
rect 166885 -17982 167658 -17971
rect 170229 -17982 171002 -17971
rect 173573 -17982 174346 -17971
rect 176917 -17982 177690 -17971
rect 180261 -17982 181034 -17971
rect 183605 -17982 184378 -17971
rect 186949 -17982 187722 -17971
rect 190293 -17982 191066 -17971
rect 193637 -17982 194410 -17971
rect 196981 -17982 197754 -17971
rect 200325 -17982 201098 -17971
rect 203669 -17982 204442 -17971
rect 207013 -17982 207786 -17971
rect 210357 -17982 211130 -17971
rect 213701 -17982 214474 -17971
rect 217046 -17982 217818 -17971
rect 220390 -17982 221162 -17971
rect 223734 -17982 224506 -17971
rect 227078 -17982 227850 -17971
rect 230422 -17982 231194 -17971
rect 233766 -17982 234538 -17971
rect 237110 -17982 237882 -17971
rect 240454 -17982 241226 -17971
rect 243798 -17982 244570 -17971
rect 247142 -17982 247914 -17971
rect 250486 -17982 251258 -17971
rect 253830 -17982 254602 -17971
rect 257174 -17982 257946 -17971
rect 260518 -17982 261290 -17971
rect 263862 -17982 264634 -17971
rect 267206 -17982 267978 -17971
rect 270550 -17982 271322 -17971
rect 273894 -17982 274666 -17971
rect 277238 -17982 278010 -17971
rect 280582 -17982 281354 -17971
rect 283926 -17982 284698 -17971
rect 287270 -17982 288042 -17971
rect 290614 -17982 291386 -17971
rect 293958 -17982 294730 -17971
rect 297302 -17982 298074 -17971
rect 300646 -17982 301418 -17971
rect 303990 -17982 304762 -17971
rect 307334 -17982 308106 -17971
rect 310678 -17982 311450 -17971
rect 314022 -17982 314794 -17971
rect 317366 -17982 318138 -17971
rect 320710 -17982 321482 -17971
rect 324054 -17982 324826 -17971
rect 327398 -17982 328170 -17971
rect 330742 -17982 331514 -17971
rect 334086 -17982 334858 -17971
rect 337430 -17982 338202 -17971
rect 340774 -17982 341546 -17971
rect 344118 -17982 344890 -17971
rect 347462 -17982 348234 -17971
rect 350806 -17982 351578 -17971
rect 354150 -17982 354922 -17971
rect 357494 -17982 358266 -17971
rect 360838 -17982 361610 -17971
rect 364182 -17982 364954 -17971
rect 367526 -17982 368298 -17971
rect 370870 -17982 371642 -17971
rect 374214 -17982 374986 -17971
rect 377558 -17982 378330 -17971
rect 380902 -17982 381674 -17971
rect 384246 -17982 385018 -17971
rect 387590 -17982 388362 -17971
rect 390934 -17982 391706 -17971
rect 394278 -17982 395050 -17971
rect 397622 -17982 398394 -17971
rect 400966 -17982 401738 -17971
rect 404310 -17982 405082 -17971
rect 407654 -17982 408426 -17971
rect 410998 -17982 411770 -17971
rect 414342 -17982 415114 -17971
rect 417686 -17982 418458 -17971
rect 421030 -17982 421802 -17971
rect 424374 -17982 425146 -17971
rect 427718 -17982 428490 -17971
rect 39892 -18007 40586 -17982
rect 43236 -18007 43930 -17982
rect 46580 -18007 47274 -17982
rect 49924 -18007 50618 -17982
rect 53268 -18007 53962 -17982
rect 56613 -18007 57306 -17982
rect 59957 -18007 60650 -17982
rect 63301 -18007 63994 -17982
rect 66645 -18007 67338 -17982
rect 69989 -18007 70682 -17982
rect 73333 -18007 74026 -17982
rect 76677 -18007 77370 -17982
rect 80021 -18007 80714 -17982
rect 83365 -18007 84058 -17982
rect 86709 -18007 87402 -17982
rect 90053 -18007 90746 -17982
rect 93397 -18007 94090 -17982
rect 96741 -18007 97434 -17982
rect 100085 -18007 100778 -17982
rect 103429 -18007 104122 -17982
rect 106773 -18007 107466 -17982
rect 110123 -18007 110810 -17982
rect 113467 -18007 114154 -17982
rect 116811 -18007 117498 -17982
rect 120155 -18007 120842 -17982
rect 123499 -18007 124186 -17982
rect 126843 -18007 127530 -17982
rect 130187 -18007 130874 -17982
rect 133531 -18007 134218 -17982
rect 136875 -18007 137562 -17982
rect 140219 -18007 140906 -17982
rect 143563 -18007 144250 -17982
rect 146907 -18007 147594 -17982
rect 150251 -18007 150938 -17982
rect 153595 -18007 154282 -17982
rect 156939 -18007 157626 -17982
rect 160283 -18007 160970 -17982
rect 163627 -18007 164314 -17982
rect 166971 -18007 167658 -17982
rect 170315 -18007 171002 -17982
rect 173659 -18007 174346 -17982
rect 177003 -18007 177690 -17982
rect 180347 -18007 181034 -17982
rect 183691 -18007 184378 -17982
rect 187035 -18007 187722 -17982
rect 190379 -18007 191066 -17982
rect 193723 -18007 194410 -17982
rect 197067 -18007 197754 -17982
rect 200411 -18007 201098 -17982
rect 203755 -18007 204442 -17982
rect 207099 -18007 207786 -17982
rect 210443 -18007 211130 -17982
rect 213787 -18007 214474 -17982
rect 217132 -18007 217818 -17982
rect 220476 -18007 221162 -17982
rect 223820 -18007 224506 -17982
rect 227164 -18007 227850 -17982
rect 230508 -18007 231194 -17982
rect 233852 -18007 234538 -17982
rect 237196 -18007 237882 -17982
rect 240540 -18007 241226 -17982
rect 243884 -18007 244570 -17982
rect 247228 -18007 247914 -17982
rect 250572 -18007 251258 -17982
rect 253916 -18007 254602 -17982
rect 257260 -18007 257946 -17982
rect 260604 -18007 261290 -17982
rect 263948 -18007 264634 -17982
rect 267292 -18007 267978 -17982
rect 270636 -18007 271322 -17982
rect 273980 -18007 274666 -17982
rect 277324 -18007 278010 -17982
rect 280668 -18007 281354 -17982
rect 284012 -18007 284698 -17982
rect 287356 -18007 288042 -17982
rect 290700 -18007 291386 -17982
rect 294044 -18007 294730 -17982
rect 297388 -18007 298074 -17982
rect 300732 -18007 301418 -17982
rect 304076 -18007 304762 -17982
rect 307420 -18007 308106 -17982
rect 310764 -18007 311450 -17982
rect 314108 -18007 314794 -17982
rect 317452 -18007 318138 -17982
rect 320796 -18007 321482 -17982
rect 324140 -18007 324826 -17982
rect 327484 -18007 328170 -17982
rect 330828 -18007 331514 -17982
rect 334172 -18007 334858 -17982
rect 337516 -18007 338202 -17982
rect 340860 -18007 341546 -17982
rect 344204 -18007 344890 -17982
rect 347548 -18007 348234 -17982
rect 350892 -18007 351578 -17982
rect 354236 -18007 354922 -17982
rect 357580 -18007 358266 -17982
rect 360924 -18007 361610 -17982
rect 364268 -18007 364954 -17982
rect 367612 -18007 368298 -17982
rect 370956 -18007 371642 -17982
rect 374300 -18007 374986 -17982
rect 377644 -18007 378330 -17982
rect 380988 -18007 381674 -17982
rect 384332 -18007 385018 -17982
rect 387676 -18007 388362 -17982
rect 391020 -18007 391706 -17982
rect 394364 -18007 395050 -17982
rect 397708 -18007 398394 -17982
rect 401052 -18007 401738 -17982
rect 404396 -18007 405082 -17982
rect 407740 -18007 408426 -17982
rect 411084 -18007 411770 -17982
rect 414428 -18007 415114 -17982
rect 417772 -18007 418458 -17982
rect 421116 -18007 421802 -17982
rect 424460 -18007 425146 -17982
rect 427804 -18007 428490 -17982
rect 39922 -18032 40586 -18007
rect 43266 -18032 43930 -18007
rect 46610 -18032 47274 -18007
rect 49954 -18032 50618 -18007
rect 53298 -18032 53962 -18007
rect 38274 -18183 38280 -18149
rect 38322 -18543 38328 -18285
rect 38334 -18543 38376 -18245
rect 39378 -18506 39420 -18032
rect 39904 -18036 40586 -18032
rect 39574 -18108 39750 -18074
rect 39512 -18506 39554 -18167
rect 39558 -18506 39565 -18156
rect 39759 -18167 39766 -18156
rect 39770 -18506 39812 -18167
rect 39904 -18448 40645 -18036
rect 40657 -18118 41033 -18084
rect 41118 -18180 41129 -18118
rect 40757 -18256 40933 -18222
rect 40683 -18448 40689 -18294
rect 40695 -18448 40737 -18306
rect 40741 -18448 40748 -18295
rect 40942 -18306 40949 -18295
rect 40953 -18448 40995 -18306
rect 41001 -18448 41007 -18294
rect 41075 -18448 41081 -18220
rect 41087 -18448 41129 -18180
rect 41152 -18245 41163 -18149
rect 41248 -18183 41624 -18149
rect 41152 -18448 41194 -18245
rect 41200 -18448 41206 -18285
rect 41348 -18321 41524 -18287
rect 39904 -18506 41266 -18448
rect 38424 -19781 38477 -18667
rect 39534 -18543 41266 -18506
rect 41274 -18543 41280 -18359
rect 41286 -18543 41328 -18371
rect 41332 -18543 41339 -18360
rect 41533 -18371 41540 -18360
rect 41544 -18543 41586 -18371
rect 41592 -18543 41598 -18359
rect 41666 -18543 41672 -18285
rect 41678 -18543 41720 -18245
rect 42722 -18506 42764 -18032
rect 43248 -18036 43930 -18032
rect 42918 -18108 43094 -18074
rect 42856 -18506 42898 -18167
rect 42902 -18506 42909 -18156
rect 43103 -18167 43110 -18156
rect 43114 -18506 43156 -18167
rect 43248 -18448 43989 -18036
rect 44001 -18118 44377 -18084
rect 44462 -18180 44473 -18118
rect 44101 -18256 44277 -18222
rect 44027 -18448 44033 -18294
rect 44039 -18448 44081 -18306
rect 44085 -18448 44092 -18295
rect 44286 -18306 44293 -18295
rect 44297 -18448 44339 -18306
rect 44345 -18448 44351 -18294
rect 44419 -18448 44425 -18220
rect 44431 -18448 44473 -18180
rect 44496 -18245 44507 -18149
rect 44592 -18183 44968 -18149
rect 44496 -18448 44538 -18245
rect 44544 -18448 44550 -18285
rect 44692 -18321 44868 -18287
rect 43248 -18506 44610 -18448
rect 42675 -18543 44610 -18506
rect 44618 -18543 44624 -18359
rect 44630 -18543 44672 -18371
rect 44676 -18543 44683 -18360
rect 44877 -18371 44884 -18360
rect 44888 -18543 44930 -18371
rect 44936 -18543 44942 -18359
rect 45010 -18543 45016 -18285
rect 45022 -18543 45064 -18245
rect 46066 -18506 46108 -18032
rect 46592 -18036 47274 -18032
rect 46262 -18108 46438 -18074
rect 46200 -18506 46242 -18167
rect 46246 -18506 46253 -18156
rect 46447 -18167 46454 -18156
rect 46458 -18506 46500 -18167
rect 46592 -18448 47333 -18036
rect 47345 -18118 47721 -18084
rect 47806 -18180 47817 -18118
rect 47445 -18256 47621 -18222
rect 47371 -18448 47377 -18294
rect 47383 -18448 47425 -18306
rect 47429 -18448 47436 -18295
rect 47630 -18306 47637 -18295
rect 47641 -18448 47683 -18306
rect 47689 -18448 47695 -18294
rect 47763 -18448 47769 -18220
rect 47775 -18448 47817 -18180
rect 47840 -18245 47851 -18149
rect 47936 -18183 48312 -18149
rect 47840 -18448 47882 -18245
rect 47888 -18448 47894 -18285
rect 48036 -18321 48212 -18287
rect 46592 -18506 47954 -18448
rect 46019 -18543 47954 -18506
rect 47962 -18543 47968 -18359
rect 47974 -18543 48016 -18371
rect 48020 -18543 48027 -18360
rect 48221 -18371 48228 -18360
rect 48232 -18543 48274 -18371
rect 48280 -18543 48286 -18359
rect 48354 -18543 48360 -18285
rect 48366 -18543 48408 -18245
rect 49410 -18506 49452 -18032
rect 49936 -18036 50618 -18032
rect 49606 -18108 49782 -18074
rect 49544 -18506 49586 -18167
rect 49590 -18506 49597 -18156
rect 49791 -18167 49798 -18156
rect 49802 -18506 49844 -18167
rect 49936 -18448 50677 -18036
rect 50689 -18118 51065 -18084
rect 51150 -18180 51161 -18118
rect 50789 -18256 50965 -18222
rect 50715 -18448 50721 -18294
rect 50727 -18448 50769 -18306
rect 50773 -18448 50780 -18295
rect 50974 -18306 50981 -18295
rect 50985 -18448 51027 -18306
rect 51033 -18448 51039 -18294
rect 51107 -18448 51113 -18220
rect 51119 -18448 51161 -18180
rect 51184 -18245 51195 -18149
rect 51280 -18183 51656 -18149
rect 51184 -18448 51226 -18245
rect 51232 -18448 51238 -18285
rect 51380 -18321 51556 -18287
rect 49936 -18506 51298 -18448
rect 49363 -18543 51298 -18506
rect 51306 -18543 51312 -18359
rect 51318 -18543 51360 -18371
rect 51364 -18543 51371 -18360
rect 51565 -18371 51572 -18360
rect 51576 -18543 51618 -18371
rect 51624 -18543 51630 -18359
rect 51698 -18543 51704 -18285
rect 51710 -18543 51752 -18245
rect 52754 -18506 52796 -18032
rect 53280 -18036 53962 -18032
rect 52950 -18108 53126 -18074
rect 52888 -18506 52930 -18167
rect 52934 -18506 52941 -18156
rect 53135 -18167 53142 -18156
rect 53146 -18506 53188 -18167
rect 53280 -18448 54021 -18036
rect 54033 -18118 54409 -18084
rect 54494 -18180 54505 -18118
rect 54133 -18256 54309 -18222
rect 54059 -18448 54065 -18294
rect 54071 -18448 54113 -18306
rect 54117 -18448 54124 -18295
rect 54318 -18306 54325 -18295
rect 54329 -18448 54371 -18306
rect 54377 -18448 54383 -18294
rect 54451 -18448 54457 -18220
rect 54463 -18448 54505 -18180
rect 54528 -18245 54539 -18149
rect 54624 -18183 55000 -18149
rect 54528 -18448 54570 -18245
rect 54576 -18448 54582 -18285
rect 54724 -18321 54900 -18287
rect 53280 -18506 54642 -18448
rect 52707 -18543 54642 -18506
rect 54650 -18543 54656 -18359
rect 54662 -18543 54704 -18371
rect 54708 -18543 54715 -18360
rect 54909 -18371 54916 -18360
rect 54920 -18543 54962 -18371
rect 54968 -18543 54974 -18359
rect 55042 -18543 55048 -18285
rect 55054 -18543 55096 -18245
rect 56099 -18506 56140 -18032
rect 56625 -18036 57306 -18007
rect 56295 -18108 56470 -18074
rect 56233 -18506 56274 -18167
rect 56279 -18506 56285 -18156
rect 56480 -18167 56486 -18156
rect 56491 -18506 56532 -18167
rect 56625 -18448 57365 -18036
rect 57378 -18118 57753 -18084
rect 57839 -18180 57849 -18118
rect 57478 -18256 57653 -18222
rect 57404 -18448 57409 -18294
rect 57416 -18448 57457 -18306
rect 57462 -18448 57468 -18295
rect 57663 -18306 57669 -18295
rect 57674 -18448 57715 -18306
rect 57722 -18448 57727 -18294
rect 57796 -18448 57801 -18220
rect 57808 -18448 57849 -18180
rect 57873 -18245 57883 -18149
rect 57969 -18183 58344 -18149
rect 57873 -18448 57914 -18245
rect 57921 -18448 57926 -18285
rect 58069 -18321 58244 -18287
rect 56625 -18506 57986 -18448
rect 56052 -18543 57986 -18506
rect 57995 -18543 58000 -18359
rect 58007 -18543 58048 -18371
rect 58053 -18543 58059 -18360
rect 58254 -18371 58260 -18360
rect 58265 -18543 58306 -18371
rect 58313 -18543 58318 -18359
rect 58387 -18543 58392 -18285
rect 58399 -18543 58440 -18245
rect 59443 -18506 59484 -18032
rect 59969 -18036 60650 -18007
rect 59639 -18108 59814 -18074
rect 59577 -18506 59618 -18167
rect 59623 -18506 59629 -18156
rect 59824 -18167 59830 -18156
rect 59835 -18506 59876 -18167
rect 59969 -18448 60709 -18036
rect 60722 -18118 61097 -18084
rect 61183 -18180 61193 -18118
rect 60822 -18256 60997 -18222
rect 60748 -18448 60753 -18294
rect 60760 -18448 60801 -18306
rect 60806 -18448 60812 -18295
rect 61007 -18306 61013 -18295
rect 61018 -18448 61059 -18306
rect 61066 -18448 61071 -18294
rect 61140 -18448 61145 -18220
rect 61152 -18448 61193 -18180
rect 61217 -18245 61227 -18149
rect 61313 -18183 61688 -18149
rect 61217 -18448 61258 -18245
rect 61265 -18448 61270 -18285
rect 61413 -18321 61588 -18287
rect 59969 -18506 61330 -18448
rect 59396 -18543 61330 -18506
rect 61339 -18543 61344 -18359
rect 61351 -18543 61392 -18371
rect 61397 -18543 61403 -18360
rect 61598 -18371 61604 -18360
rect 61609 -18543 61650 -18371
rect 61657 -18543 61662 -18359
rect 61731 -18543 61736 -18285
rect 61743 -18543 61784 -18245
rect 62787 -18506 62828 -18032
rect 63313 -18036 63994 -18007
rect 62983 -18108 63158 -18074
rect 62921 -18506 62962 -18167
rect 62967 -18506 62973 -18156
rect 63168 -18167 63174 -18156
rect 63179 -18506 63220 -18167
rect 63313 -18448 64053 -18036
rect 64066 -18118 64441 -18084
rect 64527 -18180 64537 -18118
rect 64166 -18256 64341 -18222
rect 64092 -18448 64097 -18294
rect 64104 -18448 64145 -18306
rect 64150 -18448 64156 -18295
rect 64351 -18306 64357 -18295
rect 64362 -18448 64403 -18306
rect 64410 -18448 64415 -18294
rect 64484 -18448 64489 -18220
rect 64496 -18448 64537 -18180
rect 64561 -18245 64571 -18149
rect 64657 -18183 65032 -18149
rect 64561 -18448 64602 -18245
rect 64609 -18448 64614 -18285
rect 64757 -18321 64932 -18287
rect 63313 -18506 64674 -18448
rect 62740 -18543 64674 -18506
rect 64683 -18543 64688 -18359
rect 64695 -18543 64736 -18371
rect 64741 -18543 64747 -18360
rect 64942 -18371 64948 -18360
rect 64953 -18543 64994 -18371
rect 65001 -18543 65006 -18359
rect 65075 -18543 65080 -18285
rect 65087 -18543 65128 -18245
rect 66131 -18506 66172 -18032
rect 66657 -18036 67338 -18007
rect 66327 -18108 66502 -18074
rect 66265 -18506 66306 -18167
rect 66311 -18506 66317 -18156
rect 66512 -18167 66518 -18156
rect 66523 -18506 66564 -18167
rect 66657 -18448 67397 -18036
rect 67410 -18118 67785 -18084
rect 67871 -18180 67881 -18118
rect 67510 -18256 67685 -18222
rect 67436 -18448 67441 -18294
rect 67448 -18448 67489 -18306
rect 67494 -18448 67500 -18295
rect 67695 -18306 67701 -18295
rect 67706 -18448 67747 -18306
rect 67754 -18448 67759 -18294
rect 67828 -18448 67833 -18220
rect 67840 -18448 67881 -18180
rect 67905 -18245 67915 -18149
rect 68001 -18183 68376 -18149
rect 67905 -18448 67946 -18245
rect 67953 -18448 67958 -18285
rect 68101 -18321 68276 -18287
rect 66657 -18506 68018 -18448
rect 66084 -18543 68018 -18506
rect 68027 -18543 68032 -18359
rect 68039 -18543 68080 -18371
rect 68085 -18543 68091 -18360
rect 68286 -18371 68292 -18360
rect 68297 -18543 68338 -18371
rect 68345 -18543 68350 -18359
rect 68419 -18543 68424 -18285
rect 68431 -18543 68472 -18245
rect 69475 -18506 69516 -18032
rect 70001 -18036 70682 -18007
rect 69671 -18108 69846 -18074
rect 69609 -18506 69650 -18167
rect 69655 -18506 69661 -18156
rect 69856 -18167 69862 -18156
rect 69867 -18506 69908 -18167
rect 70001 -18448 70741 -18036
rect 70754 -18118 71129 -18084
rect 71215 -18180 71225 -18118
rect 70854 -18256 71029 -18222
rect 70780 -18448 70785 -18294
rect 70792 -18448 70833 -18306
rect 70838 -18448 70844 -18295
rect 71039 -18306 71045 -18295
rect 71050 -18448 71091 -18306
rect 71098 -18448 71103 -18294
rect 71172 -18448 71177 -18220
rect 71184 -18448 71225 -18180
rect 71249 -18245 71259 -18149
rect 71345 -18183 71720 -18149
rect 71249 -18448 71290 -18245
rect 71297 -18448 71302 -18285
rect 71445 -18321 71620 -18287
rect 70001 -18506 71362 -18448
rect 69428 -18543 71362 -18506
rect 71371 -18543 71376 -18359
rect 71383 -18543 71424 -18371
rect 71429 -18543 71435 -18360
rect 71630 -18371 71636 -18360
rect 71641 -18543 71682 -18371
rect 71689 -18543 71694 -18359
rect 71763 -18543 71768 -18285
rect 71775 -18543 71816 -18245
rect 72819 -18506 72860 -18032
rect 73345 -18036 74026 -18007
rect 73015 -18108 73190 -18074
rect 72953 -18506 72994 -18167
rect 72999 -18506 73005 -18156
rect 73200 -18167 73206 -18156
rect 73211 -18506 73252 -18167
rect 73345 -18448 74085 -18036
rect 74098 -18118 74473 -18084
rect 74559 -18180 74569 -18118
rect 74198 -18256 74373 -18222
rect 74124 -18448 74129 -18294
rect 74136 -18448 74177 -18306
rect 74182 -18448 74188 -18295
rect 74383 -18306 74389 -18295
rect 74394 -18448 74435 -18306
rect 74442 -18448 74447 -18294
rect 74516 -18448 74521 -18220
rect 74528 -18448 74569 -18180
rect 74593 -18245 74603 -18149
rect 74689 -18183 75064 -18149
rect 74593 -18448 74634 -18245
rect 74641 -18448 74646 -18285
rect 74789 -18321 74964 -18287
rect 73345 -18506 74706 -18448
rect 72772 -18543 74706 -18506
rect 74715 -18543 74720 -18359
rect 74727 -18543 74768 -18371
rect 74773 -18543 74779 -18360
rect 74974 -18371 74980 -18360
rect 74985 -18543 75026 -18371
rect 75033 -18543 75038 -18359
rect 75107 -18543 75112 -18285
rect 75119 -18543 75160 -18245
rect 76163 -18506 76204 -18032
rect 76689 -18036 77370 -18007
rect 76359 -18108 76534 -18074
rect 76297 -18506 76338 -18167
rect 76343 -18506 76349 -18156
rect 76544 -18167 76550 -18156
rect 76555 -18506 76596 -18167
rect 76689 -18448 77429 -18036
rect 77442 -18118 77817 -18084
rect 77903 -18180 77913 -18118
rect 77542 -18256 77717 -18222
rect 77468 -18448 77473 -18294
rect 77480 -18448 77521 -18306
rect 77526 -18448 77532 -18295
rect 77727 -18306 77733 -18295
rect 77738 -18448 77779 -18306
rect 77786 -18448 77791 -18294
rect 77860 -18448 77865 -18220
rect 77872 -18448 77913 -18180
rect 77937 -18245 77947 -18149
rect 78033 -18183 78408 -18149
rect 77937 -18448 77978 -18245
rect 77985 -18448 77990 -18285
rect 78133 -18321 78308 -18287
rect 76689 -18506 78050 -18448
rect 76116 -18543 78050 -18506
rect 78059 -18543 78064 -18359
rect 78071 -18543 78112 -18371
rect 78117 -18543 78123 -18360
rect 78318 -18371 78324 -18360
rect 78329 -18543 78370 -18371
rect 78377 -18543 78382 -18359
rect 78451 -18543 78456 -18285
rect 78463 -18543 78504 -18245
rect 79507 -18506 79548 -18032
rect 80033 -18036 80714 -18007
rect 79703 -18108 79878 -18074
rect 79641 -18506 79682 -18167
rect 79687 -18506 79693 -18156
rect 79888 -18167 79894 -18156
rect 79899 -18506 79940 -18167
rect 80033 -18448 80773 -18036
rect 80786 -18118 81161 -18084
rect 81247 -18180 81257 -18118
rect 80886 -18256 81061 -18222
rect 80812 -18448 80817 -18294
rect 80824 -18448 80865 -18306
rect 80870 -18448 80876 -18295
rect 81071 -18306 81077 -18295
rect 81082 -18448 81123 -18306
rect 81130 -18448 81135 -18294
rect 81204 -18448 81209 -18220
rect 81216 -18448 81257 -18180
rect 81281 -18245 81291 -18149
rect 81377 -18183 81752 -18149
rect 81281 -18448 81322 -18245
rect 81329 -18448 81334 -18285
rect 81477 -18321 81652 -18287
rect 80033 -18506 81394 -18448
rect 79460 -18543 81394 -18506
rect 81403 -18543 81408 -18359
rect 81415 -18543 81456 -18371
rect 81461 -18543 81467 -18360
rect 81662 -18371 81668 -18360
rect 81673 -18543 81714 -18371
rect 81721 -18543 81726 -18359
rect 81795 -18543 81800 -18285
rect 81807 -18543 81848 -18245
rect 82851 -18506 82892 -18032
rect 83377 -18036 84058 -18007
rect 83047 -18108 83222 -18074
rect 82985 -18506 83026 -18167
rect 83031 -18506 83037 -18156
rect 83232 -18167 83238 -18156
rect 83243 -18506 83284 -18167
rect 83377 -18448 84117 -18036
rect 84130 -18118 84505 -18084
rect 84591 -18180 84601 -18118
rect 84230 -18256 84405 -18222
rect 84156 -18448 84161 -18294
rect 84168 -18448 84209 -18306
rect 84214 -18448 84220 -18295
rect 84415 -18306 84421 -18295
rect 84426 -18448 84467 -18306
rect 84474 -18448 84479 -18294
rect 84548 -18448 84553 -18220
rect 84560 -18448 84601 -18180
rect 84625 -18245 84635 -18149
rect 84721 -18183 85096 -18149
rect 84625 -18448 84666 -18245
rect 84673 -18448 84678 -18285
rect 84821 -18321 84996 -18287
rect 83377 -18506 84738 -18448
rect 82804 -18543 84738 -18506
rect 84747 -18543 84752 -18359
rect 84759 -18543 84800 -18371
rect 84805 -18543 84811 -18360
rect 85006 -18371 85012 -18360
rect 85017 -18543 85058 -18371
rect 85065 -18543 85070 -18359
rect 85139 -18543 85144 -18285
rect 85151 -18543 85192 -18245
rect 86195 -18506 86236 -18032
rect 86721 -18036 87402 -18007
rect 86391 -18108 86566 -18074
rect 86329 -18506 86370 -18167
rect 86375 -18506 86381 -18156
rect 86576 -18167 86582 -18156
rect 86587 -18506 86628 -18167
rect 86721 -18448 87461 -18036
rect 87474 -18118 87849 -18084
rect 87935 -18180 87945 -18118
rect 87574 -18256 87749 -18222
rect 87500 -18448 87505 -18294
rect 87512 -18448 87553 -18306
rect 87558 -18448 87564 -18295
rect 87759 -18306 87765 -18295
rect 87770 -18448 87811 -18306
rect 87818 -18448 87823 -18294
rect 87892 -18448 87897 -18220
rect 87904 -18448 87945 -18180
rect 87969 -18245 87979 -18149
rect 88065 -18183 88440 -18149
rect 87969 -18448 88010 -18245
rect 88017 -18448 88022 -18285
rect 88165 -18321 88340 -18287
rect 86721 -18506 88082 -18448
rect 86148 -18543 88082 -18506
rect 88091 -18543 88096 -18359
rect 88103 -18543 88144 -18371
rect 88149 -18543 88155 -18360
rect 88350 -18371 88356 -18360
rect 88361 -18543 88402 -18371
rect 88409 -18543 88414 -18359
rect 88483 -18543 88488 -18285
rect 88495 -18543 88536 -18245
rect 89539 -18506 89580 -18032
rect 90065 -18036 90746 -18007
rect 89735 -18108 89910 -18074
rect 89673 -18506 89714 -18167
rect 89719 -18506 89725 -18156
rect 89920 -18167 89926 -18156
rect 89931 -18506 89972 -18167
rect 90065 -18448 90805 -18036
rect 90818 -18118 91193 -18084
rect 91279 -18180 91289 -18118
rect 90918 -18256 91093 -18222
rect 90844 -18448 90849 -18294
rect 90856 -18448 90897 -18306
rect 90902 -18448 90908 -18295
rect 91103 -18306 91109 -18295
rect 91114 -18448 91155 -18306
rect 91162 -18448 91167 -18294
rect 91236 -18448 91241 -18220
rect 91248 -18448 91289 -18180
rect 91313 -18245 91323 -18149
rect 91409 -18183 91784 -18149
rect 91313 -18448 91354 -18245
rect 91361 -18448 91366 -18285
rect 91509 -18321 91684 -18287
rect 90065 -18506 91426 -18448
rect 89492 -18543 91426 -18506
rect 91435 -18543 91440 -18359
rect 91447 -18543 91488 -18371
rect 91493 -18543 91499 -18360
rect 91694 -18371 91700 -18360
rect 91705 -18543 91746 -18371
rect 91753 -18543 91758 -18359
rect 91827 -18543 91832 -18285
rect 91839 -18543 91880 -18245
rect 92883 -18506 92924 -18032
rect 93409 -18036 94090 -18007
rect 93079 -18108 93254 -18074
rect 93017 -18506 93058 -18167
rect 93063 -18506 93069 -18156
rect 93264 -18167 93270 -18156
rect 93275 -18506 93316 -18167
rect 93409 -18448 94149 -18036
rect 94162 -18118 94537 -18084
rect 94623 -18180 94633 -18118
rect 94262 -18256 94437 -18222
rect 94188 -18448 94193 -18294
rect 94200 -18448 94241 -18306
rect 94246 -18448 94252 -18295
rect 94447 -18306 94453 -18295
rect 94458 -18448 94499 -18306
rect 94506 -18448 94511 -18294
rect 94580 -18448 94585 -18220
rect 94592 -18448 94633 -18180
rect 94657 -18245 94667 -18149
rect 94753 -18183 95128 -18149
rect 94657 -18448 94698 -18245
rect 94705 -18448 94710 -18285
rect 94853 -18321 95028 -18287
rect 93409 -18506 94770 -18448
rect 92836 -18543 94770 -18506
rect 94779 -18543 94784 -18359
rect 94791 -18543 94832 -18371
rect 94837 -18543 94843 -18360
rect 95038 -18371 95044 -18360
rect 95049 -18543 95090 -18371
rect 95097 -18543 95102 -18359
rect 95171 -18543 95176 -18285
rect 95183 -18543 95224 -18245
rect 96227 -18506 96268 -18032
rect 96753 -18036 97434 -18007
rect 96423 -18108 96598 -18074
rect 96361 -18506 96402 -18167
rect 96407 -18506 96413 -18156
rect 96608 -18167 96614 -18156
rect 96619 -18506 96660 -18167
rect 96753 -18448 97493 -18036
rect 97506 -18118 97881 -18084
rect 97967 -18180 97977 -18118
rect 97606 -18256 97781 -18222
rect 97532 -18448 97537 -18294
rect 97544 -18448 97585 -18306
rect 97590 -18448 97596 -18295
rect 97791 -18306 97797 -18295
rect 97802 -18448 97843 -18306
rect 97850 -18448 97855 -18294
rect 97924 -18448 97929 -18220
rect 97936 -18448 97977 -18180
rect 98001 -18245 98011 -18149
rect 98097 -18183 98472 -18149
rect 98001 -18448 98042 -18245
rect 98049 -18448 98054 -18285
rect 98197 -18321 98372 -18287
rect 96753 -18506 98114 -18448
rect 96180 -18543 98114 -18506
rect 98123 -18543 98128 -18359
rect 98135 -18543 98176 -18371
rect 98181 -18543 98187 -18360
rect 98382 -18371 98388 -18360
rect 98393 -18543 98434 -18371
rect 98441 -18543 98446 -18359
rect 98515 -18543 98520 -18285
rect 98527 -18543 98568 -18245
rect 99571 -18506 99612 -18032
rect 100097 -18036 100778 -18007
rect 99767 -18108 99942 -18074
rect 99705 -18506 99746 -18167
rect 99751 -18506 99757 -18156
rect 99952 -18167 99958 -18156
rect 99963 -18506 100004 -18167
rect 100097 -18448 100837 -18036
rect 100850 -18118 101225 -18084
rect 101311 -18180 101321 -18118
rect 100950 -18256 101125 -18222
rect 100876 -18448 100881 -18294
rect 100888 -18448 100929 -18306
rect 100934 -18448 100940 -18295
rect 101135 -18306 101141 -18295
rect 101146 -18448 101187 -18306
rect 101194 -18448 101199 -18294
rect 101268 -18448 101273 -18220
rect 101280 -18448 101321 -18180
rect 101345 -18245 101355 -18149
rect 101441 -18183 101816 -18149
rect 101345 -18448 101386 -18245
rect 101393 -18448 101398 -18285
rect 101541 -18321 101716 -18287
rect 100097 -18506 101458 -18448
rect 99524 -18543 101458 -18506
rect 101467 -18543 101472 -18359
rect 101479 -18543 101520 -18371
rect 101525 -18543 101531 -18360
rect 101726 -18371 101732 -18360
rect 101737 -18543 101778 -18371
rect 101785 -18543 101790 -18359
rect 101859 -18543 101864 -18285
rect 101871 -18543 101912 -18245
rect 102915 -18506 102956 -18032
rect 103441 -18036 104122 -18007
rect 103111 -18108 103286 -18074
rect 103049 -18506 103090 -18167
rect 103095 -18506 103101 -18156
rect 103296 -18167 103302 -18156
rect 103307 -18506 103348 -18167
rect 103441 -18448 104181 -18036
rect 104194 -18118 104569 -18084
rect 104655 -18180 104665 -18118
rect 104294 -18256 104469 -18222
rect 104220 -18448 104225 -18294
rect 104232 -18448 104273 -18306
rect 104278 -18448 104284 -18295
rect 104479 -18306 104485 -18295
rect 104490 -18448 104531 -18306
rect 104538 -18448 104543 -18294
rect 104612 -18448 104617 -18220
rect 104624 -18448 104665 -18180
rect 104689 -18245 104699 -18149
rect 104785 -18183 105160 -18149
rect 104689 -18448 104730 -18245
rect 104737 -18448 104742 -18285
rect 104885 -18321 105060 -18287
rect 103441 -18506 104802 -18448
rect 102868 -18543 104802 -18506
rect 104811 -18543 104816 -18359
rect 104823 -18543 104864 -18371
rect 104869 -18543 104875 -18360
rect 105070 -18371 105076 -18360
rect 105081 -18543 105122 -18371
rect 105129 -18543 105134 -18359
rect 105203 -18543 105208 -18285
rect 105215 -18543 105256 -18245
rect 106259 -18506 106300 -18032
rect 106785 -18036 107466 -18007
rect 106455 -18108 106630 -18074
rect 106393 -18506 106434 -18167
rect 106439 -18506 106445 -18156
rect 106640 -18167 106646 -18156
rect 106651 -18506 106692 -18167
rect 106785 -18448 107525 -18036
rect 107538 -18118 107913 -18084
rect 107999 -18180 108009 -18118
rect 107638 -18256 107813 -18222
rect 107564 -18448 107569 -18294
rect 107576 -18448 107617 -18306
rect 107622 -18448 107628 -18295
rect 107823 -18306 107829 -18295
rect 107834 -18448 107875 -18306
rect 107882 -18448 107887 -18294
rect 107956 -18448 107961 -18220
rect 107968 -18448 108009 -18180
rect 108033 -18245 108043 -18149
rect 108129 -18183 108504 -18149
rect 108033 -18448 108074 -18245
rect 108081 -18448 108086 -18285
rect 108229 -18321 108404 -18287
rect 106785 -18506 108146 -18448
rect 106212 -18543 108146 -18506
rect 108155 -18543 108160 -18359
rect 108167 -18543 108208 -18371
rect 108213 -18543 108219 -18360
rect 108414 -18371 108420 -18360
rect 108425 -18543 108466 -18371
rect 108473 -18543 108478 -18359
rect 108547 -18543 108552 -18285
rect 108559 -18543 108600 -18245
rect 109609 -18506 109644 -18032
rect 110135 -18036 110810 -18007
rect 109805 -18108 109974 -18074
rect 109743 -18506 109778 -18167
rect 110001 -18506 110036 -18167
rect 110135 -18448 110869 -18036
rect 110888 -18118 111257 -18084
rect 110988 -18256 111157 -18222
rect 110926 -18448 110961 -18306
rect 111184 -18448 111219 -18306
rect 111317 -18448 111365 -18083
rect 111371 -18448 111419 -18137
rect 111479 -18183 111848 -18149
rect 111579 -18321 111748 -18287
rect 110135 -18506 111490 -18448
rect 109562 -18543 111490 -18506
rect 111517 -18543 111552 -18371
rect 111775 -18543 111810 -18371
rect 111909 -18543 111944 -18245
rect 112953 -18506 112988 -18032
rect 113479 -18036 114154 -18007
rect 113149 -18108 113318 -18074
rect 113087 -18506 113122 -18167
rect 113345 -18506 113380 -18167
rect 113479 -18448 114213 -18036
rect 114232 -18118 114601 -18084
rect 114332 -18256 114501 -18222
rect 114270 -18448 114305 -18306
rect 114528 -18448 114563 -18306
rect 114661 -18448 114709 -18083
rect 114715 -18448 114763 -18137
rect 114823 -18183 115192 -18149
rect 114923 -18321 115092 -18287
rect 113479 -18506 114834 -18448
rect 112906 -18543 114834 -18506
rect 114861 -18543 114896 -18371
rect 115119 -18543 115154 -18371
rect 115253 -18543 115288 -18245
rect 116297 -18506 116332 -18032
rect 116823 -18036 117498 -18007
rect 116493 -18108 116662 -18074
rect 116431 -18506 116466 -18167
rect 116689 -18506 116724 -18167
rect 116823 -18448 117557 -18036
rect 117576 -18118 117945 -18084
rect 117676 -18256 117845 -18222
rect 117614 -18448 117649 -18306
rect 117872 -18448 117907 -18306
rect 118005 -18448 118053 -18083
rect 118059 -18448 118107 -18137
rect 118167 -18183 118536 -18149
rect 118267 -18321 118436 -18287
rect 116823 -18506 118178 -18448
rect 116250 -18543 118178 -18506
rect 118205 -18543 118240 -18371
rect 118463 -18543 118498 -18371
rect 118597 -18543 118632 -18245
rect 119641 -18506 119676 -18032
rect 120167 -18036 120842 -18007
rect 119837 -18108 120006 -18074
rect 119775 -18506 119810 -18167
rect 120033 -18506 120068 -18167
rect 120167 -18448 120901 -18036
rect 120920 -18118 121289 -18084
rect 121020 -18256 121189 -18222
rect 120958 -18448 120993 -18306
rect 121216 -18448 121251 -18306
rect 121349 -18448 121397 -18083
rect 121403 -18448 121451 -18137
rect 121511 -18183 121880 -18149
rect 121611 -18321 121780 -18287
rect 120167 -18506 121522 -18448
rect 119594 -18543 121522 -18506
rect 121549 -18543 121584 -18371
rect 121807 -18543 121842 -18371
rect 121941 -18543 121976 -18245
rect 122985 -18506 123020 -18032
rect 123511 -18036 124186 -18007
rect 123181 -18108 123350 -18074
rect 123119 -18506 123154 -18167
rect 123377 -18506 123412 -18167
rect 123511 -18448 124245 -18036
rect 124264 -18118 124633 -18084
rect 124364 -18256 124533 -18222
rect 124302 -18448 124337 -18306
rect 124560 -18448 124595 -18306
rect 124693 -18448 124741 -18083
rect 124747 -18448 124795 -18137
rect 124855 -18183 125224 -18149
rect 124955 -18321 125124 -18287
rect 123511 -18506 124866 -18448
rect 122938 -18543 124866 -18506
rect 124893 -18543 124928 -18371
rect 125151 -18543 125186 -18371
rect 125285 -18543 125320 -18245
rect 126329 -18506 126364 -18032
rect 126855 -18036 127530 -18007
rect 126525 -18108 126694 -18074
rect 126463 -18506 126498 -18167
rect 126721 -18506 126756 -18167
rect 126855 -18448 127589 -18036
rect 127608 -18118 127977 -18084
rect 127708 -18256 127877 -18222
rect 127646 -18448 127681 -18306
rect 127904 -18448 127939 -18306
rect 128037 -18448 128085 -18083
rect 128091 -18448 128139 -18137
rect 128199 -18183 128568 -18149
rect 128299 -18321 128468 -18287
rect 126855 -18506 128210 -18448
rect 126282 -18543 128210 -18506
rect 128237 -18543 128272 -18371
rect 128495 -18543 128530 -18371
rect 128629 -18543 128664 -18245
rect 129673 -18506 129708 -18032
rect 130199 -18036 130874 -18007
rect 129869 -18108 130038 -18074
rect 129807 -18506 129842 -18167
rect 130065 -18506 130100 -18167
rect 130199 -18448 130933 -18036
rect 130952 -18118 131321 -18084
rect 131052 -18256 131221 -18222
rect 130990 -18448 131025 -18306
rect 131248 -18448 131283 -18306
rect 131381 -18448 131429 -18083
rect 131435 -18448 131483 -18137
rect 131543 -18183 131912 -18149
rect 131643 -18321 131812 -18287
rect 130199 -18506 131554 -18448
rect 129626 -18543 131554 -18506
rect 131581 -18543 131616 -18371
rect 131839 -18543 131874 -18371
rect 131973 -18543 132008 -18245
rect 133017 -18506 133052 -18032
rect 133543 -18036 134218 -18007
rect 133213 -18108 133382 -18074
rect 133151 -18506 133186 -18167
rect 133409 -18506 133444 -18167
rect 133543 -18448 134277 -18036
rect 134296 -18118 134665 -18084
rect 134396 -18256 134565 -18222
rect 134334 -18448 134369 -18306
rect 134592 -18448 134627 -18306
rect 134725 -18448 134773 -18083
rect 134779 -18448 134827 -18137
rect 134887 -18183 135256 -18149
rect 134987 -18321 135156 -18287
rect 133543 -18506 134898 -18448
rect 132970 -18543 134898 -18506
rect 134925 -18543 134960 -18371
rect 135183 -18543 135218 -18371
rect 135317 -18543 135352 -18245
rect 136361 -18506 136396 -18032
rect 136887 -18036 137562 -18007
rect 136557 -18108 136726 -18074
rect 136495 -18506 136530 -18167
rect 136753 -18506 136788 -18167
rect 136887 -18448 137621 -18036
rect 137640 -18118 138009 -18084
rect 137740 -18256 137909 -18222
rect 137678 -18448 137713 -18306
rect 137936 -18448 137971 -18306
rect 138069 -18448 138117 -18083
rect 138123 -18448 138171 -18137
rect 138231 -18183 138600 -18149
rect 138331 -18321 138500 -18287
rect 136887 -18506 138242 -18448
rect 136314 -18543 138242 -18506
rect 138269 -18543 138304 -18371
rect 138527 -18543 138562 -18371
rect 138661 -18543 138696 -18245
rect 139705 -18506 139740 -18032
rect 140231 -18036 140906 -18007
rect 139901 -18108 140070 -18074
rect 139839 -18506 139874 -18167
rect 140097 -18506 140132 -18167
rect 140231 -18448 140965 -18036
rect 140984 -18118 141353 -18084
rect 141084 -18256 141253 -18222
rect 141022 -18448 141057 -18306
rect 141280 -18448 141315 -18306
rect 141413 -18448 141461 -18083
rect 141467 -18448 141515 -18137
rect 141575 -18183 141944 -18149
rect 141675 -18321 141844 -18287
rect 140231 -18506 141586 -18448
rect 139658 -18543 141586 -18506
rect 141613 -18543 141648 -18371
rect 141871 -18543 141906 -18371
rect 142005 -18543 142040 -18245
rect 143049 -18506 143084 -18032
rect 143575 -18036 144250 -18007
rect 143245 -18108 143414 -18074
rect 143183 -18506 143218 -18167
rect 143441 -18506 143476 -18167
rect 143575 -18448 144309 -18036
rect 144328 -18118 144697 -18084
rect 144428 -18256 144597 -18222
rect 144366 -18448 144401 -18306
rect 144624 -18448 144659 -18306
rect 144757 -18448 144805 -18083
rect 144811 -18448 144859 -18137
rect 144919 -18183 145288 -18149
rect 145019 -18321 145188 -18287
rect 143575 -18506 144930 -18448
rect 143002 -18543 144930 -18506
rect 144957 -18543 144992 -18371
rect 145215 -18543 145250 -18371
rect 145349 -18543 145384 -18245
rect 146393 -18506 146428 -18032
rect 146919 -18036 147594 -18007
rect 146589 -18108 146758 -18074
rect 146527 -18506 146562 -18167
rect 146785 -18506 146820 -18167
rect 146919 -18448 147653 -18036
rect 147672 -18118 148041 -18084
rect 147772 -18256 147941 -18222
rect 147710 -18448 147745 -18306
rect 147968 -18448 148003 -18306
rect 148101 -18448 148149 -18083
rect 148155 -18448 148203 -18137
rect 148263 -18183 148632 -18149
rect 148363 -18321 148532 -18287
rect 146919 -18506 148274 -18448
rect 146346 -18543 148274 -18506
rect 148301 -18543 148336 -18371
rect 148559 -18543 148594 -18371
rect 148693 -18543 148728 -18245
rect 149737 -18506 149772 -18032
rect 150263 -18036 150938 -18007
rect 149933 -18108 150102 -18074
rect 149871 -18506 149906 -18167
rect 150129 -18506 150164 -18167
rect 150263 -18448 150997 -18036
rect 151016 -18118 151385 -18084
rect 151116 -18256 151285 -18222
rect 151054 -18448 151089 -18306
rect 151312 -18448 151347 -18306
rect 151445 -18448 151493 -18083
rect 151499 -18448 151547 -18137
rect 151607 -18183 151976 -18149
rect 151707 -18321 151876 -18287
rect 150263 -18506 151618 -18448
rect 149690 -18543 151618 -18506
rect 151645 -18543 151680 -18371
rect 151903 -18543 151938 -18371
rect 152037 -18543 152072 -18245
rect 153081 -18506 153116 -18032
rect 153607 -18036 154282 -18007
rect 153277 -18108 153446 -18074
rect 153215 -18506 153250 -18167
rect 153473 -18506 153508 -18167
rect 153607 -18448 154341 -18036
rect 154360 -18118 154729 -18084
rect 154460 -18256 154629 -18222
rect 154398 -18448 154433 -18306
rect 154656 -18448 154691 -18306
rect 154789 -18448 154837 -18083
rect 154843 -18448 154891 -18137
rect 154951 -18183 155320 -18149
rect 155051 -18321 155220 -18287
rect 153607 -18506 154962 -18448
rect 153034 -18543 154962 -18506
rect 154989 -18543 155024 -18371
rect 155247 -18543 155282 -18371
rect 155381 -18543 155416 -18245
rect 156425 -18506 156460 -18032
rect 156951 -18036 157626 -18007
rect 156621 -18108 156790 -18074
rect 156559 -18506 156594 -18167
rect 156817 -18506 156852 -18167
rect 156951 -18448 157685 -18036
rect 157704 -18118 158073 -18084
rect 157804 -18256 157973 -18222
rect 157742 -18448 157777 -18306
rect 158000 -18448 158035 -18306
rect 158133 -18448 158181 -18083
rect 158187 -18448 158235 -18137
rect 158295 -18183 158664 -18149
rect 158395 -18321 158564 -18287
rect 156951 -18506 158306 -18448
rect 156378 -18543 158306 -18506
rect 158333 -18543 158368 -18371
rect 158591 -18543 158626 -18371
rect 158725 -18543 158760 -18245
rect 159769 -18506 159804 -18032
rect 160295 -18036 160970 -18007
rect 159965 -18108 160134 -18074
rect 159903 -18506 159938 -18167
rect 160161 -18506 160196 -18167
rect 160295 -18448 161029 -18036
rect 161048 -18118 161417 -18084
rect 161148 -18256 161317 -18222
rect 161086 -18448 161121 -18306
rect 161344 -18448 161379 -18306
rect 161477 -18448 161525 -18083
rect 161531 -18448 161579 -18137
rect 161639 -18183 162008 -18149
rect 161739 -18321 161908 -18287
rect 160295 -18506 161650 -18448
rect 159722 -18543 161650 -18506
rect 161677 -18543 161712 -18371
rect 161935 -18543 161970 -18371
rect 162069 -18543 162104 -18245
rect 163113 -18506 163148 -18032
rect 163639 -18036 164314 -18007
rect 163309 -18108 163478 -18074
rect 163247 -18506 163282 -18167
rect 163505 -18506 163540 -18167
rect 163639 -18448 164373 -18036
rect 164392 -18118 164761 -18084
rect 164492 -18256 164661 -18222
rect 164430 -18448 164465 -18306
rect 164688 -18448 164723 -18306
rect 164821 -18448 164869 -18083
rect 164875 -18448 164923 -18137
rect 164983 -18183 165352 -18149
rect 165083 -18321 165252 -18287
rect 163639 -18506 164994 -18448
rect 163066 -18543 164994 -18506
rect 165021 -18543 165056 -18371
rect 165279 -18543 165314 -18371
rect 165413 -18543 165448 -18245
rect 166457 -18506 166492 -18032
rect 166983 -18036 167658 -18007
rect 166653 -18108 166822 -18074
rect 166591 -18506 166626 -18167
rect 166849 -18506 166884 -18167
rect 166983 -18448 167717 -18036
rect 167736 -18118 168105 -18084
rect 167836 -18256 168005 -18222
rect 167774 -18448 167809 -18306
rect 168032 -18448 168067 -18306
rect 168165 -18448 168213 -18083
rect 168219 -18448 168267 -18137
rect 168327 -18183 168696 -18149
rect 168427 -18321 168596 -18287
rect 166983 -18506 168338 -18448
rect 166410 -18543 168338 -18506
rect 168365 -18543 168400 -18371
rect 168623 -18543 168658 -18371
rect 168757 -18543 168792 -18245
rect 169801 -18506 169836 -18032
rect 170327 -18036 171002 -18007
rect 169997 -18108 170166 -18074
rect 169935 -18506 169970 -18167
rect 170193 -18506 170228 -18167
rect 170327 -18448 171061 -18036
rect 171080 -18118 171449 -18084
rect 171180 -18256 171349 -18222
rect 171118 -18448 171153 -18306
rect 171376 -18448 171411 -18306
rect 171509 -18448 171557 -18083
rect 171563 -18448 171611 -18137
rect 171671 -18183 172040 -18149
rect 171771 -18321 171940 -18287
rect 170327 -18506 171682 -18448
rect 169754 -18543 171682 -18506
rect 171709 -18543 171744 -18371
rect 171967 -18543 172002 -18371
rect 172101 -18543 172136 -18245
rect 173145 -18506 173180 -18032
rect 173671 -18036 174346 -18007
rect 173341 -18108 173510 -18074
rect 173279 -18506 173314 -18167
rect 173537 -18506 173572 -18167
rect 173671 -18448 174405 -18036
rect 174424 -18118 174793 -18084
rect 174524 -18256 174693 -18222
rect 174462 -18448 174497 -18306
rect 174720 -18448 174755 -18306
rect 174853 -18448 174901 -18083
rect 174907 -18448 174955 -18137
rect 175015 -18183 175384 -18149
rect 175115 -18321 175284 -18287
rect 173671 -18506 175026 -18448
rect 173098 -18543 175026 -18506
rect 175053 -18543 175088 -18371
rect 175311 -18543 175346 -18371
rect 175445 -18543 175480 -18245
rect 176489 -18506 176524 -18032
rect 177015 -18036 177690 -18007
rect 176685 -18108 176854 -18074
rect 176623 -18506 176658 -18167
rect 176881 -18506 176916 -18167
rect 177015 -18448 177749 -18036
rect 177768 -18118 178137 -18084
rect 177868 -18256 178037 -18222
rect 177806 -18448 177841 -18306
rect 178064 -18448 178099 -18306
rect 178197 -18448 178245 -18083
rect 178251 -18448 178299 -18137
rect 178359 -18183 178728 -18149
rect 178459 -18321 178628 -18287
rect 177015 -18506 178370 -18448
rect 176442 -18543 178370 -18506
rect 178397 -18543 178432 -18371
rect 178655 -18543 178690 -18371
rect 178789 -18543 178824 -18245
rect 179833 -18506 179868 -18032
rect 180359 -18036 181034 -18007
rect 180029 -18108 180198 -18074
rect 179967 -18506 180002 -18167
rect 180225 -18506 180260 -18167
rect 180359 -18448 181093 -18036
rect 181112 -18118 181481 -18084
rect 181212 -18256 181381 -18222
rect 181150 -18448 181185 -18306
rect 181408 -18448 181443 -18306
rect 181541 -18448 181589 -18083
rect 181595 -18448 181643 -18137
rect 181703 -18183 182072 -18149
rect 181803 -18321 181972 -18287
rect 180359 -18506 181714 -18448
rect 179786 -18543 181714 -18506
rect 181741 -18543 181776 -18371
rect 181999 -18543 182034 -18371
rect 182133 -18543 182168 -18245
rect 183177 -18506 183212 -18032
rect 183703 -18036 184378 -18007
rect 183373 -18108 183542 -18074
rect 183311 -18506 183346 -18167
rect 183569 -18506 183604 -18167
rect 183703 -18448 184437 -18036
rect 184456 -18118 184825 -18084
rect 184556 -18256 184725 -18222
rect 184494 -18448 184529 -18306
rect 184752 -18448 184787 -18306
rect 184885 -18448 184933 -18083
rect 184939 -18448 184987 -18137
rect 185047 -18183 185416 -18149
rect 185147 -18321 185316 -18287
rect 183703 -18506 185058 -18448
rect 183130 -18543 185058 -18506
rect 185085 -18543 185120 -18371
rect 185343 -18543 185378 -18371
rect 185477 -18543 185512 -18245
rect 186521 -18506 186556 -18032
rect 187047 -18036 187722 -18007
rect 186717 -18108 186886 -18074
rect 186655 -18506 186690 -18167
rect 186913 -18506 186948 -18167
rect 187047 -18448 187781 -18036
rect 187800 -18118 188169 -18084
rect 187900 -18256 188069 -18222
rect 187838 -18448 187873 -18306
rect 188096 -18448 188131 -18306
rect 188229 -18448 188277 -18083
rect 188283 -18448 188331 -18137
rect 188391 -18183 188760 -18149
rect 188491 -18321 188660 -18287
rect 187047 -18506 188402 -18448
rect 186474 -18543 188402 -18506
rect 188429 -18543 188464 -18371
rect 188687 -18543 188722 -18371
rect 188821 -18543 188856 -18245
rect 189865 -18506 189900 -18032
rect 190391 -18036 191066 -18007
rect 190061 -18108 190230 -18074
rect 189999 -18506 190034 -18167
rect 190257 -18506 190292 -18167
rect 190391 -18448 191125 -18036
rect 191144 -18118 191513 -18084
rect 191244 -18256 191413 -18222
rect 191182 -18448 191217 -18306
rect 191440 -18448 191475 -18306
rect 191573 -18448 191621 -18083
rect 191627 -18448 191675 -18137
rect 191735 -18183 192104 -18149
rect 191835 -18321 192004 -18287
rect 190391 -18506 191746 -18448
rect 189818 -18543 191746 -18506
rect 191773 -18543 191808 -18371
rect 192031 -18543 192066 -18371
rect 192165 -18543 192200 -18245
rect 193209 -18506 193244 -18032
rect 193735 -18036 194410 -18007
rect 193405 -18108 193574 -18074
rect 193343 -18506 193378 -18167
rect 193601 -18506 193636 -18167
rect 193735 -18448 194469 -18036
rect 194488 -18118 194857 -18084
rect 194588 -18256 194757 -18222
rect 194526 -18448 194561 -18306
rect 194784 -18448 194819 -18306
rect 194917 -18448 194965 -18083
rect 194971 -18448 195019 -18137
rect 195079 -18183 195448 -18149
rect 195179 -18321 195348 -18287
rect 193735 -18506 195090 -18448
rect 193162 -18543 195090 -18506
rect 195117 -18543 195152 -18371
rect 195375 -18543 195410 -18371
rect 195509 -18543 195544 -18245
rect 196553 -18506 196588 -18032
rect 197079 -18036 197754 -18007
rect 196749 -18108 196918 -18074
rect 196687 -18506 196722 -18167
rect 196945 -18506 196980 -18167
rect 197079 -18448 197813 -18036
rect 197832 -18118 198201 -18084
rect 197932 -18256 198101 -18222
rect 197870 -18448 197905 -18306
rect 198128 -18448 198163 -18306
rect 198261 -18448 198309 -18083
rect 198315 -18448 198363 -18137
rect 198423 -18183 198792 -18149
rect 198523 -18321 198692 -18287
rect 197079 -18506 198434 -18448
rect 196506 -18543 198434 -18506
rect 198461 -18543 198496 -18371
rect 198719 -18543 198754 -18371
rect 198853 -18543 198888 -18245
rect 199897 -18506 199932 -18032
rect 200423 -18036 201098 -18007
rect 200093 -18108 200262 -18074
rect 200031 -18506 200066 -18167
rect 200289 -18506 200324 -18167
rect 200423 -18448 201157 -18036
rect 201176 -18118 201545 -18084
rect 201276 -18256 201445 -18222
rect 201214 -18448 201249 -18306
rect 201472 -18448 201507 -18306
rect 201605 -18448 201653 -18083
rect 201659 -18448 201707 -18137
rect 201767 -18183 202136 -18149
rect 201867 -18321 202036 -18287
rect 200423 -18506 201778 -18448
rect 199850 -18543 201778 -18506
rect 201805 -18543 201840 -18371
rect 202063 -18543 202098 -18371
rect 202197 -18543 202232 -18245
rect 203241 -18506 203276 -18032
rect 203767 -18036 204442 -18007
rect 203437 -18108 203606 -18074
rect 203375 -18506 203410 -18167
rect 203633 -18506 203668 -18167
rect 203767 -18448 204501 -18036
rect 204520 -18118 204889 -18084
rect 204620 -18256 204789 -18222
rect 204558 -18448 204593 -18306
rect 204816 -18448 204851 -18306
rect 204949 -18448 204997 -18083
rect 205003 -18448 205051 -18137
rect 205111 -18183 205480 -18149
rect 205211 -18321 205380 -18287
rect 203767 -18506 205122 -18448
rect 203194 -18543 205122 -18506
rect 205149 -18543 205184 -18371
rect 205407 -18543 205442 -18371
rect 205541 -18543 205576 -18245
rect 206585 -18506 206620 -18032
rect 207111 -18036 207786 -18007
rect 206781 -18108 206950 -18074
rect 206719 -18506 206754 -18167
rect 206977 -18506 207012 -18167
rect 207111 -18448 207845 -18036
rect 207864 -18118 208233 -18084
rect 207964 -18256 208133 -18222
rect 207902 -18448 207937 -18306
rect 208160 -18448 208195 -18306
rect 208293 -18448 208341 -18083
rect 208347 -18448 208395 -18137
rect 208455 -18183 208824 -18149
rect 208555 -18321 208724 -18287
rect 207111 -18506 208466 -18448
rect 206538 -18543 208466 -18506
rect 208493 -18543 208528 -18371
rect 208751 -18543 208786 -18371
rect 208885 -18543 208920 -18245
rect 209929 -18506 209964 -18032
rect 210455 -18036 211130 -18007
rect 210125 -18108 210294 -18074
rect 210063 -18506 210098 -18167
rect 210321 -18506 210356 -18167
rect 210455 -18448 211189 -18036
rect 211208 -18118 211577 -18084
rect 211308 -18256 211477 -18222
rect 211246 -18448 211281 -18306
rect 211504 -18448 211539 -18306
rect 211637 -18448 211685 -18083
rect 211691 -18448 211739 -18137
rect 211799 -18183 212168 -18149
rect 211899 -18321 212068 -18287
rect 210455 -18506 211810 -18448
rect 209882 -18543 211810 -18506
rect 211837 -18543 211872 -18371
rect 212095 -18543 212130 -18371
rect 212229 -18543 212264 -18245
rect 213273 -18506 213308 -18032
rect 213799 -18036 214474 -18007
rect 217144 -18036 217818 -18007
rect 220488 -18036 221162 -18007
rect 223832 -18036 224506 -18007
rect 227176 -18036 227850 -18007
rect 230520 -18036 231194 -18007
rect 233864 -18036 234538 -18007
rect 237208 -18036 237882 -18007
rect 240552 -18036 241226 -18007
rect 243896 -18036 244570 -18007
rect 247240 -18036 247914 -18007
rect 250584 -18036 251258 -18007
rect 253928 -18036 254602 -18007
rect 257272 -18036 257946 -18007
rect 260616 -18036 261290 -18007
rect 263960 -18036 264634 -18007
rect 267304 -18036 267978 -18007
rect 270648 -18036 271322 -18007
rect 273992 -18036 274666 -18007
rect 277336 -18036 278010 -18007
rect 280680 -18036 281354 -18007
rect 284024 -18036 284698 -18007
rect 287368 -18036 288042 -18007
rect 290712 -18036 291386 -18007
rect 294056 -18036 294730 -18007
rect 297400 -18036 298074 -18007
rect 300744 -18036 301418 -18007
rect 304088 -18036 304762 -18007
rect 307432 -18036 308106 -18007
rect 310776 -18036 311450 -18007
rect 314120 -18036 314794 -18007
rect 317464 -18036 318138 -18007
rect 320808 -18036 321482 -18007
rect 324152 -18036 324826 -18007
rect 327496 -18036 328170 -18007
rect 330840 -18036 331514 -18007
rect 334184 -18036 334858 -18007
rect 337528 -18036 338202 -18007
rect 340872 -18036 341546 -18007
rect 344216 -18036 344890 -18007
rect 347560 -18036 348234 -18007
rect 350904 -18036 351578 -18007
rect 354248 -18036 354922 -18007
rect 357592 -18036 358266 -18007
rect 360936 -18036 361610 -18007
rect 364280 -18036 364954 -18007
rect 367624 -18036 368298 -18007
rect 370968 -18036 371642 -18007
rect 374312 -18036 374986 -18007
rect 377656 -18036 378330 -18007
rect 381000 -18036 381674 -18007
rect 384344 -18036 385018 -18007
rect 387688 -18036 388362 -18007
rect 391032 -18036 391706 -18007
rect 394376 -18036 395050 -18007
rect 397720 -18036 398394 -18007
rect 401064 -18036 401738 -18007
rect 404408 -18036 405082 -18007
rect 407752 -18036 408426 -18007
rect 411096 -18036 411770 -18007
rect 414440 -18036 415114 -18007
rect 417784 -18036 418458 -18007
rect 421128 -18036 421802 -18007
rect 424472 -18036 425146 -18007
rect 427816 -18036 428490 -18007
rect 213469 -18108 213638 -18074
rect 213407 -18506 213442 -18167
rect 213665 -18506 213700 -18167
rect 213799 -18448 214533 -18036
rect 214552 -18118 214921 -18084
rect 214652 -18256 214821 -18222
rect 214590 -18448 214625 -18306
rect 214848 -18448 214883 -18306
rect 214981 -18448 215029 -18083
rect 215035 -18448 215083 -18137
rect 215143 -18183 215512 -18149
rect 215243 -18321 215412 -18287
rect 213799 -18506 215154 -18448
rect 213226 -18543 215154 -18506
rect 215181 -18543 215216 -18371
rect 215439 -18543 215474 -18371
rect 215573 -18543 215608 -18245
rect 217144 -18448 217877 -18036
rect 218326 -18448 218373 -18083
rect 218380 -18448 218427 -18137
rect 220488 -18448 221221 -18036
rect 221670 -18448 221717 -18083
rect 221724 -18448 221771 -18137
rect 223832 -18448 224565 -18036
rect 225014 -18448 225061 -18083
rect 225068 -18448 225115 -18137
rect 227176 -18448 227909 -18036
rect 228358 -18448 228405 -18083
rect 228412 -18448 228459 -18137
rect 230520 -18448 231253 -18036
rect 231702 -18448 231749 -18083
rect 231756 -18448 231803 -18137
rect 233864 -18448 234597 -18036
rect 235046 -18448 235093 -18083
rect 235100 -18448 235147 -18137
rect 237208 -18448 237941 -18036
rect 238390 -18448 238437 -18083
rect 238444 -18448 238491 -18137
rect 240552 -18448 241285 -18036
rect 241734 -18448 241781 -18083
rect 241788 -18448 241835 -18137
rect 243896 -18448 244629 -18036
rect 245078 -18448 245125 -18083
rect 245132 -18448 245179 -18137
rect 247240 -18448 247973 -18036
rect 248422 -18448 248469 -18083
rect 248476 -18448 248523 -18137
rect 250584 -18448 251317 -18036
rect 251766 -18448 251813 -18083
rect 251820 -18448 251867 -18137
rect 253928 -18448 254661 -18036
rect 255110 -18448 255157 -18083
rect 255164 -18448 255211 -18137
rect 257272 -18448 258005 -18036
rect 258454 -18448 258501 -18083
rect 258508 -18448 258555 -18137
rect 260616 -18448 261349 -18036
rect 261798 -18448 261845 -18083
rect 261852 -18448 261899 -18137
rect 263960 -18448 264693 -18036
rect 265142 -18448 265189 -18083
rect 265196 -18448 265243 -18137
rect 267304 -18448 268037 -18036
rect 268486 -18448 268533 -18083
rect 268540 -18448 268587 -18137
rect 270648 -18448 271381 -18036
rect 271830 -18448 271877 -18083
rect 271884 -18448 271931 -18137
rect 273992 -18448 274725 -18036
rect 275174 -18448 275221 -18083
rect 275228 -18448 275275 -18137
rect 277336 -18448 278069 -18036
rect 278518 -18448 278565 -18083
rect 278572 -18448 278619 -18137
rect 280680 -18448 281413 -18036
rect 281862 -18448 281909 -18083
rect 281916 -18448 281963 -18137
rect 284024 -18448 284757 -18036
rect 285206 -18448 285253 -18083
rect 285260 -18448 285307 -18137
rect 287368 -18448 288101 -18036
rect 288550 -18448 288597 -18083
rect 288604 -18448 288651 -18137
rect 290712 -18448 291445 -18036
rect 291894 -18448 291941 -18083
rect 291948 -18448 291995 -18137
rect 294056 -18448 294789 -18036
rect 295238 -18448 295285 -18083
rect 295292 -18448 295339 -18137
rect 297400 -18448 298133 -18036
rect 298582 -18448 298629 -18083
rect 298636 -18448 298683 -18137
rect 300744 -18448 301477 -18036
rect 301926 -18448 301973 -18083
rect 301980 -18448 302027 -18137
rect 304088 -18448 304821 -18036
rect 305270 -18448 305317 -18083
rect 305324 -18448 305371 -18137
rect 307432 -18448 308165 -18036
rect 308614 -18448 308661 -18083
rect 308668 -18448 308715 -18137
rect 310776 -18448 311509 -18036
rect 311958 -18448 312005 -18083
rect 312012 -18448 312059 -18137
rect 314120 -18448 314853 -18036
rect 315302 -18448 315349 -18083
rect 315356 -18448 315403 -18137
rect 317464 -18448 318197 -18036
rect 318646 -18448 318693 -18083
rect 318700 -18448 318747 -18137
rect 320808 -18448 321541 -18036
rect 321990 -18448 322037 -18083
rect 322044 -18448 322091 -18137
rect 324152 -18448 324885 -18036
rect 325334 -18448 325381 -18083
rect 325388 -18448 325435 -18137
rect 327496 -18448 328229 -18036
rect 328678 -18448 328725 -18083
rect 328732 -18448 328779 -18137
rect 330840 -18448 331573 -18036
rect 332022 -18448 332069 -18083
rect 332076 -18448 332123 -18137
rect 334184 -18448 334917 -18036
rect 335366 -18448 335413 -18083
rect 335420 -18448 335467 -18137
rect 337528 -18448 338261 -18036
rect 338710 -18448 338757 -18083
rect 338764 -18448 338811 -18137
rect 340872 -18448 341605 -18036
rect 342054 -18448 342101 -18083
rect 342108 -18448 342155 -18137
rect 344216 -18448 344949 -18036
rect 345398 -18448 345445 -18083
rect 345452 -18448 345499 -18137
rect 347560 -18448 348293 -18036
rect 348742 -18448 348789 -18083
rect 348796 -18448 348843 -18137
rect 350904 -18448 351637 -18036
rect 352086 -18448 352133 -18083
rect 352140 -18448 352187 -18137
rect 354248 -18448 354981 -18036
rect 355430 -18448 355477 -18083
rect 355484 -18448 355531 -18137
rect 357592 -18448 358325 -18036
rect 358774 -18448 358821 -18083
rect 358828 -18448 358875 -18137
rect 360936 -18448 361669 -18036
rect 362118 -18448 362165 -18083
rect 362172 -18448 362219 -18137
rect 364280 -18448 365013 -18036
rect 365462 -18448 365509 -18083
rect 365516 -18448 365563 -18137
rect 367624 -18448 368357 -18036
rect 368806 -18448 368853 -18083
rect 368860 -18448 368907 -18137
rect 370968 -18448 371701 -18036
rect 372150 -18448 372197 -18083
rect 372204 -18448 372251 -18137
rect 374312 -18448 375045 -18036
rect 375494 -18448 375541 -18083
rect 375548 -18448 375595 -18137
rect 377656 -18448 378389 -18036
rect 378838 -18448 378885 -18083
rect 378892 -18448 378939 -18137
rect 381000 -18448 381733 -18036
rect 382182 -18448 382229 -18083
rect 382236 -18448 382283 -18137
rect 384344 -18448 385077 -18036
rect 385526 -18448 385573 -18083
rect 385580 -18448 385627 -18137
rect 387688 -18448 388421 -18036
rect 388870 -18448 388917 -18083
rect 388924 -18448 388971 -18137
rect 391032 -18448 391765 -18036
rect 392214 -18448 392261 -18083
rect 392268 -18448 392315 -18137
rect 394376 -18448 395109 -18036
rect 395558 -18448 395605 -18083
rect 395612 -18448 395659 -18137
rect 397720 -18448 398453 -18036
rect 398902 -18448 398949 -18083
rect 398956 -18448 399003 -18137
rect 401064 -18448 401797 -18036
rect 402246 -18448 402293 -18083
rect 402300 -18448 402347 -18137
rect 404408 -18448 405141 -18036
rect 405590 -18448 405637 -18083
rect 405644 -18448 405691 -18137
rect 407752 -18448 408485 -18036
rect 408934 -18448 408981 -18083
rect 408988 -18448 409035 -18137
rect 411096 -18448 411829 -18036
rect 412278 -18448 412325 -18083
rect 412332 -18448 412379 -18137
rect 414440 -18448 415173 -18036
rect 415622 -18448 415669 -18083
rect 415676 -18448 415723 -18137
rect 417784 -18448 418517 -18036
rect 418966 -18448 419013 -18083
rect 419020 -18448 419067 -18137
rect 421128 -18448 421861 -18036
rect 422310 -18448 422357 -18083
rect 422364 -18448 422411 -18137
rect 424472 -18448 425205 -18036
rect 425654 -18448 425701 -18083
rect 425708 -18448 425755 -18137
rect 427816 -18448 428549 -18036
rect 428998 -18448 429045 -18083
rect 429052 -18448 429099 -18137
rect 217144 -18506 218498 -18448
rect 220488 -18506 221842 -18448
rect 223832 -18506 225186 -18448
rect 227176 -18506 228530 -18448
rect 230520 -18506 231874 -18448
rect 233864 -18506 235218 -18448
rect 237208 -18506 238562 -18448
rect 240552 -18506 241906 -18448
rect 243896 -18506 245250 -18448
rect 247240 -18506 248594 -18448
rect 250584 -18506 251938 -18448
rect 253928 -18506 255282 -18448
rect 257272 -18506 258626 -18448
rect 260616 -18506 261970 -18448
rect 263960 -18506 265314 -18448
rect 267304 -18506 268658 -18448
rect 270648 -18506 272002 -18448
rect 273992 -18506 275346 -18448
rect 277336 -18506 278690 -18448
rect 280680 -18506 282034 -18448
rect 284024 -18506 285378 -18448
rect 287368 -18506 288722 -18448
rect 290712 -18506 292066 -18448
rect 294056 -18506 295410 -18448
rect 297400 -18506 298754 -18448
rect 300744 -18506 302098 -18448
rect 304088 -18506 305442 -18448
rect 307432 -18506 308786 -18448
rect 310776 -18506 312130 -18448
rect 314120 -18506 315474 -18448
rect 317464 -18506 318818 -18448
rect 320808 -18506 322162 -18448
rect 324152 -18506 325506 -18448
rect 327496 -18506 328850 -18448
rect 330840 -18506 332194 -18448
rect 334184 -18506 335538 -18448
rect 337528 -18506 338882 -18448
rect 340872 -18506 342226 -18448
rect 344216 -18506 345570 -18448
rect 347560 -18506 348914 -18448
rect 350904 -18506 352258 -18448
rect 354248 -18506 355602 -18448
rect 357592 -18506 358946 -18448
rect 360936 -18506 362290 -18448
rect 364280 -18506 365634 -18448
rect 367624 -18506 368978 -18448
rect 370968 -18506 372322 -18448
rect 374312 -18506 375666 -18448
rect 377656 -18506 379010 -18448
rect 381000 -18506 382354 -18448
rect 384344 -18506 385698 -18448
rect 387688 -18506 389042 -18448
rect 391032 -18506 392386 -18448
rect 394376 -18506 395730 -18448
rect 397720 -18506 399074 -18448
rect 401064 -18506 402418 -18448
rect 404408 -18506 405762 -18448
rect 407752 -18506 409106 -18448
rect 411096 -18506 412450 -18448
rect 414440 -18506 415794 -18448
rect 417784 -18506 419138 -18448
rect 421128 -18506 422482 -18448
rect 424472 -18506 425826 -18448
rect 427816 -18506 429170 -18448
rect 216571 -18543 218498 -18506
rect 219915 -18543 221842 -18506
rect 223259 -18543 225186 -18506
rect 226603 -18543 228530 -18506
rect 229947 -18543 231874 -18506
rect 233291 -18543 235218 -18506
rect 236635 -18543 238562 -18506
rect 239979 -18543 241906 -18506
rect 243323 -18543 245250 -18506
rect 246667 -18543 248594 -18506
rect 250011 -18543 251938 -18506
rect 253355 -18543 255282 -18506
rect 256699 -18543 258626 -18506
rect 260043 -18543 261970 -18506
rect 263387 -18543 265314 -18506
rect 266731 -18543 268658 -18506
rect 270075 -18543 272002 -18506
rect 273419 -18543 275346 -18506
rect 276763 -18543 278690 -18506
rect 280107 -18543 282034 -18506
rect 283451 -18543 285378 -18506
rect 286795 -18543 288722 -18506
rect 290139 -18543 292066 -18506
rect 293483 -18543 295410 -18506
rect 296827 -18543 298754 -18506
rect 300171 -18543 302098 -18506
rect 303515 -18543 305442 -18506
rect 306859 -18543 308786 -18506
rect 310203 -18543 312130 -18506
rect 313547 -18543 315474 -18506
rect 316891 -18543 318818 -18506
rect 320235 -18543 322162 -18506
rect 323579 -18543 325506 -18506
rect 326923 -18543 328850 -18506
rect 330267 -18543 332194 -18506
rect 333611 -18543 335538 -18506
rect 336955 -18543 338882 -18506
rect 340299 -18543 342226 -18506
rect 343643 -18543 345570 -18506
rect 346987 -18543 348914 -18506
rect 350331 -18543 352258 -18506
rect 353675 -18543 355602 -18506
rect 357019 -18543 358946 -18506
rect 360363 -18543 362290 -18506
rect 363707 -18543 365634 -18506
rect 367051 -18543 368978 -18506
rect 370395 -18543 372322 -18506
rect 373739 -18543 375666 -18506
rect 377083 -18543 379010 -18506
rect 380427 -18543 382354 -18506
rect 383771 -18543 385698 -18506
rect 387115 -18543 389042 -18506
rect 390459 -18543 392386 -18506
rect 393803 -18543 395730 -18506
rect 397147 -18543 399074 -18506
rect 400491 -18543 402418 -18506
rect 403835 -18543 405762 -18506
rect 407179 -18543 409106 -18506
rect 410523 -18543 412450 -18506
rect 413867 -18543 415794 -18506
rect 417211 -18543 419138 -18506
rect 420555 -18543 422482 -18506
rect 423899 -18543 425826 -18506
rect 427243 -18543 429170 -18506
rect 39534 -18667 41768 -18543
rect 42675 -18667 45112 -18543
rect 46019 -18667 48456 -18543
rect 49363 -18667 51800 -18543
rect 52707 -18667 55144 -18543
rect 56052 -18667 58488 -18543
rect 59396 -18667 61832 -18543
rect 62740 -18667 65176 -18543
rect 66084 -18667 68520 -18543
rect 69428 -18667 71864 -18543
rect 72772 -18667 75208 -18543
rect 76116 -18667 78552 -18543
rect 79460 -18667 81896 -18543
rect 82804 -18667 85240 -18543
rect 86148 -18667 88584 -18543
rect 89492 -18667 91928 -18543
rect 92836 -18667 95272 -18543
rect 96180 -18667 98616 -18543
rect 99524 -18667 101960 -18543
rect 102868 -18667 105304 -18543
rect 106212 -18667 108648 -18543
rect 109562 -18667 111992 -18543
rect 112906 -18667 115336 -18543
rect 116250 -18667 118680 -18543
rect 119594 -18667 122024 -18543
rect 122938 -18667 125368 -18543
rect 126282 -18667 128712 -18543
rect 129626 -18667 132056 -18543
rect 132970 -18667 135400 -18543
rect 136314 -18667 138744 -18543
rect 139658 -18667 142088 -18543
rect 143002 -18667 145432 -18543
rect 146346 -18667 148776 -18543
rect 149690 -18667 152120 -18543
rect 153034 -18667 155464 -18543
rect 156378 -18667 158808 -18543
rect 159722 -18667 162152 -18543
rect 163066 -18667 165496 -18543
rect 166410 -18667 168840 -18543
rect 169754 -18667 172184 -18543
rect 173098 -18667 175528 -18543
rect 176442 -18667 178872 -18543
rect 179786 -18667 182216 -18543
rect 183130 -18667 185560 -18543
rect 186474 -18667 188904 -18543
rect 189818 -18667 192248 -18543
rect 193162 -18667 195592 -18543
rect 196506 -18667 198936 -18543
rect 199850 -18667 202280 -18543
rect 203194 -18667 205624 -18543
rect 206538 -18667 208968 -18543
rect 209882 -18667 212312 -18543
rect 213226 -18667 215656 -18543
rect 216571 -18667 219000 -18543
rect 219915 -18667 222344 -18543
rect 223259 -18667 225688 -18543
rect 226603 -18667 229032 -18543
rect 229947 -18667 232376 -18543
rect 233291 -18667 235720 -18543
rect 236635 -18667 239064 -18543
rect 239979 -18667 242408 -18543
rect 243323 -18667 245752 -18543
rect 246667 -18667 249096 -18543
rect 250011 -18667 252440 -18543
rect 253355 -18667 255784 -18543
rect 256699 -18667 259128 -18543
rect 260043 -18667 262472 -18543
rect 263387 -18667 265816 -18543
rect 266731 -18667 269160 -18543
rect 270075 -18667 272504 -18543
rect 273419 -18667 275848 -18543
rect 276763 -18667 279192 -18543
rect 280107 -18667 282536 -18543
rect 283451 -18667 285880 -18543
rect 286795 -18667 289224 -18543
rect 290139 -18667 292568 -18543
rect 293483 -18667 295912 -18543
rect 296827 -18667 299256 -18543
rect 300171 -18667 302600 -18543
rect 303515 -18667 305944 -18543
rect 306859 -18667 309288 -18543
rect 310203 -18667 312632 -18543
rect 313547 -18667 315976 -18543
rect 316891 -18667 319320 -18543
rect 320235 -18667 322664 -18543
rect 323579 -18667 326008 -18543
rect 326923 -18667 329352 -18543
rect 330267 -18667 332696 -18543
rect 333611 -18667 336040 -18543
rect 336955 -18667 339384 -18543
rect 340299 -18667 342728 -18543
rect 343643 -18667 346072 -18543
rect 346987 -18667 349416 -18543
rect 350331 -18667 352760 -18543
rect 353675 -18667 356104 -18543
rect 357019 -18667 359448 -18543
rect 360363 -18667 362792 -18543
rect 363707 -18667 366136 -18543
rect 367051 -18667 369480 -18543
rect 370395 -18667 372824 -18543
rect 373739 -18667 376168 -18543
rect 377083 -18667 379512 -18543
rect 380427 -18667 382856 -18543
rect 383771 -18667 386200 -18543
rect 387115 -18667 389544 -18543
rect 390459 -18667 392888 -18543
rect 393803 -18667 396232 -18543
rect 397147 -18667 399576 -18543
rect 400491 -18667 402920 -18543
rect 403835 -18667 406264 -18543
rect 407179 -18667 409608 -18543
rect 410523 -18667 412952 -18543
rect 413867 -18667 416296 -18543
rect 417211 -18667 419640 -18543
rect 420555 -18667 422984 -18543
rect 423899 -18667 426328 -18543
rect 427243 -18667 429672 -18543
rect 39534 -19622 41821 -18667
rect 42675 -19622 45165 -18667
rect 46019 -19622 48509 -18667
rect 49363 -19622 51853 -18667
rect 52707 -19622 55197 -18667
rect 56052 -19622 58541 -18667
rect 59396 -19622 61885 -18667
rect 62740 -19622 65229 -18667
rect 66084 -19622 68573 -18667
rect 69428 -19622 71917 -18667
rect 72772 -19622 75261 -18667
rect 76116 -19622 78605 -18667
rect 79460 -19622 81949 -18667
rect 82804 -19622 85293 -18667
rect 86148 -19622 88637 -18667
rect 89492 -19622 91981 -18667
rect 92836 -19622 95325 -18667
rect 96180 -19622 98669 -18667
rect 99524 -19622 102013 -18667
rect 102868 -19622 105357 -18667
rect 106212 -19622 108701 -18667
rect 109562 -19622 112045 -18667
rect 112906 -19622 115389 -18667
rect 116250 -19622 118733 -18667
rect 119594 -19622 122077 -18667
rect 122938 -19622 125421 -18667
rect 126282 -19622 128765 -18667
rect 129626 -19622 132109 -18667
rect 132970 -19622 135453 -18667
rect 136314 -19622 138797 -18667
rect 139658 -19622 142141 -18667
rect 143002 -19622 145485 -18667
rect 146346 -19622 148829 -18667
rect 149690 -19622 152173 -18667
rect 153034 -19622 155517 -18667
rect 156378 -19622 158861 -18667
rect 159722 -19622 162205 -18667
rect 163066 -19622 165549 -18667
rect 166410 -19622 168893 -18667
rect 169754 -19622 172237 -18667
rect 173098 -19622 175581 -18667
rect 176442 -19622 178925 -18667
rect 179786 -19622 182269 -18667
rect 183130 -19622 185613 -18667
rect 186474 -19622 188957 -18667
rect 189818 -19622 192301 -18667
rect 193162 -19622 195645 -18667
rect 196506 -19622 198989 -18667
rect 199850 -19622 202333 -18667
rect 203194 -19622 205677 -18667
rect 206538 -19622 209021 -18667
rect 209882 -19622 212365 -18667
rect 213226 -19622 215709 -18667
rect 216571 -19622 219053 -18667
rect 219915 -19622 222397 -18667
rect 223259 -19622 225741 -18667
rect 226603 -19622 229085 -18667
rect 229947 -19622 232429 -18667
rect 233291 -19622 235773 -18667
rect 236635 -19622 239117 -18667
rect 239979 -19622 242461 -18667
rect 243323 -19622 245805 -18667
rect 246667 -19622 249149 -18667
rect 250011 -19622 252493 -18667
rect 253355 -19622 255837 -18667
rect 256699 -19622 259181 -18667
rect 260043 -19622 262525 -18667
rect 263387 -19622 265869 -18667
rect 266731 -19622 269213 -18667
rect 270075 -19622 272557 -18667
rect 273419 -19622 275901 -18667
rect 276763 -19622 279245 -18667
rect 280107 -19622 282589 -18667
rect 283451 -19622 285933 -18667
rect 286795 -19622 289277 -18667
rect 290139 -19622 292621 -18667
rect 293483 -19622 295965 -18667
rect 296827 -19622 299309 -18667
rect 300171 -19622 302653 -18667
rect 303515 -19622 305997 -18667
rect 306859 -19622 309341 -18667
rect 310203 -19622 312685 -18667
rect 313547 -19622 316029 -18667
rect 316891 -19622 319373 -18667
rect 320235 -19622 322717 -18667
rect 323579 -19622 326061 -18667
rect 326923 -19622 329405 -18667
rect 330267 -19622 332749 -18667
rect 333611 -19622 336093 -18667
rect 336955 -19622 339437 -18667
rect 340299 -19622 342781 -18667
rect 343643 -19622 346125 -18667
rect 346987 -19622 349469 -18667
rect 350331 -19622 352813 -18667
rect 353675 -19622 356157 -18667
rect 357019 -19622 359501 -18667
rect 360363 -19622 362845 -18667
rect 363707 -19622 366189 -18667
rect 367051 -19622 369533 -18667
rect 370395 -19622 372877 -18667
rect 373739 -19622 376221 -18667
rect 377083 -19622 379565 -18667
rect 380427 -19622 382909 -18667
rect 383771 -19622 386253 -18667
rect 387115 -19622 389597 -18667
rect 390459 -19622 392941 -18667
rect 393803 -19622 396285 -18667
rect 397147 -19622 399629 -18667
rect 400491 -19622 402973 -18667
rect 403835 -19622 406317 -18667
rect 407179 -19622 409661 -18667
rect 410523 -19622 413005 -18667
rect 413867 -19622 416349 -18667
rect 417211 -19622 419693 -18667
rect 420555 -19622 423037 -18667
rect 423899 -19622 426381 -18667
rect 427243 -19622 429725 -18667
rect 39922 -19687 41821 -19622
rect 43266 -19687 45165 -19622
rect 46610 -19687 48509 -19622
rect 49954 -19687 51853 -19622
rect 53298 -19687 55197 -19622
rect 56643 -19687 58541 -19622
rect 59987 -19687 61885 -19622
rect 63331 -19687 65229 -19622
rect 66675 -19687 68573 -19622
rect 70019 -19687 71917 -19622
rect 73363 -19687 75261 -19622
rect 76707 -19687 78605 -19622
rect 80051 -19687 81949 -19622
rect 83395 -19687 85293 -19622
rect 86739 -19687 88637 -19622
rect 90083 -19687 91981 -19622
rect 93427 -19687 95325 -19622
rect 96771 -19687 98669 -19622
rect 100115 -19687 102013 -19622
rect 103459 -19687 105357 -19622
rect 106803 -19687 108701 -19622
rect 110153 -19687 112045 -19622
rect 113497 -19687 115389 -19622
rect 116841 -19687 118733 -19622
rect 120185 -19687 122077 -19622
rect 123529 -19687 125421 -19622
rect 126873 -19687 128765 -19622
rect 130217 -19687 132109 -19622
rect 133561 -19687 135453 -19622
rect 136905 -19687 138797 -19622
rect 140249 -19687 142141 -19622
rect 143593 -19687 145485 -19622
rect 146937 -19687 148829 -19622
rect 150281 -19687 152173 -19622
rect 153625 -19687 155517 -19622
rect 156969 -19687 158861 -19622
rect 160313 -19687 162205 -19622
rect 163657 -19687 165549 -19622
rect 167001 -19687 168893 -19622
rect 170345 -19687 172237 -19622
rect 173689 -19687 175581 -19622
rect 177033 -19687 178925 -19622
rect 180377 -19687 182269 -19622
rect 183721 -19687 185613 -19622
rect 187065 -19687 188957 -19622
rect 190409 -19687 192301 -19622
rect 193753 -19687 195645 -19622
rect 197097 -19687 198989 -19622
rect 200441 -19687 202333 -19622
rect 203785 -19687 205677 -19622
rect 207129 -19687 209021 -19622
rect 210473 -19687 212365 -19622
rect 213817 -19687 215709 -19622
rect 217162 -19687 219053 -19622
rect 220506 -19687 222397 -19622
rect 223850 -19687 225741 -19622
rect 227194 -19687 229085 -19622
rect 230538 -19687 232429 -19622
rect 233882 -19687 235773 -19622
rect 237226 -19687 239117 -19622
rect 240570 -19687 242461 -19622
rect 243914 -19687 245805 -19622
rect 247258 -19687 249149 -19622
rect 250602 -19687 252493 -19622
rect 253946 -19687 255837 -19622
rect 257290 -19687 259181 -19622
rect 260634 -19687 262525 -19622
rect 263978 -19687 265869 -19622
rect 267322 -19687 269213 -19622
rect 270666 -19687 272557 -19622
rect 274010 -19687 275901 -19622
rect 277354 -19687 279245 -19622
rect 280698 -19687 282589 -19622
rect 284042 -19687 285933 -19622
rect 287386 -19687 289277 -19622
rect 290730 -19687 292621 -19622
rect 294074 -19687 295965 -19622
rect 297418 -19687 299309 -19622
rect 300762 -19687 302653 -19622
rect 304106 -19687 305997 -19622
rect 307450 -19687 309341 -19622
rect 310794 -19687 312685 -19622
rect 314138 -19687 316029 -19622
rect 317482 -19687 319373 -19622
rect 320826 -19687 322717 -19622
rect 324170 -19687 326061 -19622
rect 327514 -19687 329405 -19622
rect 330858 -19687 332749 -19622
rect 334202 -19687 336093 -19622
rect 337546 -19687 339437 -19622
rect 340890 -19687 342781 -19622
rect 344234 -19687 346125 -19622
rect 347578 -19687 349469 -19622
rect 350922 -19687 352813 -19622
rect 354266 -19687 356157 -19622
rect 357610 -19687 359501 -19622
rect 360954 -19687 362845 -19622
rect 364298 -19687 366189 -19622
rect 367642 -19687 369533 -19622
rect 370986 -19687 372877 -19622
rect 374330 -19687 376221 -19622
rect 377674 -19687 379565 -19622
rect 381018 -19687 382909 -19622
rect 384362 -19687 386253 -19622
rect 387706 -19687 389597 -19622
rect 391050 -19687 392941 -19622
rect 394394 -19687 396285 -19622
rect 397738 -19687 399629 -19622
rect 401082 -19687 402973 -19622
rect 404426 -19687 406317 -19622
rect 407770 -19687 409661 -19622
rect 411114 -19687 413005 -19622
rect 414458 -19687 416349 -19622
rect 417802 -19687 419693 -19622
rect 421146 -19687 423037 -19622
rect 424490 -19687 426381 -19622
rect 427834 -19687 429725 -19622
rect 40513 -19747 41821 -19687
rect 43857 -19747 45165 -19687
rect 47201 -19747 48509 -19687
rect 50545 -19747 51853 -19687
rect 53889 -19747 55197 -19687
rect 57234 -19747 58541 -19687
rect 60578 -19747 61885 -19687
rect 63922 -19747 65229 -19687
rect 67266 -19747 68573 -19687
rect 70610 -19747 71917 -19687
rect 73954 -19747 75261 -19687
rect 77298 -19747 78605 -19687
rect 80642 -19747 81949 -19687
rect 83986 -19747 85293 -19687
rect 87330 -19747 88637 -19687
rect 90674 -19747 91981 -19687
rect 94018 -19747 95325 -19687
rect 97362 -19747 98669 -19687
rect 100706 -19747 102013 -19687
rect 104050 -19747 105357 -19687
rect 107394 -19747 108701 -19687
rect 110744 -19747 112045 -19687
rect 114088 -19747 115389 -19687
rect 117432 -19747 118733 -19687
rect 120776 -19747 122077 -19687
rect 124120 -19747 125421 -19687
rect 127464 -19747 128765 -19687
rect 130808 -19747 132109 -19687
rect 134152 -19747 135453 -19687
rect 137496 -19747 138797 -19687
rect 140840 -19747 142141 -19687
rect 144184 -19747 145485 -19687
rect 147528 -19747 148829 -19687
rect 150872 -19747 152173 -19687
rect 154216 -19747 155517 -19687
rect 157560 -19747 158861 -19687
rect 160904 -19747 162205 -19687
rect 164248 -19747 165549 -19687
rect 167592 -19747 168893 -19687
rect 170936 -19747 172237 -19687
rect 174280 -19747 175581 -19687
rect 177624 -19747 178925 -19687
rect 180968 -19747 182269 -19687
rect 184312 -19747 185613 -19687
rect 187656 -19747 188957 -19687
rect 191000 -19747 192301 -19687
rect 194344 -19747 195645 -19687
rect 197688 -19747 198989 -19687
rect 201032 -19747 202333 -19687
rect 204376 -19747 205677 -19687
rect 207720 -19747 209021 -19687
rect 211064 -19747 212365 -19687
rect 214408 -19747 215709 -19687
rect 217753 -19747 219053 -19687
rect 221097 -19747 222397 -19687
rect 224441 -19747 225741 -19687
rect 227785 -19747 229085 -19687
rect 231129 -19747 232429 -19687
rect 234473 -19747 235773 -19687
rect 237817 -19747 239117 -19687
rect 241161 -19747 242461 -19687
rect 244505 -19747 245805 -19687
rect 247849 -19747 249149 -19687
rect 251193 -19747 252493 -19687
rect 254537 -19747 255837 -19687
rect 257881 -19747 259181 -19687
rect 261225 -19747 262525 -19687
rect 264569 -19747 265869 -19687
rect 267913 -19747 269213 -19687
rect 271257 -19747 272557 -19687
rect 274601 -19747 275901 -19687
rect 277945 -19747 279245 -19687
rect 281289 -19747 282589 -19687
rect 284633 -19747 285933 -19687
rect 287977 -19747 289277 -19687
rect 291321 -19747 292621 -19687
rect 294665 -19747 295965 -19687
rect 298009 -19747 299309 -19687
rect 301353 -19747 302653 -19687
rect 304697 -19747 305997 -19687
rect 308041 -19747 309341 -19687
rect 311385 -19747 312685 -19687
rect 314729 -19747 316029 -19687
rect 318073 -19747 319373 -19687
rect 321417 -19747 322717 -19687
rect 324761 -19747 326061 -19687
rect 328105 -19747 329405 -19687
rect 331449 -19747 332749 -19687
rect 334793 -19747 336093 -19687
rect 338137 -19747 339437 -19687
rect 341481 -19747 342781 -19687
rect 344825 -19747 346125 -19687
rect 348169 -19747 349469 -19687
rect 351513 -19747 352813 -19687
rect 354857 -19747 356157 -19687
rect 358201 -19747 359501 -19687
rect 361545 -19747 362845 -19687
rect 364889 -19747 366189 -19687
rect 368233 -19747 369533 -19687
rect 371577 -19747 372877 -19687
rect 374921 -19747 376221 -19687
rect 378265 -19747 379565 -19687
rect 381609 -19747 382909 -19687
rect 384953 -19747 386253 -19687
rect 388297 -19747 389597 -19687
rect 391641 -19747 392941 -19687
rect 394985 -19747 396285 -19687
rect 398329 -19747 399629 -19687
rect 401673 -19747 402973 -19687
rect 405017 -19747 406317 -19687
rect 408361 -19747 409661 -19687
rect 411705 -19747 413005 -19687
rect 415049 -19747 416349 -19687
rect 418393 -19747 419693 -19687
rect 421737 -19747 423037 -19687
rect 425081 -19747 426381 -19687
rect 428425 -19747 429725 -19687
rect 40542 -19752 41821 -19747
rect 43886 -19752 45165 -19747
rect 47230 -19752 48509 -19747
rect 50574 -19752 51853 -19747
rect 53918 -19752 55197 -19747
rect 57263 -19752 58541 -19747
rect 60607 -19752 61885 -19747
rect 63951 -19752 65229 -19747
rect 67295 -19752 68573 -19747
rect 70639 -19752 71917 -19747
rect 73983 -19752 75261 -19747
rect 77327 -19752 78605 -19747
rect 80671 -19752 81949 -19747
rect 84015 -19752 85293 -19747
rect 87359 -19752 88637 -19747
rect 90703 -19752 91981 -19747
rect 94047 -19752 95325 -19747
rect 97391 -19752 98669 -19747
rect 100735 -19752 102013 -19747
rect 104079 -19752 105357 -19747
rect 107423 -19752 108701 -19747
rect 110773 -19752 112045 -19747
rect 114117 -19752 115389 -19747
rect 117461 -19752 118733 -19747
rect 120805 -19752 122077 -19747
rect 124149 -19752 125421 -19747
rect 127493 -19752 128765 -19747
rect 130837 -19752 132109 -19747
rect 134181 -19752 135453 -19747
rect 137525 -19752 138797 -19747
rect 140869 -19752 142141 -19747
rect 144213 -19752 145485 -19747
rect 147557 -19752 148829 -19747
rect 150901 -19752 152173 -19747
rect 154245 -19752 155517 -19747
rect 157589 -19752 158861 -19747
rect 160933 -19752 162205 -19747
rect 164277 -19752 165549 -19747
rect 167621 -19752 168893 -19747
rect 170965 -19752 172237 -19747
rect 174309 -19752 175581 -19747
rect 177653 -19752 178925 -19747
rect 180997 -19752 182269 -19747
rect 184341 -19752 185613 -19747
rect 187685 -19752 188957 -19747
rect 191029 -19752 192301 -19747
rect 194373 -19752 195645 -19747
rect 197717 -19752 198989 -19747
rect 201061 -19752 202333 -19747
rect 204405 -19752 205677 -19747
rect 207749 -19752 209021 -19747
rect 211093 -19752 212365 -19747
rect 214437 -19752 215709 -19747
rect 217782 -19752 219053 -19747
rect 221126 -19752 222397 -19747
rect 224470 -19752 225741 -19747
rect 227814 -19752 229085 -19747
rect 231158 -19752 232429 -19747
rect 234502 -19752 235773 -19747
rect 237846 -19752 239117 -19747
rect 241190 -19752 242461 -19747
rect 244534 -19752 245805 -19747
rect 247878 -19752 249149 -19747
rect 251222 -19752 252493 -19747
rect 254566 -19752 255837 -19747
rect 257910 -19752 259181 -19747
rect 261254 -19752 262525 -19747
rect 264598 -19752 265869 -19747
rect 267942 -19752 269213 -19747
rect 271286 -19752 272557 -19747
rect 274630 -19752 275901 -19747
rect 277974 -19752 279245 -19747
rect 281318 -19752 282589 -19747
rect 284662 -19752 285933 -19747
rect 288006 -19752 289277 -19747
rect 291350 -19752 292621 -19747
rect 294694 -19752 295965 -19747
rect 298038 -19752 299309 -19747
rect 301382 -19752 302653 -19747
rect 304726 -19752 305997 -19747
rect 308070 -19752 309341 -19747
rect 311414 -19752 312685 -19747
rect 314758 -19752 316029 -19747
rect 318102 -19752 319373 -19747
rect 321446 -19752 322717 -19747
rect 324790 -19752 326061 -19747
rect 328134 -19752 329405 -19747
rect 331478 -19752 332749 -19747
rect 334822 -19752 336093 -19747
rect 338166 -19752 339437 -19747
rect 341510 -19752 342781 -19747
rect 344854 -19752 346125 -19747
rect 348198 -19752 349469 -19747
rect 351542 -19752 352813 -19747
rect 354886 -19752 356157 -19747
rect 358230 -19752 359501 -19747
rect 361574 -19752 362845 -19747
rect 364918 -19752 366189 -19747
rect 368262 -19752 369533 -19747
rect 371606 -19752 372877 -19747
rect 374950 -19752 376221 -19747
rect 378294 -19752 379565 -19747
rect 381638 -19752 382909 -19747
rect 384982 -19752 386253 -19747
rect 388326 -19752 389597 -19747
rect 391670 -19752 392941 -19747
rect 395014 -19752 396285 -19747
rect 398358 -19752 399629 -19747
rect 401702 -19752 402973 -19747
rect 405046 -19752 406317 -19747
rect 408390 -19752 409661 -19747
rect 411734 -19752 413005 -19747
rect 415078 -19752 416349 -19747
rect 418422 -19752 419693 -19747
rect 421766 -19752 423037 -19747
rect 425110 -19752 426381 -19747
rect 428454 -19752 429725 -19747
rect 40674 -19770 41821 -19752
rect 44018 -19770 45165 -19752
rect 47362 -19770 48509 -19752
rect 50706 -19770 51853 -19752
rect 54050 -19770 55197 -19752
rect 57394 -19770 58541 -19752
rect 60738 -19770 61885 -19752
rect 64082 -19770 65229 -19752
rect 67426 -19770 68573 -19752
rect 70770 -19770 71917 -19752
rect 74114 -19770 75261 -19752
rect 77458 -19770 78605 -19752
rect 80802 -19770 81949 -19752
rect 84146 -19770 85293 -19752
rect 87490 -19770 88637 -19752
rect 90834 -19770 91981 -19752
rect 94178 -19770 95325 -19752
rect 97522 -19770 98669 -19752
rect 100866 -19770 102013 -19752
rect 104210 -19770 105357 -19752
rect 107554 -19770 108701 -19752
rect 110898 -19770 112045 -19752
rect 114242 -19770 115389 -19752
rect 117586 -19770 118733 -19752
rect 120930 -19770 122077 -19752
rect 124274 -19770 125421 -19752
rect 127618 -19770 128765 -19752
rect 130962 -19770 132109 -19752
rect 134306 -19770 135453 -19752
rect 137650 -19770 138797 -19752
rect 140994 -19770 142141 -19752
rect 144338 -19770 145485 -19752
rect 147682 -19770 148829 -19752
rect 151026 -19770 152173 -19752
rect 154370 -19770 155517 -19752
rect 157714 -19770 158861 -19752
rect 161058 -19770 162205 -19752
rect 164402 -19770 165549 -19752
rect 167746 -19770 168893 -19752
rect 171090 -19770 172237 -19752
rect 174434 -19770 175581 -19752
rect 177778 -19770 178925 -19752
rect 181122 -19770 182269 -19752
rect 184466 -19770 185613 -19752
rect 187810 -19770 188957 -19752
rect 191154 -19770 192301 -19752
rect 194498 -19770 195645 -19752
rect 197842 -19770 198989 -19752
rect 201186 -19770 202333 -19752
rect 204530 -19770 205677 -19752
rect 207874 -19770 209021 -19752
rect 211218 -19770 212365 -19752
rect 214562 -19770 215709 -19752
rect 217906 -19770 219053 -19752
rect 221250 -19770 222397 -19752
rect 224594 -19770 225741 -19752
rect 227938 -19770 229085 -19752
rect 231282 -19770 232429 -19752
rect 234626 -19770 235773 -19752
rect 237970 -19770 239117 -19752
rect 241314 -19770 242461 -19752
rect 244658 -19770 245805 -19752
rect 248002 -19770 249149 -19752
rect 251346 -19770 252493 -19752
rect 254690 -19770 255837 -19752
rect 258034 -19770 259181 -19752
rect 261378 -19770 262525 -19752
rect 264722 -19770 265869 -19752
rect 268066 -19770 269213 -19752
rect 271410 -19770 272557 -19752
rect 274754 -19770 275901 -19752
rect 278098 -19770 279245 -19752
rect 281442 -19770 282589 -19752
rect 284786 -19770 285933 -19752
rect 288130 -19770 289277 -19752
rect 291474 -19770 292621 -19752
rect 294818 -19770 295965 -19752
rect 298162 -19770 299309 -19752
rect 301506 -19770 302653 -19752
rect 304850 -19770 305997 -19752
rect 308194 -19770 309341 -19752
rect 311538 -19770 312685 -19752
rect 314882 -19770 316029 -19752
rect 318226 -19770 319373 -19752
rect 321570 -19770 322717 -19752
rect 324914 -19770 326061 -19752
rect 328258 -19770 329405 -19752
rect 331602 -19770 332749 -19752
rect 334946 -19770 336093 -19752
rect 338290 -19770 339437 -19752
rect 341634 -19770 342781 -19752
rect 344978 -19770 346125 -19752
rect 348322 -19770 349469 -19752
rect 351666 -19770 352813 -19752
rect 355010 -19770 356157 -19752
rect 358354 -19770 359501 -19752
rect 361698 -19770 362845 -19752
rect 365042 -19770 366189 -19752
rect 368386 -19770 369533 -19752
rect 371730 -19770 372877 -19752
rect 375074 -19770 376221 -19752
rect 378418 -19770 379565 -19752
rect 381762 -19770 382909 -19752
rect 385106 -19770 386253 -19752
rect 388450 -19770 389597 -19752
rect 391794 -19770 392941 -19752
rect 395138 -19770 396285 -19752
rect 398482 -19770 399629 -19752
rect 401826 -19770 402973 -19752
rect 405170 -19770 406317 -19752
rect 408514 -19770 409661 -19752
rect 411858 -19770 413005 -19752
rect 415202 -19770 416349 -19752
rect 418546 -19770 419693 -19752
rect 421890 -19770 423037 -19752
rect 425234 -19770 426381 -19752
rect 428578 -19770 429725 -19752
rect 41104 -19781 41821 -19770
rect 44448 -19781 45165 -19770
rect 47792 -19781 48509 -19770
rect 51136 -19781 51853 -19770
rect 54480 -19781 55197 -19770
rect 57825 -19781 58541 -19770
rect 61169 -19781 61885 -19770
rect 64513 -19781 65229 -19770
rect 67857 -19781 68573 -19770
rect 71201 -19781 71917 -19770
rect 74545 -19781 75261 -19770
rect 77889 -19781 78605 -19770
rect 81233 -19781 81949 -19770
rect 84577 -19781 85293 -19770
rect 87921 -19781 88637 -19770
rect 91265 -19781 91981 -19770
rect 94609 -19781 95325 -19770
rect 97953 -19781 98669 -19770
rect 101297 -19781 102013 -19770
rect 104641 -19781 105357 -19770
rect 107985 -19781 108701 -19770
rect 111335 -19781 112045 -19770
rect 114679 -19781 115389 -19770
rect 118023 -19781 118733 -19770
rect 121367 -19781 122077 -19770
rect 124711 -19781 125421 -19770
rect 128055 -19781 128765 -19770
rect 131399 -19781 132109 -19770
rect 134743 -19781 135453 -19770
rect 138087 -19781 138797 -19770
rect 141431 -19781 142141 -19770
rect 144775 -19781 145485 -19770
rect 148119 -19781 148829 -19770
rect 151463 -19781 152173 -19770
rect 154807 -19781 155517 -19770
rect 158151 -19781 158861 -19770
rect 161495 -19781 162205 -19770
rect 164839 -19781 165549 -19770
rect 168183 -19781 168893 -19770
rect 171527 -19781 172237 -19770
rect 174871 -19781 175581 -19770
rect 178215 -19781 178925 -19770
rect 181559 -19781 182269 -19770
rect 184903 -19781 185613 -19770
rect 188247 -19781 188957 -19770
rect 191591 -19781 192301 -19770
rect 194935 -19781 195645 -19770
rect 198279 -19781 198989 -19770
rect 201623 -19781 202333 -19770
rect 204967 -19781 205677 -19770
rect 208311 -19781 209021 -19770
rect 211655 -19781 212365 -19770
rect 214999 -19781 215709 -19770
rect 218344 -19781 219053 -19770
rect 221688 -19781 222397 -19770
rect 225032 -19781 225741 -19770
rect 228376 -19781 229085 -19770
rect 231720 -19781 232429 -19770
rect 235064 -19781 235773 -19770
rect 238408 -19781 239117 -19770
rect 241752 -19781 242461 -19770
rect 245096 -19781 245805 -19770
rect 248440 -19781 249149 -19770
rect 251784 -19781 252493 -19770
rect 255128 -19781 255837 -19770
rect 258472 -19781 259181 -19770
rect 261816 -19781 262525 -19770
rect 265160 -19781 265869 -19770
rect 268504 -19781 269213 -19770
rect 271848 -19781 272557 -19770
rect 275192 -19781 275901 -19770
rect 278536 -19781 279245 -19770
rect 281880 -19781 282589 -19770
rect 285224 -19781 285933 -19770
rect 288568 -19781 289277 -19770
rect 291912 -19781 292621 -19770
rect 295256 -19781 295965 -19770
rect 298600 -19781 299309 -19770
rect 301944 -19781 302653 -19770
rect 305288 -19781 305997 -19770
rect 308632 -19781 309341 -19770
rect 311976 -19781 312685 -19770
rect 315320 -19781 316029 -19770
rect 318664 -19781 319373 -19770
rect 322008 -19781 322717 -19770
rect 325352 -19781 326061 -19770
rect 328696 -19781 329405 -19770
rect 332040 -19781 332749 -19770
rect 335384 -19781 336093 -19770
rect 338728 -19781 339437 -19770
rect 342072 -19781 342781 -19770
rect 345416 -19781 346125 -19770
rect 348760 -19781 349469 -19770
rect 352104 -19781 352813 -19770
rect 355448 -19781 356157 -19770
rect 358792 -19781 359501 -19770
rect 362136 -19781 362845 -19770
rect 365480 -19781 366189 -19770
rect 368824 -19781 369533 -19770
rect 372168 -19781 372877 -19770
rect 375512 -19781 376221 -19770
rect 378856 -19781 379565 -19770
rect 382200 -19781 382909 -19770
rect 385544 -19781 386253 -19770
rect 388888 -19781 389597 -19770
rect 392232 -19781 392941 -19770
rect 395576 -19781 396285 -19770
rect 398920 -19781 399629 -19770
rect 402264 -19781 402973 -19770
rect 405608 -19781 406317 -19770
rect 408952 -19781 409661 -19770
rect 412296 -19781 413005 -19770
rect 415640 -19781 416349 -19770
rect 418984 -19781 419693 -19770
rect 422328 -19781 423037 -19770
rect 425672 -19781 426381 -19770
rect 429016 -19781 429725 -19770
rect 38424 -19817 38442 -19781
rect 41104 -19817 41786 -19781
rect 44448 -19817 45130 -19781
rect 47792 -19817 48474 -19781
rect 51136 -19817 51818 -19781
rect 54480 -19817 55162 -19781
rect 57825 -19817 58506 -19781
rect 61169 -19817 61850 -19781
rect 64513 -19817 65194 -19781
rect 67857 -19817 68538 -19781
rect 71201 -19817 71882 -19781
rect 74545 -19817 75226 -19781
rect 77889 -19817 78570 -19781
rect 81233 -19817 81914 -19781
rect 84577 -19817 85258 -19781
rect 87921 -19817 88602 -19781
rect 91265 -19817 91946 -19781
rect 94609 -19817 95290 -19781
rect 97953 -19817 98634 -19781
rect 101297 -19817 101978 -19781
rect 104641 -19817 105322 -19781
rect 107985 -19817 108666 -19781
rect 111335 -19817 112010 -19781
rect 114679 -19817 115354 -19781
rect 118023 -19817 118698 -19781
rect 121367 -19817 122042 -19781
rect 124711 -19817 125386 -19781
rect 128055 -19817 128730 -19781
rect 131399 -19817 132074 -19781
rect 134743 -19817 135418 -19781
rect 138087 -19817 138762 -19781
rect 141431 -19817 142106 -19781
rect 144775 -19817 145450 -19781
rect 148119 -19817 148794 -19781
rect 151463 -19817 152138 -19781
rect 154807 -19817 155482 -19781
rect 158151 -19817 158826 -19781
rect 161495 -19817 162170 -19781
rect 164839 -19817 165514 -19781
rect 168183 -19817 168858 -19781
rect 171527 -19817 172202 -19781
rect 174871 -19817 175546 -19781
rect 178215 -19817 178890 -19781
rect 181559 -19817 182234 -19781
rect 184903 -19817 185578 -19781
rect 188247 -19817 188922 -19781
rect 191591 -19817 192266 -19781
rect 194935 -19817 195610 -19781
rect 198279 -19817 198954 -19781
rect 201623 -19817 202298 -19781
rect 204967 -19817 205642 -19781
rect 208311 -19817 208986 -19781
rect 211655 -19817 212330 -19781
rect 214999 -19817 215674 -19781
rect 218344 -19817 219018 -19781
rect 221688 -19817 222362 -19781
rect 225032 -19817 225706 -19781
rect 228376 -19817 229050 -19781
rect 231720 -19817 232394 -19781
rect 235064 -19817 235738 -19781
rect 238408 -19817 239082 -19781
rect 241752 -19817 242426 -19781
rect 245096 -19817 245770 -19781
rect 248440 -19817 249114 -19781
rect 251784 -19817 252458 -19781
rect 255128 -19817 255802 -19781
rect 258472 -19817 259146 -19781
rect 261816 -19817 262490 -19781
rect 265160 -19817 265834 -19781
rect 268504 -19817 269178 -19781
rect 271848 -19817 272522 -19781
rect 275192 -19817 275866 -19781
rect 278536 -19817 279210 -19781
rect 281880 -19817 282554 -19781
rect 285224 -19817 285898 -19781
rect 288568 -19817 289242 -19781
rect 291912 -19817 292586 -19781
rect 295256 -19817 295930 -19781
rect 298600 -19817 299274 -19781
rect 301944 -19817 302618 -19781
rect 305288 -19817 305962 -19781
rect 308632 -19817 309306 -19781
rect 311976 -19817 312650 -19781
rect 315320 -19817 315994 -19781
rect 318664 -19817 319338 -19781
rect 322008 -19817 322682 -19781
rect 325352 -19817 326026 -19781
rect 328696 -19817 329370 -19781
rect 332040 -19817 332714 -19781
rect 335384 -19817 336058 -19781
rect 338728 -19817 339402 -19781
rect 342072 -19817 342746 -19781
rect 345416 -19817 346090 -19781
rect 348760 -19817 349434 -19781
rect 352104 -19817 352778 -19781
rect 355448 -19817 356122 -19781
rect 358792 -19817 359466 -19781
rect 362136 -19817 362810 -19781
rect 365480 -19817 366154 -19781
rect 368824 -19817 369498 -19781
rect 372168 -19817 372842 -19781
rect 375512 -19817 376186 -19781
rect 378856 -19817 379530 -19781
rect 382200 -19817 382874 -19781
rect 385544 -19817 386218 -19781
rect 388888 -19817 389562 -19781
rect 392232 -19817 392906 -19781
rect 395576 -19817 396250 -19781
rect 398920 -19817 399594 -19781
rect 402264 -19817 402938 -19781
rect 405608 -19817 406282 -19781
rect 408952 -19817 409626 -19781
rect 412296 -19817 412970 -19781
rect 415640 -19817 416314 -19781
rect 418984 -19817 419658 -19781
rect 422328 -19817 423002 -19781
rect 425672 -19817 426346 -19781
rect 429016 -19817 429690 -19781
rect 38274 -19835 38442 -19817
rect 41295 -19835 41786 -19817
rect 44639 -19835 45130 -19817
rect 47983 -19835 48474 -19817
rect 51327 -19835 51818 -19817
rect 54671 -19835 55162 -19817
rect 58015 -19835 58506 -19817
rect 61359 -19835 61850 -19817
rect 64703 -19835 65194 -19817
rect 68047 -19835 68538 -19817
rect 71391 -19835 71882 -19817
rect 74735 -19835 75226 -19817
rect 78079 -19835 78570 -19817
rect 81423 -19835 81914 -19817
rect 84767 -19835 85258 -19817
rect 88111 -19835 88602 -19817
rect 91455 -19835 91946 -19817
rect 94799 -19835 95290 -19817
rect 98143 -19835 98634 -19817
rect 101487 -19835 101978 -19817
rect 104831 -19835 105322 -19817
rect 108175 -19835 108666 -19817
rect 111519 -19835 112010 -19817
rect 114863 -19835 115354 -19817
rect 118207 -19835 118698 -19817
rect 121551 -19835 122042 -19817
rect 124895 -19835 125386 -19817
rect 128239 -19835 128730 -19817
rect 131583 -19835 132074 -19817
rect 134927 -19835 135418 -19817
rect 138271 -19835 138762 -19817
rect 141615 -19835 142106 -19817
rect 144959 -19835 145450 -19817
rect 148303 -19835 148794 -19817
rect 151647 -19835 152138 -19817
rect 154991 -19835 155482 -19817
rect 158335 -19835 158826 -19817
rect 161679 -19835 162170 -19817
rect 165023 -19835 165514 -19817
rect 168367 -19835 168858 -19817
rect 171711 -19835 172202 -19817
rect 175055 -19835 175546 -19817
rect 178399 -19835 178890 -19817
rect 181743 -19835 182234 -19817
rect 185087 -19835 185578 -19817
rect 188431 -19835 188922 -19817
rect 191775 -19835 192266 -19817
rect 195119 -19835 195610 -19817
rect 198463 -19835 198954 -19817
rect 201807 -19835 202298 -19817
rect 205151 -19835 205642 -19817
rect 208495 -19835 208986 -19817
rect 211839 -19835 212330 -19817
rect 215183 -19835 215674 -19817
rect 218527 -19835 219018 -19817
rect 221871 -19835 222362 -19817
rect 225215 -19835 225706 -19817
rect 228559 -19835 229050 -19817
rect 231903 -19835 232394 -19817
rect 235247 -19835 235738 -19817
rect 238591 -19835 239082 -19817
rect 241935 -19835 242426 -19817
rect 245279 -19835 245770 -19817
rect 248623 -19835 249114 -19817
rect 251967 -19835 252458 -19817
rect 255311 -19835 255802 -19817
rect 258655 -19835 259146 -19817
rect 261999 -19835 262490 -19817
rect 265343 -19835 265834 -19817
rect 268687 -19835 269178 -19817
rect 272031 -19835 272522 -19817
rect 275375 -19835 275866 -19817
rect 278719 -19835 279210 -19817
rect 282063 -19835 282554 -19817
rect 285407 -19835 285898 -19817
rect 288751 -19835 289242 -19817
rect 292095 -19835 292586 -19817
rect 295439 -19835 295930 -19817
rect 298783 -19835 299274 -19817
rect 302127 -19835 302618 -19817
rect 305471 -19835 305962 -19817
rect 308815 -19835 309306 -19817
rect 312159 -19835 312650 -19817
rect 315503 -19835 315994 -19817
rect 318847 -19835 319338 -19817
rect 322191 -19835 322682 -19817
rect 325535 -19835 326026 -19817
rect 328879 -19835 329370 -19817
rect 332223 -19835 332714 -19817
rect 335567 -19835 336058 -19817
rect 338911 -19835 339402 -19817
rect 342255 -19835 342746 -19817
rect 345599 -19835 346090 -19817
rect 348943 -19835 349434 -19817
rect 352287 -19835 352778 -19817
rect 355631 -19835 356122 -19817
rect 358975 -19835 359466 -19817
rect 362319 -19835 362810 -19817
rect 365663 -19835 366154 -19817
rect 369007 -19835 369498 -19817
rect 372351 -19835 372842 -19817
rect 375695 -19835 376186 -19817
rect 379039 -19835 379530 -19817
rect 382383 -19835 382874 -19817
rect 385727 -19835 386218 -19817
rect 389071 -19835 389562 -19817
rect 392415 -19835 392906 -19817
rect 395759 -19835 396250 -19817
rect 399103 -19835 399594 -19817
rect 402447 -19835 402938 -19817
rect 405791 -19835 406282 -19817
rect 409135 -19835 409626 -19817
rect 412479 -19835 412970 -19817
rect 415823 -19835 416314 -19817
rect 419167 -19835 419658 -19817
rect 422511 -19835 423002 -19817
rect 425855 -19835 426346 -19817
rect 429199 -19835 429690 -19817
rect 38274 -19859 38369 -19835
rect 41337 -19859 41713 -19835
rect 44681 -19859 45057 -19835
rect 48025 -19859 48401 -19835
rect 51369 -19859 51745 -19835
rect 54713 -19859 55089 -19835
rect 58058 -19859 58433 -19835
rect 61402 -19859 61777 -19835
rect 64746 -19859 65121 -19835
rect 68090 -19859 68465 -19835
rect 71434 -19859 71809 -19835
rect 74778 -19859 75153 -19835
rect 78122 -19859 78497 -19835
rect 81466 -19859 81841 -19835
rect 84810 -19859 85185 -19835
rect 88154 -19859 88529 -19835
rect 91498 -19859 91873 -19835
rect 94842 -19859 95217 -19835
rect 98186 -19859 98561 -19835
rect 101530 -19859 101905 -19835
rect 104874 -19859 105249 -19835
rect 108218 -19859 108593 -19835
rect 111568 -19859 111937 -19835
rect 114912 -19859 115281 -19835
rect 118256 -19859 118625 -19835
rect 121600 -19859 121969 -19835
rect 124944 -19859 125313 -19835
rect 128288 -19859 128657 -19835
rect 131632 -19859 132001 -19835
rect 134976 -19859 135345 -19835
rect 138320 -19859 138689 -19835
rect 141664 -19859 142033 -19835
rect 145008 -19859 145377 -19835
rect 148352 -19859 148721 -19835
rect 151696 -19859 152065 -19835
rect 155040 -19859 155409 -19835
rect 158384 -19859 158753 -19835
rect 161728 -19859 162097 -19835
rect 165072 -19859 165441 -19835
rect 168416 -19859 168785 -19835
rect 171760 -19859 172129 -19835
rect 175104 -19859 175473 -19835
rect 178448 -19859 178817 -19835
rect 181792 -19859 182161 -19835
rect 185136 -19859 185505 -19835
rect 188480 -19859 188849 -19835
rect 191824 -19859 192193 -19835
rect 195168 -19859 195537 -19835
rect 198512 -19859 198881 -19835
rect 201856 -19859 202225 -19835
rect 205200 -19859 205569 -19835
rect 208544 -19859 208913 -19835
rect 211888 -19859 212257 -19835
rect 215232 -19859 215601 -19835
rect 2424 -25666 2462 -25641
rect 4890 -25709 4928 -25684
rect 7356 -25752 7394 -25727
rect 9822 -25795 9860 -25770
rect 12288 -25838 12326 -25813
rect 14754 -25881 14792 -25856
rect 17220 -25924 17258 -25899
rect 19686 -25967 19724 -25942
rect 22152 -26010 22190 -25985
rect 24618 -26053 24656 -26028
rect 27084 -26096 27122 -26071
rect 29550 -26139 29588 -26114
rect 32016 -26182 32054 -26157
rect 34482 -26225 34520 -26200
<< error_s >>
rect -9 -11275 25 -10475
rect 125 -11167 159 -11145
rect 383 -11167 417 -11145
rect 113 -11179 429 -11167
rect 95 -11213 429 -11179
rect 113 -11225 429 -11213
rect -9 -12475 33 -11275
rect 125 -11283 159 -11225
rect 383 -11270 417 -11225
rect 125 -11385 165 -11283
rect 363 -11311 417 -11270
rect 183 -11317 193 -11311
rect 349 -11317 417 -11311
rect 179 -11351 193 -11317
rect 195 -11351 417 -11317
rect 183 -11357 193 -11351
rect 349 -11357 417 -11351
rect 371 -11385 417 -11357
rect 125 -11410 159 -11385
rect 371 -11398 379 -11385
rect 125 -12367 167 -11410
rect 171 -12367 178 -11399
rect 383 -11410 417 -11385
rect 517 -11275 551 -10475
rect 383 -12367 425 -11410
rect 113 -12379 437 -12367
rect 517 -12379 559 -11275
rect 3220 -12079 5718 0
rect 3191 -12127 5718 -12079
rect 1268 -12161 5718 -12127
rect 113 -12413 671 -12379
rect 113 -12425 437 -12413
rect -11 -13129 33 -12475
rect 125 -12610 167 -12425
rect 171 -12501 178 -12425
rect 383 -12470 425 -12425
rect 383 -12486 430 -12470
rect 383 -12501 437 -12486
rect 123 -13121 167 -12610
rect 169 -12517 178 -12501
rect 371 -12517 437 -12501
rect 169 -12551 437 -12517
rect 169 -12998 178 -12551
rect 371 -12598 437 -12551
rect 505 -12501 516 -12490
rect 517 -12501 559 -12413
rect 560 -12501 571 -12490
rect 383 -12986 425 -12598
rect 391 -12998 425 -12986
rect 169 -13045 179 -12998
rect 355 -13045 425 -12998
rect 169 -13079 425 -13045
rect 169 -13095 179 -13079
rect 357 -13085 367 -13079
rect 169 -13121 178 -13095
rect 385 -13113 425 -13079
rect 391 -13121 425 -13113
rect 94 -13129 199 -13121
rect 382 -13129 425 -13121
rect 505 -12814 571 -12501
rect 1124 -12796 2827 -12301
rect 3191 -12394 5718 -12161
rect 3191 -12488 5784 -12394
rect 3191 -12796 5836 -12488
rect 1124 -12814 5836 -12796
rect 505 -13129 5836 -12814
rect 6434 -12954 6579 -12943
rect 6434 -12988 6542 -12954
rect 6434 -13000 6579 -12988
rect 6434 -13059 6492 -13000
rect -25 -13215 5836 -13129
rect -11 -13223 33 -13215
rect 87 -13217 5836 -13215
rect -11 -13228 70 -13223
rect -11 -13275 33 -13228
rect 111 -13229 5836 -13217
rect -11 -13349 34 -13275
rect 123 -13342 167 -13229
rect 169 -13342 178 -13229
rect 318 -13230 5836 -13229
rect 5843 -13230 5890 -13095
rect 318 -13251 5784 -13230
rect 326 -13257 5784 -13251
rect 324 -13270 5784 -13257
rect 318 -13283 5784 -13270
rect 281 -13288 5784 -13283
rect 5790 -13242 5824 -13230
rect 5790 -13288 5835 -13242
rect 5855 -13288 5889 -13230
rect 281 -13297 5889 -13288
rect 318 -13311 5889 -13297
rect 281 -13317 5889 -13311
rect 123 -13349 178 -13342
rect 180 -13349 5889 -13317
rect -58 -14003 5889 -13349
rect 6368 -13742 6492 -13059
rect 6731 -13132 6822 -13114
rect 6759 -13160 6850 -13142
rect 6568 -13742 6579 -13173
rect 6368 -13800 6884 -13742
rect 6368 -13895 6503 -13800
rect 6568 -13895 6579 -13800
rect 6580 -13858 6614 -13800
rect 6838 -13845 6872 -13800
rect 5977 -13946 6293 -13895
rect 5912 -13953 6293 -13946
rect -58 -14032 5900 -14003
rect 5903 -14032 5912 -13953
rect 5977 -14032 5986 -13953
rect 5989 -14011 6023 -13953
rect 6247 -14007 6281 -13953
rect 5989 -14032 6029 -14011
rect -58 -14113 6029 -14032
rect 6050 -14045 6057 -14039
rect 6230 -14045 6281 -14007
rect 6046 -14079 6057 -14045
rect 6062 -14079 6281 -14045
rect 6050 -14085 6057 -14079
rect -58 -14129 6028 -14113
rect 6235 -14117 6246 -14079
rect -58 -14465 6034 -14129
rect -47 -14552 6034 -14465
rect -47 -14638 5900 -14552
rect 5903 -14638 5934 -14552
rect -47 -14650 5934 -14638
rect 5977 -14578 5986 -14552
rect 5989 -14578 6034 -14552
rect -47 -14724 5912 -14650
rect 5977 -14705 6034 -14578
rect 5977 -14717 5989 -14705
rect -47 -14758 5921 -14724
rect -47 -14788 5912 -14758
rect 5988 -14788 5989 -14717
rect -47 -14816 5900 -14788
rect -47 -14819 5784 -14816
rect 5801 -14819 5835 -14816
rect 5855 -14819 5900 -14816
rect -47 -14853 5799 -14819
rect 5801 -14853 5900 -14819
rect 5906 -14853 5943 -14819
rect -47 -14858 5784 -14853
rect -47 -14874 5789 -14858
rect 5801 -14874 5835 -14853
rect 5855 -14874 5900 -14853
rect -47 -14912 5784 -14874
rect 5789 -14912 5900 -14874
rect 6000 -14881 6034 -14705
rect 6035 -14717 6045 -14118
rect 6247 -14129 6281 -14079
rect 6247 -14705 6292 -14129
rect 6035 -14755 6046 -14717
rect 6219 -14721 6257 -14717
rect 6258 -14721 6292 -14705
rect 6219 -14755 6292 -14721
rect 6035 -14789 6292 -14755
rect 6035 -14805 6046 -14789
rect 6224 -14795 6231 -14789
rect 6252 -14823 6292 -14789
rect 6258 -14881 6292 -14823
rect 6295 -14881 6304 -14117
rect 5988 -14893 6304 -14881
rect -47 -14928 5789 -14912
rect -47 -15249 5784 -14928
rect 5798 -14946 5835 -14912
rect 5866 -14939 5931 -14912
rect 5951 -14927 5965 -14893
rect 5966 -14927 6304 -14893
rect 6319 -14927 6326 -14893
rect 5988 -14939 6304 -14927
rect 5866 -14946 5962 -14939
rect -78 -15295 5784 -15249
rect 1171 -15348 1218 -15295
rect 2743 -15301 5784 -15295
rect 2124 -15313 5784 -15301
rect 1279 -15347 5784 -15313
rect 2743 -15390 5784 -15347
rect 3191 -15395 5784 -15390
rect 40 -15603 88 -15569
rect 136 -15603 184 -15569
rect 232 -15603 280 -15569
rect 328 -15603 376 -15569
rect 424 -15603 472 -15569
rect 501 -15603 503 -15569
rect 555 -15646 557 -15612
rect 586 -15646 634 -15612
rect 682 -15646 730 -15612
rect 778 -15646 826 -15612
rect 874 -15646 922 -15612
rect 970 -15646 1018 -15612
rect 1066 -15646 1114 -15612
rect 1162 -15646 1210 -15612
rect 1239 -15646 1241 -15612
rect 142 -15665 156 -15657
rect 219 -15665 231 -15649
rect 253 -15657 265 -15649
rect 307 -15657 317 -15649
rect 242 -15665 265 -15657
rect 298 -15665 317 -15657
rect 33 -15699 81 -15665
rect 97 -15699 156 -15665
rect 177 -15699 231 -15665
rect 142 -15748 156 -15737
rect 97 -15782 156 -15748
rect 219 -15791 231 -15699
rect 253 -15699 317 -15665
rect 253 -15737 265 -15699
rect 307 -15737 317 -15699
rect 242 -15748 265 -15737
rect 298 -15748 317 -15737
rect 253 -15782 317 -15748
rect 253 -15791 265 -15782
rect 307 -15791 317 -15782
rect 341 -15665 351 -15649
rect 398 -15665 412 -15657
rect 341 -15699 395 -15665
rect 409 -15699 467 -15665
rect 1293 -15689 1295 -15655
rect 1324 -15689 1372 -15655
rect 1420 -15689 1468 -15655
rect 1516 -15689 1564 -15655
rect 1593 -15689 1595 -15655
rect 341 -15791 351 -15699
rect 1117 -15708 1129 -15692
rect 1151 -15700 1163 -15692
rect 1140 -15708 1163 -15700
rect 398 -15748 412 -15737
rect 577 -15742 625 -15708
rect 649 -15742 697 -15708
rect 721 -15742 769 -15708
rect 865 -15742 913 -15708
rect 937 -15742 1057 -15708
rect 1081 -15742 1129 -15708
rect 409 -15782 457 -15748
rect -57 -16023 489 -15791
rect 974 -15825 1022 -15791
rect 1117 -15834 1129 -15742
rect 1151 -15742 1199 -15708
rect 1647 -15732 1649 -15698
rect 1678 -15732 1726 -15698
rect 1774 -15732 1822 -15698
rect 1870 -15732 1918 -15698
rect 1947 -15732 1949 -15698
rect 3220 -15710 5784 -15395
rect 5789 -15616 5847 -14946
rect 5800 -15674 5847 -15616
rect 1151 -15780 1163 -15742
rect 1390 -15751 1404 -15743
rect 1490 -15751 1504 -15743
rect 1140 -15791 1163 -15780
rect 1317 -15785 1437 -15751
rect 1501 -15785 1549 -15751
rect 2001 -15775 2003 -15741
rect 2032 -15775 2080 -15741
rect 2128 -15775 2176 -15741
rect 2224 -15775 2272 -15741
rect 2320 -15775 2368 -15741
rect 2416 -15775 2464 -15741
rect 2493 -15775 2495 -15741
rect 3220 -15784 5718 -15710
rect 5854 -15718 5901 -14946
rect 5988 -15020 6036 -14939
rect 6368 -15004 6491 -13895
rect 6580 -13960 6620 -13858
rect 6641 -13892 6648 -13886
rect 6821 -13892 6872 -13845
rect 6637 -13926 6648 -13892
rect 6653 -13926 6872 -13892
rect 6641 -13932 6648 -13926
rect 6580 -13985 6614 -13960
rect 6826 -13973 6837 -13926
rect 6580 -14761 6625 -13985
rect 6591 -14946 6625 -14761
rect 6626 -14773 6636 -13974
rect 6838 -13985 6872 -13926
rect 6972 -13850 7006 -13050
rect 6838 -14761 6883 -13985
rect 6849 -14773 6883 -14761
rect 6626 -14820 6637 -14773
rect 6693 -14800 6759 -14786
rect 6665 -14820 6759 -14814
rect 6810 -14820 6883 -14773
rect 6626 -14854 6883 -14820
rect 6626 -14870 6637 -14854
rect 6849 -14946 6883 -14854
rect 6972 -14896 7017 -13850
rect 6579 -14958 6895 -14946
rect 6557 -14992 6895 -14958
rect 6910 -14992 6917 -14958
rect 6579 -15004 6895 -14992
rect 6368 -15070 6503 -15004
rect 6379 -15718 6503 -15070
rect 6579 -15573 6590 -15004
rect 6693 -15600 6759 -15586
rect 6665 -15628 6759 -15614
rect 6983 -15696 7017 -14896
rect 5854 -15739 6503 -15718
rect 6379 -15775 6492 -15739
rect 1151 -15825 1199 -15791
rect 1744 -15794 1758 -15786
rect 1844 -15794 1858 -15786
rect 1151 -15834 1163 -15825
rect 1390 -15834 1404 -15823
rect 1490 -15834 1504 -15823
rect 1671 -15828 1791 -15794
rect 1855 -15828 1903 -15794
rect 2547 -15818 2549 -15784
rect 2578 -15818 2626 -15784
rect 2674 -15818 2722 -15784
rect 2770 -15818 2818 -15784
rect 2866 -15818 2914 -15784
rect 2962 -15818 3010 -15784
rect 3058 -15818 3106 -15784
rect 3154 -15818 5718 -15784
rect 6445 -15793 6492 -15775
rect 162 -16063 210 -16029
rect 219 -16077 226 -16023
rect 36 -16090 226 -16077
rect 253 -16077 260 -16023
rect 284 -16077 298 -16023
rect 404 -16045 416 -16029
rect 459 -16045 489 -16023
rect 253 -16095 325 -16077
rect 284 -16111 298 -16095
rect 370 -16111 382 -16061
rect 404 -16077 462 -16045
rect 627 -16066 1227 -15834
rect 1345 -15868 1404 -15834
rect 1501 -15868 1549 -15834
rect 2134 -15837 2148 -15829
rect 2211 -15837 2223 -15821
rect 2245 -15829 2257 -15821
rect 2299 -15829 2309 -15821
rect 2234 -15837 2257 -15829
rect 2290 -15837 2309 -15829
rect 1744 -15877 1758 -15866
rect 1844 -15877 1858 -15866
rect 2025 -15871 2073 -15837
rect 2089 -15871 2148 -15837
rect 2169 -15871 2223 -15837
rect 1365 -15918 1581 -15877
rect 1699 -15911 1758 -15877
rect 1855 -15911 1903 -15877
rect 1345 -15952 1581 -15918
rect 2134 -15920 2148 -15909
rect 1365 -16001 1581 -15952
rect 1719 -15961 1935 -15920
rect 2089 -15954 2148 -15920
rect 1699 -15995 1935 -15961
rect 2211 -15963 2223 -15871
rect 2245 -15871 2309 -15837
rect 2245 -15909 2257 -15871
rect 2299 -15909 2309 -15871
rect 2234 -15920 2257 -15909
rect 2290 -15920 2309 -15909
rect 2245 -15954 2309 -15920
rect 2245 -15963 2257 -15954
rect 2299 -15963 2309 -15954
rect 2333 -15837 2343 -15821
rect 2390 -15837 2404 -15829
rect 2333 -15871 2387 -15837
rect 2401 -15871 2459 -15837
rect 2333 -15963 2343 -15871
rect 3109 -15880 3121 -15864
rect 3143 -15872 3155 -15864
rect 3220 -15870 5718 -15818
rect 3132 -15880 3155 -15872
rect 2390 -15920 2404 -15909
rect 2569 -15914 2617 -15880
rect 2641 -15914 2689 -15880
rect 2713 -15914 2761 -15880
rect 2857 -15914 2905 -15880
rect 2929 -15914 3049 -15880
rect 3073 -15914 3121 -15880
rect 2401 -15954 2449 -15920
rect 1345 -16035 1581 -16001
rect 404 -16095 478 -16077
rect 70 -16113 530 -16111
rect 59 -16129 530 -16113
rect 59 -16145 481 -16129
rect 485 -16145 530 -16129
rect 546 -16145 561 -16111
rect 59 -16173 523 -16145
rect 59 -16191 481 -16173
rect 580 -16179 595 -16077
rect 615 -16124 663 -16090
rect 664 -16124 676 -16074
rect 664 -16154 682 -16124
rect 698 -16154 710 -16066
rect 734 -16095 752 -16066
rect 1060 -16082 1108 -16066
rect 734 -16154 746 -16095
rect 780 -16098 794 -16095
rect 1117 -16098 1124 -16066
rect 768 -16154 794 -16098
rect 796 -16146 844 -16112
rect 1151 -16132 1158 -16066
rect 1197 -16088 1227 -16066
rect 1365 -16109 1581 -16035
rect 1719 -16044 1935 -15995
rect 1699 -16078 1935 -16044
rect 839 -16154 874 -16146
rect 616 -16158 980 -16154
rect 615 -16160 980 -16158
rect 1029 -16160 1172 -16154
rect 1223 -16160 1268 -16154
rect 615 -16184 1268 -16160
rect 1284 -16161 1299 -16154
rect 1318 -16161 1333 -16120
rect 1410 -16149 1458 -16115
rect 517 -16188 1268 -16184
rect 1269 -16163 1354 -16161
rect 1462 -16163 1474 -16109
rect 1269 -16176 1474 -16163
rect 1269 -16188 1354 -16176
rect 517 -16191 1354 -16188
rect 59 -16197 1354 -16191
rect 1496 -16197 1508 -16109
rect 1551 -16131 1619 -16109
rect 1719 -16152 1935 -16078
rect 59 -16199 1526 -16197
rect 59 -16207 481 -16199
rect 517 -16203 1526 -16199
rect 1577 -16203 1622 -16197
rect 517 -16207 1622 -16203
rect 1638 -16204 1653 -16197
rect 1672 -16204 1687 -16163
rect 1764 -16192 1812 -16158
rect 59 -16216 1622 -16207
rect 59 -16234 1237 -16216
rect 1269 -16229 1622 -16216
rect 1311 -16231 1622 -16229
rect 1623 -16206 1708 -16204
rect 1816 -16206 1828 -16152
rect 1623 -16219 1828 -16206
rect 1623 -16231 1708 -16219
rect 59 -16241 1262 -16234
rect 59 -16247 481 -16241
rect 517 -16242 1262 -16241
rect 517 -16247 1237 -16242
rect 59 -16250 1237 -16247
rect 59 -16252 1257 -16250
rect 59 -16253 531 -16252
rect 59 -16275 481 -16253
rect 59 -16281 503 -16275
rect 59 -16287 481 -16281
rect 33 -16290 481 -16287
rect 559 -16284 1257 -16252
rect 559 -16290 1237 -16284
rect 33 -16321 515 -16290
rect 59 -16324 515 -16321
rect 559 -16296 1269 -16290
rect 559 -16318 1237 -16296
rect 559 -16324 1241 -16318
rect 59 -16335 481 -16324
rect 559 -16333 1237 -16324
rect 59 -16349 503 -16335
rect 6 -16357 506 -16349
rect -17 -16378 529 -16357
rect 559 -16367 1257 -16333
rect 559 -16378 1237 -16367
rect -17 -16400 531 -16378
rect 555 -16392 1241 -16378
rect 552 -16400 1237 -16392
rect -17 -16401 1267 -16400
rect -17 -16421 1269 -16401
rect 1277 -16421 1278 -16234
rect 1311 -16240 1708 -16231
rect 1850 -16240 1862 -16152
rect 1905 -16174 1973 -16152
rect 2073 -16195 2481 -15963
rect 2966 -15997 3014 -15963
rect 3109 -16006 3121 -15914
rect 3143 -15914 3191 -15880
rect 3143 -15952 3155 -15914
rect 3132 -15963 3155 -15952
rect 3143 -15997 3191 -15963
rect 3143 -16006 3155 -15997
rect 1311 -16246 1880 -16240
rect 1931 -16246 1976 -16240
rect 1311 -16272 1976 -16246
rect 1992 -16269 2007 -16240
rect 2026 -16249 2041 -16206
rect 2154 -16235 2202 -16201
rect 2211 -16249 2218 -16195
rect 2026 -16262 2218 -16249
rect 2245 -16249 2252 -16195
rect 2276 -16249 2290 -16195
rect 2396 -16217 2408 -16201
rect 2451 -16217 2481 -16195
rect 2245 -16267 2317 -16249
rect 1311 -16277 1633 -16272
rect 1665 -16274 1976 -16272
rect 1985 -16274 2007 -16269
rect 1311 -16285 1634 -16277
rect 1311 -16293 1591 -16285
rect 1311 -16327 1607 -16293
rect 1311 -16333 1591 -16327
rect 1311 -16339 1623 -16333
rect 1311 -16361 1591 -16339
rect 1311 -16367 1595 -16361
rect 1311 -16376 1591 -16367
rect 1311 -16410 1607 -16376
rect 1311 -16421 1591 -16410
rect -17 -16443 1278 -16421
rect 1293 -16435 1595 -16421
rect 1290 -16443 1591 -16435
rect 3 -16449 70 -16443
rect 146 -16446 203 -16443
rect 3 -16451 88 -16449
rect 146 -16457 214 -16446
rect 280 -16451 483 -16443
rect 280 -16454 297 -16451
rect 79 -16471 146 -16457
rect 158 -16491 214 -16457
rect 236 -16465 297 -16454
rect 303 -16457 370 -16451
rect 247 -16499 297 -16465
rect 236 -16524 297 -16499
rect 176 -16571 297 -16524
rect 223 -16582 297 -16571
rect 314 -16491 370 -16457
rect 392 -16465 448 -16454
rect 459 -16457 470 -16451
rect 495 -16457 1621 -16443
rect 314 -16582 331 -16491
rect 403 -16499 448 -16465
rect 470 -16464 1621 -16457
rect 1631 -16464 1634 -16285
rect 1665 -16320 1987 -16274
rect 2276 -16283 2290 -16267
rect 2362 -16283 2374 -16233
rect 2396 -16249 2454 -16217
rect 2619 -16238 3191 -16006
rect 3202 -16172 3203 -15872
rect 3220 -15904 5736 -15870
rect 5784 -15904 5832 -15870
rect 5880 -15904 5928 -15870
rect 5976 -15904 6024 -15870
rect 6072 -15904 6120 -15870
rect 6168 -15904 6216 -15870
rect 6264 -15904 6312 -15870
rect 6360 -15904 6408 -15870
rect 6456 -15904 6504 -15870
rect 6552 -15904 6600 -15870
rect 6648 -15904 6696 -15870
rect 6744 -15904 6792 -15870
rect 6821 -15904 6823 -15870
rect 3220 -15958 5718 -15904
rect 6875 -15947 6877 -15913
rect 6906 -15947 6954 -15913
rect 7002 -15947 7050 -15913
rect 7098 -15947 7146 -15913
rect 7194 -15947 7242 -15913
rect 7290 -15947 7338 -15913
rect 7386 -15947 7434 -15913
rect 7482 -15947 7530 -15913
rect 7578 -15947 7626 -15913
rect 7655 -15947 7657 -15913
rect 3220 -15966 5725 -15958
rect 5767 -15966 5781 -15958
rect 3220 -16023 5718 -15966
rect 5722 -15972 5781 -15966
rect 5827 -15972 5841 -15950
rect 5721 -16000 5781 -15972
rect 5721 -16006 5769 -16000
rect 5793 -16006 5841 -15972
rect 3220 -16034 5725 -16023
rect 5767 -16034 5781 -16023
rect 3220 -16137 5718 -16034
rect 5722 -16068 5781 -16034
rect 3220 -16148 5725 -16137
rect 5767 -16148 5781 -16137
rect 3220 -16205 5718 -16148
rect 5722 -16182 5781 -16148
rect 3220 -16216 5725 -16205
rect 5767 -16216 5781 -16205
rect 2396 -16267 2470 -16249
rect 2062 -16285 2522 -16283
rect 2051 -16301 2522 -16285
rect 2019 -16308 2041 -16303
rect 1665 -16328 1988 -16320
rect 1665 -16336 1945 -16328
rect 1665 -16370 1961 -16336
rect 1665 -16376 1945 -16370
rect 1665 -16382 1977 -16376
rect 1665 -16404 1945 -16382
rect 1665 -16410 1949 -16404
rect 1665 -16419 1945 -16410
rect 1665 -16453 1961 -16419
rect 1665 -16464 1945 -16453
rect 470 -16486 1634 -16464
rect 1647 -16478 1949 -16464
rect 1644 -16486 1945 -16478
rect 470 -16491 531 -16486
rect 495 -16499 527 -16491
rect 549 -16494 1975 -16486
rect 223 -16605 331 -16582
rect 236 -16655 297 -16605
rect 314 -16637 331 -16605
rect 392 -16537 449 -16499
rect 470 -16507 520 -16499
rect 700 -16517 756 -16494
rect 822 -16534 831 -16494
rect 856 -16517 912 -16494
rect 957 -16508 1012 -16497
rect 392 -16613 453 -16537
rect 465 -16587 487 -16571
rect 465 -16613 520 -16587
rect 533 -16613 536 -16571
rect 567 -16613 570 -16542
rect 392 -16655 581 -16613
rect 120 -16823 581 -16655
rect 676 -16666 721 -16632
rect 676 -16716 721 -16700
rect 725 -16716 753 -16536
rect 856 -16568 865 -16517
rect 968 -16542 1012 -16508
rect 1034 -16500 1101 -16494
rect 1178 -16497 1200 -16494
rect 1034 -16534 1091 -16500
rect 1134 -16508 1200 -16497
rect 1201 -16500 1975 -16494
rect 1034 -16542 1054 -16534
rect 1145 -16542 1200 -16508
rect 759 -16716 787 -16570
rect 799 -16606 810 -16595
rect 795 -16637 810 -16606
rect 795 -16648 804 -16637
rect 792 -16690 810 -16648
rect 829 -16674 838 -16640
rect 841 -16674 852 -16637
rect 857 -16674 902 -16654
rect 829 -16688 902 -16674
rect 795 -16708 804 -16690
rect 795 -16716 823 -16708
rect 829 -16716 857 -16688
rect 956 -16716 1012 -16542
rect 1134 -16543 1200 -16542
rect 1074 -16590 1200 -16543
rect 1121 -16624 1200 -16590
rect 1134 -16660 1200 -16624
rect 1212 -16507 1975 -16500
rect 1985 -16507 1988 -16328
rect 2019 -16499 2022 -16308
rect 2051 -16317 2473 -16301
rect 2477 -16317 2522 -16301
rect 2538 -16317 2553 -16283
rect 2051 -16345 2515 -16317
rect 2051 -16363 2473 -16345
rect 2572 -16351 2587 -16249
rect 2607 -16296 2655 -16262
rect 2656 -16296 2668 -16246
rect 2641 -16326 2676 -16296
rect 2690 -16326 2702 -16238
rect 2726 -16267 2744 -16238
rect 3052 -16254 3100 -16238
rect 2726 -16326 2738 -16267
rect 2772 -16270 2786 -16267
rect 3109 -16270 3116 -16238
rect 2760 -16326 2786 -16270
rect 2788 -16318 2836 -16284
rect 3143 -16304 3150 -16238
rect 3220 -16249 5718 -16216
rect 5722 -16249 5781 -16216
rect 5827 -16249 5841 -16006
rect 3220 -16266 5841 -16249
rect 5861 -15958 5875 -15950
rect 5927 -15958 5941 -15950
rect 5861 -15966 5881 -15958
rect 5923 -15966 5941 -15958
rect 5861 -16023 5875 -15966
rect 5878 -16000 5941 -15966
rect 5927 -16023 5941 -16000
rect 5861 -16034 5881 -16023
rect 5923 -16034 5941 -16023
rect 5861 -16137 5875 -16034
rect 5878 -16068 5941 -16034
rect 5927 -16137 5941 -16068
rect 5861 -16148 5881 -16137
rect 5923 -16148 5941 -16137
rect 5861 -16205 5875 -16148
rect 5878 -16182 5941 -16148
rect 5878 -16205 5926 -16203
rect 5927 -16205 5941 -16182
rect 5861 -16216 5941 -16205
rect 3220 -16283 5718 -16266
rect 5861 -16283 5875 -16216
rect 5878 -16229 5941 -16216
rect 5961 -15972 5975 -15950
rect 6023 -15966 6037 -15958
rect 6079 -15966 6093 -15958
rect 6034 -15972 6093 -15966
rect 6139 -15972 6153 -15950
rect 5961 -16006 6009 -15972
rect 6033 -16000 6093 -15972
rect 6033 -16006 6081 -16000
rect 6105 -16006 6153 -15972
rect 5878 -16250 5951 -16229
rect 5881 -16258 5951 -16250
rect 3220 -16317 5897 -16283
rect 5927 -16292 5941 -16258
rect 5961 -16266 5975 -16006
rect 6023 -16034 6037 -16023
rect 6079 -16034 6093 -16023
rect 6034 -16068 6093 -16034
rect 6023 -16148 6037 -16137
rect 6079 -16148 6093 -16137
rect 6034 -16182 6093 -16148
rect 6023 -16216 6037 -16205
rect 6079 -16216 6093 -16205
rect 6034 -16250 6093 -16216
rect 6139 -16266 6153 -16006
rect 6173 -15958 6187 -15950
rect 6239 -15958 6253 -15950
rect 6173 -15966 6193 -15958
rect 6235 -15966 6253 -15958
rect 6173 -16023 6187 -15966
rect 6190 -16000 6253 -15966
rect 6239 -16023 6253 -16000
rect 6173 -16034 6193 -16023
rect 6235 -16034 6253 -16023
rect 6173 -16137 6187 -16034
rect 6190 -16068 6253 -16034
rect 6239 -16137 6253 -16068
rect 6173 -16148 6193 -16137
rect 6235 -16148 6253 -16137
rect 6173 -16205 6187 -16148
rect 6190 -16182 6253 -16148
rect 6190 -16205 6238 -16203
rect 6239 -16205 6253 -16182
rect 6173 -16216 6253 -16205
rect 2833 -16326 2868 -16318
rect 3220 -16323 5846 -16317
rect 3220 -16326 5841 -16323
rect 2610 -16330 2974 -16326
rect 2607 -16332 2974 -16330
rect 3021 -16332 3166 -16326
rect 3217 -16332 5841 -16326
rect 2607 -16351 5841 -16332
rect 2607 -16356 5734 -16351
rect 2509 -16363 5734 -16356
rect 2051 -16371 5734 -16363
rect 5755 -16371 5826 -16351
rect 5827 -16363 5841 -16351
rect 5861 -16342 5875 -16317
rect 5920 -16342 5941 -16292
rect 5961 -16326 5975 -16322
rect 5985 -16326 6020 -16304
rect 6091 -16326 6126 -16304
rect 6139 -16326 6153 -16322
rect 6173 -16326 6187 -16216
rect 6190 -16250 6253 -16216
rect 6239 -16326 6253 -16250
rect 6273 -15972 6287 -15950
rect 6335 -15966 6349 -15958
rect 6391 -15966 6405 -15958
rect 6346 -15972 6405 -15966
rect 6451 -15972 6465 -15950
rect 6273 -16006 6321 -15972
rect 6345 -16000 6405 -15972
rect 6345 -16006 6393 -16000
rect 6417 -16006 6465 -15972
rect 6273 -16266 6287 -16006
rect 6335 -16034 6349 -16023
rect 6391 -16034 6405 -16023
rect 6346 -16068 6405 -16034
rect 6335 -16148 6349 -16137
rect 6391 -16148 6405 -16137
rect 6346 -16182 6405 -16148
rect 6335 -16216 6349 -16205
rect 6391 -16216 6405 -16205
rect 6346 -16250 6405 -16216
rect 6451 -16266 6465 -16006
rect 6485 -15958 6499 -15950
rect 6551 -15958 6565 -15950
rect 6485 -15966 6505 -15958
rect 6547 -15966 6565 -15958
rect 6485 -16023 6499 -15966
rect 6502 -16000 6565 -15966
rect 6551 -16023 6565 -16000
rect 6485 -16034 6505 -16023
rect 6547 -16034 6565 -16023
rect 6485 -16137 6499 -16034
rect 6502 -16068 6565 -16034
rect 6551 -16137 6565 -16068
rect 6485 -16148 6505 -16137
rect 6547 -16148 6565 -16137
rect 6485 -16205 6499 -16148
rect 6502 -16182 6565 -16148
rect 6502 -16205 6550 -16203
rect 6551 -16205 6565 -16182
rect 6485 -16216 6565 -16205
rect 6283 -16322 6318 -16304
rect 6273 -16326 6318 -16322
rect 6379 -16326 6414 -16304
rect 6451 -16326 6465 -16322
rect 6485 -16326 6499 -16216
rect 6502 -16250 6565 -16216
rect 6551 -16300 6565 -16250
rect 6585 -15972 6599 -15966
rect 6647 -15970 6661 -15959
rect 6658 -15972 6706 -15970
rect 6585 -16006 6642 -15972
rect 6658 -16004 6714 -15972
rect 7709 -15990 7711 -15956
rect 7740 -15990 7788 -15956
rect 7836 -15990 7884 -15956
rect 7932 -15990 7980 -15956
rect 8028 -15990 8076 -15956
rect 8124 -15990 8172 -15956
rect 8220 -15990 8268 -15956
rect 8316 -15990 8364 -15956
rect 8412 -15990 8460 -15956
rect 8508 -15990 8556 -15956
rect 8604 -15990 8652 -15956
rect 8700 -15990 8748 -15956
rect 8796 -15990 8844 -15956
rect 8892 -15990 8940 -15956
rect 8988 -15990 9036 -15956
rect 9084 -15990 9132 -15956
rect 9180 -15990 9228 -15956
rect 9276 -15990 9324 -15956
rect 9372 -15990 9420 -15956
rect 9468 -15990 9516 -15956
rect 9564 -15990 9612 -15956
rect 9660 -15990 9708 -15956
rect 9756 -15990 9804 -15956
rect 9852 -15990 9900 -15956
rect 9948 -15990 9996 -15956
rect 10044 -15990 10092 -15956
rect 10140 -15990 10188 -15956
rect 10236 -15990 10284 -15956
rect 10332 -15990 10380 -15956
rect 10409 -15990 10411 -15956
rect 7151 -16001 7163 -15993
rect 6666 -16006 6714 -16004
rect 6585 -16266 6599 -16006
rect 6988 -16009 7002 -16001
rect 7088 -16009 7102 -16001
rect 7144 -16009 7163 -16001
rect 6647 -16038 6661 -16027
rect 6658 -16072 6706 -16038
rect 6899 -16043 7019 -16009
rect 7099 -16043 7163 -16009
rect 6647 -16144 6661 -16133
rect 6705 -16144 6714 -16072
rect 7151 -16077 7163 -16043
rect 6948 -16081 6991 -16077
rect 7099 -16081 7163 -16077
rect 6948 -16092 7002 -16081
rect 7088 -16092 7163 -16081
rect 6931 -16111 6942 -16099
rect 6943 -16111 7002 -16092
rect 7099 -16111 7163 -16092
rect 7185 -16009 7197 -15993
rect 7244 -16009 7258 -16001
rect 7300 -16009 7314 -16001
rect 7377 -16009 7389 -15993
rect 7411 -16001 7423 -15993
rect 7465 -16001 7475 -15993
rect 7400 -16009 7423 -16001
rect 7456 -16009 7475 -16001
rect 7185 -16043 7239 -16009
rect 7255 -16043 7314 -16009
rect 7335 -16043 7389 -16009
rect 7185 -16111 7197 -16043
rect 7244 -16090 7258 -16079
rect 7300 -16090 7314 -16079
rect 6658 -16178 6714 -16144
rect 6759 -16145 6768 -16111
rect 6790 -16145 6834 -16111
rect 6886 -16145 6930 -16111
rect 6931 -16145 7249 -16111
rect 7255 -16124 7314 -16090
rect 6931 -16173 6946 -16158
rect 7083 -16165 7097 -16157
rect 7151 -16165 7163 -16145
rect 6988 -16173 7002 -16165
rect 6931 -16196 7002 -16173
rect 7083 -16173 7102 -16165
rect 7144 -16173 7163 -16165
rect 7083 -16176 7163 -16173
rect 7049 -16196 7063 -16191
rect 6931 -16199 7063 -16196
rect 6647 -16212 6661 -16201
rect 6892 -16207 6902 -16199
rect 6943 -16207 7063 -16199
rect 6658 -16246 6706 -16212
rect 6783 -16241 6827 -16207
rect 6847 -16241 6902 -16207
rect 6927 -16210 7002 -16207
rect 6927 -16241 6971 -16210
rect 7003 -16241 7063 -16207
rect 6932 -16259 7002 -16248
rect 6943 -16279 7002 -16259
rect 7049 -16279 7063 -16241
rect 6847 -16324 6891 -16290
rect 6892 -16324 6902 -16279
rect 6943 -16290 7063 -16279
rect 6943 -16293 7002 -16290
rect 7003 -16301 7063 -16290
rect 5954 -16342 6637 -16326
rect 5861 -16360 6782 -16342
rect 6969 -16347 6977 -16309
rect 7002 -16347 7063 -16301
rect 7083 -16207 7097 -16176
rect 7099 -16191 7163 -16176
rect 7185 -16191 7197 -16145
rect 7377 -16154 7389 -16043
rect 7411 -16043 7475 -16009
rect 7411 -16081 7423 -16043
rect 7465 -16081 7475 -16043
rect 7400 -16092 7423 -16081
rect 7456 -16092 7475 -16081
rect 7411 -16126 7475 -16092
rect 7411 -16154 7423 -16126
rect 7465 -16142 7475 -16126
rect 7432 -16154 7475 -16142
rect 7499 -16009 7509 -15993
rect 7556 -16009 7570 -16001
rect 7499 -16043 7553 -16009
rect 7567 -16043 7625 -16009
rect 10463 -16033 10465 -15999
rect 10494 -16033 10542 -15999
rect 10590 -16033 10638 -15999
rect 10686 -16033 10734 -15999
rect 10782 -16033 10830 -15999
rect 10878 -16033 10926 -15999
rect 10974 -16033 11022 -15999
rect 11070 -16033 11118 -15999
rect 11166 -16033 11214 -15999
rect 11243 -16033 11245 -15999
rect 7499 -16154 7509 -16043
rect 7955 -16044 7969 -16036
rect 7795 -16056 7809 -16045
rect 7895 -16052 7909 -16044
rect 7951 -16052 7969 -16044
rect 7750 -16058 7809 -16056
rect 7556 -16090 7570 -16079
rect 7734 -16090 7854 -16058
rect 7906 -16086 7969 -16052
rect 7567 -16124 7615 -16090
rect 7734 -16092 7782 -16090
rect 7806 -16092 7854 -16090
rect 7955 -16109 7969 -16086
rect 7795 -16120 7809 -16113
rect 7895 -16120 7909 -16109
rect 7951 -16120 7969 -16109
rect 7537 -16154 7572 -16139
rect 7750 -16154 7809 -16120
rect 7906 -16154 7969 -16120
rect 7989 -16058 8003 -16036
rect 8051 -16052 8065 -16044
rect 8107 -16052 8121 -16044
rect 8062 -16058 8121 -16052
rect 8167 -16058 8181 -16036
rect 7989 -16092 8037 -16058
rect 8061 -16086 8121 -16058
rect 8061 -16092 8109 -16086
rect 8133 -16092 8181 -16058
rect 7989 -16120 8003 -16092
rect 8051 -16120 8065 -16109
rect 8107 -16120 8121 -16109
rect 7305 -16162 7668 -16154
rect 7244 -16173 7258 -16162
rect 7300 -16173 7668 -16162
rect 7255 -16188 7668 -16173
rect 7720 -16188 7987 -16154
rect 7099 -16196 7158 -16191
rect 7099 -16207 7214 -16196
rect 7255 -16207 7314 -16188
rect 7083 -16210 7158 -16207
rect 7083 -16241 7141 -16210
rect 7159 -16241 7214 -16207
rect 7083 -16248 7097 -16241
rect 7083 -16259 7158 -16248
rect 7244 -16254 7258 -16243
rect 7300 -16254 7314 -16243
rect 7377 -16244 7389 -16188
rect 7411 -16210 7475 -16188
rect 7411 -16244 7423 -16210
rect 7465 -16244 7475 -16210
rect 7499 -16244 7509 -16188
rect 7567 -16207 7615 -16188
rect 7790 -16219 7795 -16216
rect 7790 -16230 7809 -16219
rect 7750 -16234 7809 -16230
rect 7889 -16234 7909 -16200
rect 7955 -16223 7969 -16188
rect 7951 -16234 7969 -16223
rect 7400 -16250 7414 -16248
rect 7083 -16347 7097 -16259
rect 7099 -16279 7158 -16259
rect 7099 -16290 7214 -16279
rect 7255 -16288 7314 -16254
rect 7327 -16284 7371 -16250
rect 7399 -16259 7443 -16250
rect 7456 -16259 7470 -16248
rect 7399 -16284 7470 -16259
rect 7471 -16284 7515 -16250
rect 7556 -16254 7570 -16243
rect 7734 -16250 7809 -16234
rect 7855 -16250 7875 -16234
rect 7615 -16254 7659 -16250
rect 7567 -16284 7659 -16254
rect 7687 -16264 7809 -16250
rect 7687 -16284 7803 -16264
rect 7831 -16284 7875 -16250
rect 7099 -16293 7158 -16290
rect 7159 -16301 7214 -16290
rect 7411 -16293 7470 -16284
rect 7567 -16288 7615 -16284
rect 7790 -16298 7809 -16287
rect 7158 -16347 7215 -16301
rect 7750 -16332 7809 -16298
rect 5861 -16363 6504 -16360
rect 5863 -16371 6504 -16363
rect 2051 -16379 2473 -16371
rect 2509 -16372 6504 -16371
rect 2509 -16379 5734 -16372
rect 5755 -16379 6504 -16372
rect 2051 -16384 5734 -16379
rect 5744 -16384 6504 -16379
rect 6546 -16384 6782 -16360
rect 6869 -16374 7063 -16347
rect 2051 -16413 6782 -16384
rect 6847 -16394 7063 -16374
rect 7073 -16394 7215 -16347
rect 7724 -16367 7768 -16333
rect 7795 -16386 7800 -16344
rect 6847 -16408 6891 -16394
rect 6892 -16408 6902 -16394
rect 2051 -16419 2473 -16413
rect 2509 -16419 6782 -16413
rect 2051 -16424 6782 -16419
rect 2051 -16425 2523 -16424
rect 2051 -16447 2473 -16425
rect 2034 -16453 2495 -16447
rect 2051 -16459 2473 -16453
rect 2025 -16462 2473 -16459
rect 2025 -16493 2507 -16462
rect 2051 -16496 2507 -16493
rect 2051 -16507 2473 -16496
rect 2551 -16499 6782 -16424
rect 6896 -16446 6902 -16408
rect 6916 -16419 7236 -16394
rect 7256 -16419 7304 -16394
rect 7324 -16419 7372 -16394
rect 6916 -16428 7377 -16419
rect 7392 -16428 7440 -16394
rect 7548 -16416 7570 -16394
rect 6847 -16491 6891 -16457
rect 6892 -16491 6902 -16446
rect 6969 -16461 6977 -16428
rect 7002 -16446 7063 -16428
rect 6992 -16457 7063 -16446
rect 7002 -16461 7063 -16457
rect 7091 -16461 7097 -16428
rect 7158 -16446 7377 -16428
rect 7148 -16457 7377 -16446
rect 7158 -16458 7377 -16457
rect 7511 -16434 7623 -16416
rect 7158 -16461 7444 -16458
rect 7511 -16461 7526 -16434
rect 7545 -16458 7589 -16450
rect 7590 -16458 7612 -16434
rect 7544 -16461 7589 -16458
rect 7615 -16461 7623 -16434
rect 7712 -16458 7715 -16417
rect 7724 -16451 7768 -16417
rect 1212 -16529 1988 -16507
rect 2001 -16521 2495 -16507
rect 1998 -16529 2473 -16521
rect 1212 -16534 1278 -16529
rect 1212 -16542 1269 -16534
rect 1212 -16550 1262 -16542
rect 1212 -16660 1234 -16550
rect 1271 -16660 1278 -16534
rect 1287 -16537 1575 -16529
rect 1305 -16660 1312 -16537
rect 1394 -16543 1462 -16537
rect 1327 -16557 1394 -16543
rect 1406 -16577 1462 -16543
rect 1484 -16551 1540 -16540
rect 1551 -16543 1562 -16537
rect 1587 -16543 2521 -16529
rect 1495 -16585 1540 -16551
rect 1562 -16550 2521 -16543
rect 2551 -16550 6809 -16499
rect 1562 -16572 2523 -16550
rect 2547 -16564 6809 -16550
rect 2544 -16565 6809 -16564
rect 6905 -16565 7653 -16461
rect 7794 -16470 7800 -16386
rect 7855 -16470 7875 -16284
rect 7889 -16268 7969 -16234
rect 7889 -16284 7945 -16268
rect 7951 -16284 7969 -16268
rect 7889 -16289 7909 -16284
rect 7889 -16291 7954 -16289
rect 7955 -16291 7969 -16284
rect 7889 -16336 7969 -16291
rect 7889 -16344 7945 -16336
rect 7951 -16344 7969 -16336
rect 7889 -16367 7969 -16344
rect 7989 -16222 8021 -16120
rect 8062 -16154 8121 -16120
rect 8167 -16197 8181 -16092
rect 8201 -16044 8215 -16036
rect 8267 -16044 8281 -16036
rect 8201 -16052 8221 -16044
rect 8263 -16052 8281 -16044
rect 8201 -16109 8215 -16052
rect 8218 -16086 8281 -16052
rect 8267 -16109 8281 -16086
rect 8201 -16120 8221 -16109
rect 8263 -16120 8281 -16109
rect 8201 -16197 8215 -16120
rect 8218 -16154 8281 -16120
rect 8267 -16197 8281 -16154
rect 8301 -16058 8315 -16036
rect 8363 -16052 8377 -16044
rect 8419 -16052 8433 -16044
rect 8374 -16058 8433 -16052
rect 8479 -16058 8493 -16036
rect 8301 -16092 8349 -16058
rect 8373 -16086 8433 -16058
rect 8373 -16092 8421 -16086
rect 8445 -16092 8493 -16058
rect 8301 -16197 8315 -16092
rect 8363 -16120 8377 -16109
rect 8419 -16120 8433 -16109
rect 8374 -16154 8433 -16120
rect 7989 -16352 8003 -16222
rect 8043 -16231 8341 -16197
rect 8051 -16234 8065 -16231
rect 8107 -16234 8121 -16231
rect 8062 -16268 8121 -16234
rect 8167 -16277 8181 -16231
rect 8201 -16234 8221 -16231
rect 8263 -16234 8281 -16231
rect 8201 -16243 8215 -16234
rect 8218 -16243 8281 -16234
rect 8201 -16268 8281 -16243
rect 8051 -16302 8065 -16291
rect 8107 -16293 8150 -16282
rect 8167 -16293 8189 -16277
rect 8067 -16302 8189 -16293
rect 8062 -16327 8189 -16302
rect 8062 -16336 8121 -16327
rect 7889 -16386 7909 -16367
rect 7931 -16370 7969 -16367
rect 7951 -16386 7969 -16370
rect 7889 -16428 7969 -16386
rect 8083 -16376 8098 -16371
rect 8107 -16376 8150 -16344
rect 8083 -16377 8150 -16376
rect 8167 -16377 8189 -16327
rect 8201 -16285 8250 -16268
rect 8267 -16277 8281 -16268
rect 8301 -16277 8315 -16231
rect 8363 -16234 8377 -16223
rect 8419 -16234 8433 -16223
rect 8374 -16240 8433 -16234
rect 8479 -16240 8493 -16092
rect 8513 -16044 8527 -16036
rect 8579 -16044 8593 -16036
rect 8513 -16052 8533 -16044
rect 8575 -16052 8593 -16044
rect 8513 -16109 8527 -16052
rect 8530 -16086 8593 -16052
rect 8579 -16109 8593 -16086
rect 8513 -16120 8533 -16109
rect 8575 -16120 8593 -16109
rect 8513 -16223 8527 -16120
rect 8530 -16154 8593 -16120
rect 8579 -16223 8593 -16154
rect 8513 -16234 8533 -16223
rect 8575 -16234 8593 -16223
rect 8513 -16240 8527 -16234
rect 8530 -16240 8593 -16234
rect 8613 -16058 8627 -16036
rect 8675 -16052 8689 -16044
rect 8731 -16052 8745 -16044
rect 8686 -16058 8745 -16052
rect 8791 -16058 8805 -16036
rect 8613 -16092 8661 -16058
rect 8685 -16086 8745 -16058
rect 8685 -16092 8733 -16086
rect 8757 -16092 8805 -16058
rect 8613 -16240 8627 -16092
rect 8675 -16120 8689 -16109
rect 8731 -16120 8745 -16109
rect 8686 -16154 8745 -16120
rect 8675 -16234 8689 -16223
rect 8731 -16234 8745 -16223
rect 8686 -16240 8745 -16234
rect 8374 -16268 8745 -16240
rect 8397 -16280 8695 -16268
rect 8201 -16289 8223 -16285
rect 8240 -16289 8250 -16285
rect 8263 -16289 8306 -16282
rect 8479 -16289 8493 -16280
rect 8513 -16283 8527 -16280
rect 8579 -16283 8593 -16280
rect 8513 -16289 8593 -16283
rect 8613 -16289 8627 -16280
rect 8791 -16283 8805 -16092
rect 8825 -16044 8839 -16036
rect 8891 -16044 8905 -16036
rect 8825 -16052 8845 -16044
rect 8887 -16052 8905 -16044
rect 8825 -16109 8839 -16052
rect 8842 -16086 8905 -16052
rect 8891 -16109 8905 -16086
rect 8825 -16120 8845 -16109
rect 8887 -16120 8905 -16109
rect 8825 -16223 8839 -16120
rect 8842 -16154 8905 -16120
rect 8891 -16223 8905 -16154
rect 8825 -16234 8845 -16223
rect 8887 -16234 8905 -16223
rect 8825 -16283 8839 -16234
rect 8842 -16268 8905 -16234
rect 8925 -16058 8939 -16036
rect 8987 -16052 9001 -16044
rect 9043 -16052 9057 -16044
rect 8998 -16058 9057 -16052
rect 9103 -16058 9117 -16036
rect 8925 -16092 8973 -16058
rect 8997 -16086 9057 -16058
rect 8997 -16092 9045 -16086
rect 9069 -16092 9117 -16058
rect 8878 -16283 8924 -16268
rect 8925 -16283 8939 -16092
rect 8987 -16120 9001 -16109
rect 9043 -16120 9057 -16109
rect 8998 -16154 9057 -16120
rect 8987 -16234 9001 -16223
rect 9043 -16234 9057 -16223
rect 8998 -16268 9057 -16234
rect 9103 -16283 9117 -16092
rect 9137 -16044 9151 -16036
rect 9203 -16044 9217 -16036
rect 9137 -16052 9157 -16044
rect 9199 -16052 9217 -16044
rect 9137 -16109 9151 -16052
rect 9154 -16086 9217 -16052
rect 9203 -16109 9217 -16086
rect 9137 -16120 9157 -16109
rect 9199 -16120 9217 -16109
rect 9137 -16223 9151 -16120
rect 9154 -16154 9217 -16120
rect 9203 -16223 9217 -16154
rect 9137 -16234 9157 -16223
rect 9199 -16234 9217 -16223
rect 9137 -16283 9151 -16234
rect 9154 -16268 9217 -16234
rect 9237 -16058 9251 -16036
rect 9299 -16052 9313 -16044
rect 9355 -16052 9369 -16044
rect 9310 -16058 9369 -16052
rect 9415 -16058 9429 -16036
rect 9237 -16092 9285 -16058
rect 9309 -16086 9369 -16058
rect 9309 -16092 9357 -16086
rect 9381 -16092 9429 -16058
rect 9166 -16283 9236 -16268
rect 9237 -16283 9251 -16092
rect 9299 -16120 9313 -16109
rect 9355 -16120 9369 -16109
rect 9310 -16154 9369 -16120
rect 9299 -16234 9313 -16223
rect 9355 -16234 9369 -16223
rect 9310 -16268 9369 -16234
rect 8201 -16327 8306 -16289
rect 8369 -16291 8723 -16289
rect 8363 -16302 8723 -16291
rect 8731 -16302 8745 -16291
rect 8369 -16308 8745 -16302
rect 8201 -16336 8277 -16327
rect 8374 -16336 8433 -16308
rect 8479 -16320 8493 -16308
rect 8513 -16320 8593 -16308
rect 8613 -16320 8627 -16308
rect 8438 -16336 8504 -16325
rect 8519 -16328 8589 -16320
rect 8530 -16336 8589 -16328
rect 8594 -16336 8660 -16325
rect 8686 -16329 8745 -16308
rect 8751 -16317 9241 -16283
rect 9299 -16302 9313 -16291
rect 9355 -16302 9369 -16291
rect 8791 -16329 8805 -16317
rect 8686 -16336 8805 -16329
rect 8201 -16377 8223 -16336
rect 8263 -16344 8292 -16336
rect 8240 -16376 8250 -16365
rect 8263 -16376 8307 -16344
rect 8421 -16370 8537 -16336
rect 8605 -16344 8660 -16336
rect 7989 -16428 8003 -16408
rect 8005 -16428 8053 -16424
rect 8083 -16428 8223 -16377
rect 8251 -16386 8307 -16376
rect 7889 -16458 8223 -16428
rect 8250 -16428 8307 -16386
rect 8437 -16424 8504 -16370
rect 8604 -16408 8661 -16344
rect 8735 -16351 8805 -16336
rect 8825 -16323 8839 -16317
rect 8842 -16323 8994 -16317
rect 8825 -16329 8994 -16323
rect 8998 -16323 9151 -16317
rect 9154 -16323 9217 -16317
rect 8998 -16329 9217 -16323
rect 8825 -16351 8839 -16329
rect 8842 -16344 9151 -16329
rect 9154 -16336 9217 -16329
rect 9157 -16344 9199 -16336
rect 8842 -16345 8845 -16344
rect 8884 -16351 8887 -16345
rect 8891 -16351 8905 -16344
rect 8925 -16351 9117 -16344
rect 9137 -16351 9151 -16344
rect 9203 -16351 9217 -16336
rect 9237 -16351 9251 -16317
rect 9310 -16326 9369 -16302
rect 9415 -16326 9429 -16092
rect 9449 -16044 9463 -16036
rect 9515 -16044 9529 -16036
rect 9449 -16052 9469 -16044
rect 9511 -16052 9529 -16044
rect 9449 -16109 9463 -16052
rect 9466 -16086 9529 -16052
rect 9515 -16109 9529 -16086
rect 9449 -16120 9469 -16109
rect 9511 -16120 9529 -16109
rect 9449 -16223 9463 -16120
rect 9466 -16154 9529 -16120
rect 9515 -16223 9529 -16154
rect 9449 -16234 9469 -16223
rect 9511 -16234 9529 -16223
rect 9449 -16291 9463 -16234
rect 9466 -16268 9529 -16234
rect 9466 -16291 9514 -16289
rect 9515 -16291 9529 -16268
rect 9449 -16302 9529 -16291
rect 9449 -16326 9463 -16302
rect 9466 -16326 9529 -16302
rect 9549 -16058 9563 -16036
rect 9611 -16052 9625 -16044
rect 9667 -16052 9681 -16044
rect 9622 -16058 9681 -16052
rect 9727 -16058 9741 -16036
rect 9549 -16092 9597 -16058
rect 9621 -16086 9681 -16058
rect 9621 -16092 9669 -16086
rect 9693 -16092 9741 -16058
rect 9549 -16326 9563 -16092
rect 9611 -16120 9625 -16109
rect 9667 -16120 9681 -16109
rect 9622 -16154 9681 -16120
rect 9611 -16234 9625 -16223
rect 9667 -16234 9681 -16223
rect 9622 -16268 9681 -16234
rect 9611 -16302 9625 -16291
rect 9667 -16302 9681 -16291
rect 9622 -16326 9681 -16302
rect 9727 -16326 9741 -16092
rect 9761 -16044 9775 -16036
rect 9827 -16044 9841 -16036
rect 9761 -16052 9781 -16044
rect 9823 -16052 9841 -16044
rect 9761 -16109 9775 -16052
rect 9778 -16086 9841 -16052
rect 9827 -16109 9841 -16086
rect 9761 -16120 9781 -16109
rect 9823 -16120 9841 -16109
rect 9761 -16223 9775 -16120
rect 9778 -16154 9841 -16120
rect 9827 -16223 9841 -16154
rect 9761 -16234 9781 -16223
rect 9823 -16234 9841 -16223
rect 9761 -16291 9775 -16234
rect 9778 -16268 9841 -16234
rect 9778 -16291 9826 -16289
rect 9827 -16291 9841 -16268
rect 9761 -16302 9841 -16291
rect 9761 -16326 9775 -16302
rect 9778 -16326 9841 -16302
rect 9861 -16058 9875 -16036
rect 9923 -16052 9937 -16044
rect 9979 -16052 9993 -16044
rect 9934 -16058 9993 -16052
rect 10039 -16058 10053 -16036
rect 9861 -16092 9909 -16058
rect 9933 -16086 9993 -16058
rect 9933 -16092 9981 -16086
rect 10005 -16092 10053 -16058
rect 9861 -16326 9875 -16092
rect 9923 -16120 9937 -16109
rect 9979 -16120 9993 -16109
rect 9934 -16154 9993 -16120
rect 9923 -16234 9937 -16223
rect 9979 -16234 9993 -16223
rect 9934 -16268 9993 -16234
rect 9923 -16302 9937 -16291
rect 9979 -16302 9993 -16291
rect 9934 -16326 9993 -16302
rect 8735 -16352 9251 -16351
rect 9299 -16336 9993 -16326
rect 9299 -16344 9981 -16336
rect 9299 -16349 9313 -16344
rect 9330 -16349 9470 -16344
rect 9511 -16349 9662 -16344
rect 9667 -16349 9781 -16344
rect 8802 -16357 8930 -16352
rect 8825 -16363 8839 -16357
rect 8769 -16371 8839 -16363
rect 8884 -16371 8887 -16357
rect 8891 -16363 8905 -16357
rect 9040 -16363 9043 -16352
rect 9114 -16357 9241 -16352
rect 9137 -16363 9151 -16357
rect 8891 -16371 8969 -16363
rect 8995 -16371 9055 -16363
rect 8769 -16379 8860 -16371
rect 8884 -16377 8969 -16371
rect 8984 -16377 9055 -16371
rect 9083 -16371 9151 -16363
rect 9203 -16371 9217 -16357
rect 9299 -16360 9324 -16349
rect 9330 -16360 9480 -16349
rect 9500 -16360 9792 -16349
rect 9810 -16360 9950 -16344
rect 9979 -16349 9981 -16344
rect 9968 -16360 9981 -16349
rect 10039 -16352 10053 -16092
rect 10073 -16044 10087 -16036
rect 10139 -16044 10153 -16036
rect 10073 -16052 10093 -16044
rect 10135 -16052 10153 -16044
rect 10073 -16109 10087 -16052
rect 10090 -16086 10153 -16052
rect 10073 -16120 10093 -16109
rect 10139 -16111 10153 -16086
rect 10173 -16058 10187 -16052
rect 10235 -16056 10249 -16045
rect 10246 -16058 10294 -16056
rect 10173 -16092 10230 -16058
rect 10246 -16090 10302 -16058
rect 11297 -16076 11299 -16042
rect 11328 -16076 11376 -16042
rect 11424 -16076 11472 -16042
rect 11520 -16076 11568 -16042
rect 11616 -16076 11664 -16042
rect 11712 -16076 11760 -16042
rect 11808 -16076 11856 -16042
rect 11904 -16076 11952 -16042
rect 12000 -16076 12048 -16042
rect 12096 -16076 12144 -16042
rect 12192 -16076 12240 -16042
rect 12288 -16076 12336 -16042
rect 12384 -16076 12432 -16042
rect 12480 -16076 12528 -16042
rect 12576 -16076 12624 -16042
rect 12672 -16076 12720 -16042
rect 12768 -16076 12816 -16042
rect 12864 -16076 12912 -16042
rect 12960 -16076 13008 -16042
rect 13056 -16076 13104 -16042
rect 13152 -16076 13200 -16042
rect 13248 -16076 13296 -16042
rect 13344 -16076 13392 -16042
rect 13440 -16076 13488 -16042
rect 13536 -16057 13584 -16042
rect 13525 -16076 13584 -16057
rect 13632 -16076 13680 -16042
rect 13681 -16076 13723 -16057
rect 13728 -16076 13776 -16042
rect 13824 -16057 13872 -16042
rect 13920 -16057 13968 -16042
rect 13824 -16076 13991 -16057
rect 13997 -16076 13999 -16042
rect 10254 -16092 10302 -16090
rect 10173 -16111 10187 -16092
rect 10313 -16098 10411 -16077
rect 10739 -16087 10751 -16079
rect 10576 -16095 10590 -16087
rect 10676 -16095 10690 -16087
rect 10732 -16095 10751 -16087
rect 10313 -16111 10439 -16105
rect 10103 -16120 10302 -16111
rect 10073 -16223 10087 -16120
rect 10090 -16145 10302 -16120
rect 10313 -16126 10466 -16111
rect 10326 -16145 10370 -16126
rect 10422 -16145 10466 -16126
rect 10487 -16129 10607 -16095
rect 10687 -16120 10751 -16095
rect 10773 -16095 10785 -16079
rect 10832 -16095 10846 -16087
rect 10888 -16095 10902 -16087
rect 10965 -16095 10977 -16079
rect 10999 -16087 11011 -16079
rect 11053 -16087 11063 -16079
rect 10988 -16095 11011 -16087
rect 11044 -16095 11063 -16087
rect 10773 -16120 10827 -16095
rect 10843 -16120 10902 -16095
rect 10923 -16120 10977 -16095
rect 10999 -16120 11063 -16095
rect 11087 -16095 11097 -16079
rect 13657 -16082 13965 -16077
rect 11144 -16095 11158 -16087
rect 11087 -16120 11141 -16095
rect 11155 -16120 11213 -16095
rect 14051 -16100 14053 -16085
rect 14082 -16100 14130 -16085
rect 13657 -16110 13937 -16105
rect 10518 -16145 10593 -16129
rect 10621 -16141 11245 -16120
rect 11543 -16130 11557 -16122
rect 10090 -16154 10153 -16145
rect 10139 -16191 10153 -16154
rect 10173 -16191 10187 -16145
rect 10246 -16158 10294 -16145
rect 10739 -16148 10751 -16141
rect 10773 -16148 10785 -16141
rect 10965 -16148 10977 -16141
rect 10999 -16148 11011 -16141
rect 11053 -16148 11063 -16141
rect 11087 -16148 11097 -16141
rect 11383 -16142 11397 -16131
rect 11483 -16138 11497 -16130
rect 11539 -16138 11557 -16130
rect 11338 -16144 11397 -16142
rect 10649 -16154 11273 -16148
rect 10287 -16173 10302 -16158
rect 10236 -16196 10302 -16173
rect 10576 -16178 10590 -16167
rect 10180 -16199 10302 -16196
rect 10180 -16207 10246 -16199
rect 10313 -16207 10321 -16191
rect 10336 -16207 10346 -16199
rect 10347 -16207 10355 -16191
rect 10401 -16199 10407 -16191
rect 10073 -16234 10093 -16223
rect 10127 -16234 10171 -16207
rect 10073 -16291 10087 -16234
rect 10090 -16241 10171 -16234
rect 10191 -16219 10246 -16207
rect 10271 -16219 10321 -16207
rect 10191 -16241 10321 -16219
rect 10090 -16268 10149 -16241
rect 10246 -16264 10305 -16241
rect 10180 -16287 10246 -16279
rect 10090 -16291 10138 -16289
rect 10180 -16290 10305 -16287
rect 10073 -16302 10149 -16291
rect 10073 -16314 10087 -16302
rect 10090 -16314 10149 -16302
rect 10073 -16329 10150 -16314
rect 10191 -16324 10305 -16290
rect 9083 -16377 9172 -16371
rect 8884 -16379 9172 -16377
rect 9184 -16379 9217 -16371
rect 8769 -16386 9217 -16379
rect 8775 -16403 8819 -16386
rect 8594 -16419 8661 -16408
rect 8317 -16428 8365 -16424
rect 8430 -16428 8504 -16424
rect 8250 -16449 8504 -16428
rect 7889 -16470 8150 -16458
rect 8167 -16470 8189 -16458
rect 8201 -16470 8223 -16458
rect 8240 -16453 8504 -16449
rect 8604 -16424 8661 -16419
rect 8751 -16409 8819 -16403
rect 8827 -16409 9149 -16386
rect 9150 -16409 9217 -16386
rect 9234 -16408 9241 -16403
rect 9234 -16409 9251 -16408
rect 8751 -16424 9251 -16409
rect 9415 -16416 9429 -16408
rect 9449 -16416 9463 -16374
rect 9299 -16424 9437 -16422
rect 8604 -16428 8677 -16424
rect 8742 -16425 9251 -16424
rect 8742 -16428 8790 -16425
rect 8827 -16428 8894 -16425
rect 8604 -16437 8894 -16428
rect 8941 -16431 9050 -16425
rect 9054 -16431 9149 -16425
rect 8941 -16437 9149 -16431
rect 9150 -16428 9217 -16425
rect 9237 -16428 9251 -16425
rect 9253 -16428 9437 -16424
rect 9465 -16428 9509 -16422
rect 9515 -16428 9529 -16374
rect 9861 -16408 9869 -16406
rect 9895 -16408 9903 -16406
rect 9549 -16428 9563 -16408
rect 9706 -16422 9784 -16414
rect 9830 -16422 9951 -16414
rect 9600 -16424 9653 -16422
rect 9565 -16428 9653 -16424
rect 9672 -16428 9797 -16422
rect 9150 -16437 9797 -16428
rect 8604 -16453 9797 -16437
rect 8240 -16458 8525 -16453
rect 8240 -16460 8504 -16458
rect 8250 -16470 8504 -16460
rect 8604 -16470 8894 -16453
rect 8941 -16456 9797 -16453
rect 9825 -16424 9951 -16422
rect 9825 -16456 9869 -16424
rect 9877 -16428 9951 -16424
rect 9990 -16428 10038 -16424
rect 10039 -16428 10053 -16408
rect 10073 -16428 10087 -16329
rect 10090 -16336 10149 -16329
rect 10246 -16332 10305 -16324
rect 10103 -16357 10178 -16342
rect 10179 -16363 10236 -16344
rect 10179 -16408 10246 -16363
rect 10179 -16428 10236 -16408
rect 9877 -16446 10236 -16428
rect 8941 -16458 9784 -16456
rect 9877 -16458 10246 -16446
rect 8962 -16470 9082 -16458
rect 9140 -16462 9784 -16458
rect 9150 -16470 9784 -16462
rect 9894 -16470 10246 -16458
rect 10313 -16470 10321 -16241
rect 10347 -16241 10391 -16207
rect 10392 -16241 10407 -16199
rect 10336 -16290 10346 -16279
rect 10347 -16290 10355 -16241
rect 10401 -16279 10407 -16241
rect 10347 -16324 10391 -16290
rect 10392 -16324 10407 -16279
rect 10336 -16374 10346 -16363
rect 10347 -16374 10355 -16324
rect 10401 -16363 10407 -16324
rect 10347 -16408 10391 -16374
rect 10392 -16408 10407 -16363
rect 10336 -16457 10346 -16446
rect 10347 -16457 10355 -16408
rect 10401 -16446 10407 -16408
rect 2544 -16572 6703 -16565
rect 6931 -16571 6994 -16565
rect 1562 -16577 1634 -16572
rect 1587 -16580 1634 -16577
rect 1641 -16580 1929 -16572
rect 1587 -16585 1619 -16580
rect 1484 -16593 1541 -16585
rect 1562 -16593 1612 -16585
rect 1484 -16610 1556 -16593
rect 1424 -16657 1556 -16610
rect 1134 -16702 1337 -16660
rect 1471 -16691 1556 -16657
rect 641 -16722 1012 -16716
rect 641 -16731 825 -16722
rect 656 -16734 823 -16731
rect 656 -16768 678 -16734
rect 725 -16768 753 -16734
rect 759 -16768 823 -16734
rect 829 -16756 1012 -16722
rect 829 -16768 857 -16756
rect 934 -16768 1012 -16756
rect 1022 -16768 1337 -16702
rect 1484 -16703 1556 -16691
rect 1557 -16703 1590 -16593
rect 1625 -16703 1634 -16580
rect 1659 -16703 1668 -16580
rect 1748 -16586 1816 -16580
rect 1681 -16600 1748 -16586
rect 1760 -16620 1816 -16586
rect 1838 -16594 1894 -16583
rect 1905 -16586 1916 -16580
rect 1941 -16582 6703 -16572
rect 1941 -16586 6714 -16582
rect 1849 -16628 1894 -16594
rect 1916 -16615 6714 -16586
rect 6912 -16584 6994 -16571
rect 6912 -16605 7002 -16584
rect 7049 -16603 7063 -16565
rect 7083 -16584 7097 -16565
rect 7102 -16584 7653 -16565
rect 7083 -16587 7653 -16584
rect 7083 -16595 7147 -16587
rect 7083 -16603 7097 -16595
rect 1916 -16620 1988 -16615
rect 1941 -16623 1988 -16620
rect 1995 -16623 2475 -16615
rect 2489 -16616 6714 -16615
rect 1941 -16628 1973 -16623
rect 1838 -16636 1895 -16628
rect 1916 -16636 1966 -16628
rect 1838 -16653 1910 -16636
rect 1778 -16700 1910 -16653
rect 1484 -16745 1691 -16703
rect 1825 -16734 1910 -16700
rect 94 -16863 139 -16829
rect 146 -16831 228 -16823
rect 314 -16829 345 -16823
rect 166 -16863 211 -16831
rect 238 -16863 283 -16829
rect 310 -16863 355 -16829
rect 370 -16831 480 -16823
rect 483 -16831 581 -16823
rect 620 -16816 1337 -16768
rect 1372 -16816 1691 -16745
rect 1838 -16746 1910 -16734
rect 1911 -16746 1944 -16636
rect 1979 -16746 1988 -16623
rect 2013 -16746 2022 -16623
rect 2138 -16629 2206 -16623
rect 2272 -16626 2289 -16623
rect 2071 -16643 2138 -16629
rect 2150 -16663 2206 -16629
rect 2228 -16637 2289 -16626
rect 2295 -16629 2362 -16623
rect 2239 -16671 2289 -16637
rect 2228 -16696 2289 -16671
rect 2168 -16743 2289 -16696
rect 1838 -16788 2045 -16746
rect 2215 -16754 2289 -16743
rect 2306 -16663 2362 -16629
rect 2384 -16637 2440 -16626
rect 2451 -16629 2462 -16623
rect 2489 -16629 6703 -16616
rect 2306 -16754 2323 -16663
rect 2395 -16671 2440 -16637
rect 2462 -16658 6703 -16629
rect 6931 -16621 7002 -16605
rect 7099 -16621 7147 -16595
rect 7154 -16608 7653 -16587
rect 7715 -16565 10328 -16470
rect 10347 -16491 10391 -16457
rect 10392 -16491 10407 -16446
rect 10336 -16525 10346 -16496
rect 10347 -16541 10355 -16491
rect 7715 -16608 10053 -16565
rect 7154 -16621 7246 -16608
rect 6931 -16631 7258 -16621
rect 7327 -16629 7470 -16608
rect 7517 -16611 7526 -16608
rect 7551 -16611 7560 -16608
rect 7517 -16616 7560 -16611
rect 7567 -16616 7627 -16608
rect 7749 -16615 7808 -16608
rect 7327 -16631 7456 -16629
rect 6899 -16637 7295 -16631
rect 6899 -16639 6947 -16637
rect 6971 -16639 7019 -16637
rect 2462 -16663 2523 -16658
rect 2489 -16671 2519 -16663
rect 2543 -16666 6703 -16658
rect 2215 -16777 2323 -16754
rect 456 -16833 539 -16831
rect 483 -16866 539 -16833
rect 620 -16843 1691 -16816
rect 620 -16866 1337 -16843
rect 622 -16874 642 -16866
rect 646 -16878 699 -16866
rect 819 -16874 852 -16866
rect 1019 -16870 1116 -16866
rect 1019 -16872 1126 -16870
rect 752 -16878 852 -16874
rect 408 -16879 442 -16878
rect 247 -16895 319 -16891
rect 398 -16895 458 -16891
rect 70 -16929 530 -16925
rect 70 -16939 242 -16929
rect 278 -16939 378 -16929
rect 389 -16939 434 -16929
rect 70 -16959 435 -16939
rect 485 -16959 530 -16929
rect 540 -16959 561 -16925
rect 574 -16992 595 -16891
rect 834 -16895 852 -16878
rect 953 -16906 998 -16872
rect 1019 -16878 1142 -16872
rect 1025 -16906 1070 -16878
rect 1097 -16906 1142 -16878
rect 1178 -16920 1200 -16866
rect 1212 -16878 1337 -16866
rect 1372 -16859 1691 -16843
rect 1726 -16859 2045 -16788
rect 2228 -16827 2289 -16777
rect 2306 -16809 2323 -16777
rect 2384 -16709 2441 -16671
rect 2462 -16679 2512 -16671
rect 2694 -16689 2750 -16666
rect 2816 -16706 2825 -16666
rect 2850 -16689 2906 -16666
rect 2951 -16680 3006 -16669
rect 2384 -16785 2445 -16709
rect 2457 -16759 2479 -16743
rect 2457 -16785 2512 -16759
rect 2527 -16785 2528 -16743
rect 2561 -16785 2562 -16714
rect 2384 -16827 2573 -16785
rect 1212 -16886 1295 -16878
rect 1221 -16909 1295 -16886
rect 1372 -16886 2045 -16859
rect 1372 -16909 1691 -16886
rect 1398 -16915 1476 -16909
rect 1378 -16921 1495 -16915
rect 1034 -16960 1038 -16957
rect 616 -16978 732 -16968
rect 743 -16978 934 -16968
rect 935 -16978 980 -16968
rect 616 -16986 981 -16978
rect 1031 -16986 1172 -16968
rect 616 -17002 1191 -16986
rect 1223 -17002 1299 -16968
rect 1312 -16976 1333 -16934
rect 1378 -16949 1423 -16921
rect 1450 -16949 1495 -16921
rect 1523 -16963 1556 -16909
rect 1557 -16921 1691 -16909
rect 1557 -16929 1649 -16921
rect 1575 -16952 1649 -16929
rect 1726 -16952 2045 -16886
rect 2071 -16921 2083 -16902
rect 2112 -16921 2573 -16827
rect 2670 -16838 2715 -16804
rect 2670 -16888 2715 -16872
rect 2719 -16888 2747 -16708
rect 2850 -16740 2859 -16689
rect 2962 -16714 3006 -16680
rect 3028 -16672 3095 -16666
rect 3172 -16669 3194 -16666
rect 3028 -16706 3085 -16672
rect 3128 -16680 3194 -16669
rect 3195 -16672 6703 -16666
rect 6893 -16671 7025 -16639
rect 7120 -16645 7147 -16637
rect 7169 -16639 7223 -16637
rect 3028 -16714 3048 -16706
rect 3139 -16714 3194 -16680
rect 2753 -16888 2781 -16742
rect 2793 -16778 2804 -16767
rect 2789 -16809 2804 -16778
rect 2789 -16820 2798 -16809
rect 2786 -16862 2804 -16820
rect 2823 -16846 2832 -16812
rect 2835 -16846 2846 -16809
rect 2851 -16846 2896 -16826
rect 2823 -16860 2896 -16846
rect 2789 -16880 2798 -16862
rect 2789 -16888 2817 -16880
rect 2823 -16888 2851 -16860
rect 2950 -16888 3006 -16714
rect 3128 -16715 3194 -16714
rect 3068 -16762 3194 -16715
rect 3115 -16796 3194 -16762
rect 3128 -16832 3194 -16796
rect 3206 -16684 6703 -16672
rect 7034 -16673 7044 -16663
rect 6859 -16681 7049 -16673
rect 3206 -16718 6823 -16684
rect 6835 -16705 7049 -16681
rect 3206 -16737 6703 -16718
rect 3206 -16744 5784 -16737
rect 3206 -16785 5718 -16744
rect 5801 -16752 5872 -16743
rect 5888 -16744 6703 -16737
rect 6835 -16723 6902 -16705
rect 6835 -16727 6897 -16723
rect 7034 -16727 7049 -16705
rect 7075 -16693 7083 -16645
rect 7120 -16671 7128 -16645
rect 7169 -16671 7239 -16639
rect 7247 -16665 7295 -16637
rect 7319 -16637 7456 -16631
rect 7508 -16637 7627 -16616
rect 7790 -16631 7794 -16615
rect 7810 -16624 7904 -16608
rect 7905 -16612 7969 -16608
rect 7319 -16665 7409 -16637
rect 7517 -16640 7605 -16637
rect 7365 -16666 7409 -16665
rect 7128 -16679 7205 -16673
rect 7135 -16681 7205 -16679
rect 7134 -16689 7205 -16681
rect 7075 -16707 7129 -16693
rect 7135 -16705 7205 -16689
rect 7145 -16723 7189 -16705
rect 7365 -16727 7409 -16700
rect 7414 -16727 7422 -16645
rect 7448 -16727 7456 -16645
rect 7484 -16727 7492 -16645
rect 7518 -16727 7526 -16645
rect 7557 -16654 7605 -16640
rect 7775 -16646 7794 -16631
rect 7855 -16640 7870 -16624
rect 7889 -16628 7904 -16624
rect 7530 -16727 7540 -16663
rect 7546 -16665 7605 -16654
rect 7546 -16688 7590 -16665
rect 7728 -16686 7776 -16668
rect 7800 -16686 7848 -16668
rect 7901 -16674 7904 -16628
rect 7955 -16628 7969 -16612
rect 7546 -16727 7590 -16722
rect 7598 -16727 7606 -16688
rect 7728 -16712 7849 -16686
rect 7632 -16727 7640 -16720
rect 5767 -16785 5776 -16775
rect 3206 -16819 5784 -16785
rect 5801 -16809 5810 -16752
rect 5811 -16793 5856 -16759
rect 5888 -16780 6038 -16744
rect 6097 -16752 6194 -16744
rect 6239 -16752 6520 -16744
rect 3200 -16832 5784 -16819
rect 3128 -16853 5784 -16832
rect 6014 -16838 6059 -16804
rect 5792 -16853 5842 -16845
rect 3128 -16861 5792 -16853
rect 3128 -16874 5784 -16861
rect 2635 -16894 3006 -16888
rect 2635 -16903 2819 -16894
rect 2071 -16929 2573 -16921
rect 1752 -16958 1830 -16952
rect 1732 -16964 1849 -16958
rect 1384 -17003 1388 -17000
rect 1305 -17029 1333 -17021
rect 1354 -17029 1526 -17011
rect 1305 -17036 1545 -17029
rect 1331 -17045 1545 -17036
rect 1577 -17045 1653 -17011
rect 1666 -17019 1687 -16977
rect 1732 -16992 1777 -16964
rect 1804 -16992 1849 -16964
rect 1877 -17006 1910 -16952
rect 1911 -16964 2045 -16952
rect 1911 -16972 2003 -16964
rect 1929 -16995 2003 -16972
rect 2112 -16995 2573 -16929
rect 2650 -16906 2817 -16903
rect 2650 -16940 2672 -16906
rect 2719 -16940 2747 -16906
rect 2753 -16940 2817 -16906
rect 2823 -16928 3006 -16894
rect 2823 -16940 2851 -16928
rect 2928 -16940 3006 -16928
rect 3016 -16940 5784 -16874
rect 5792 -16895 5837 -16861
rect 6014 -16906 6059 -16872
rect 6063 -16922 6072 -16788
rect 732 -17076 774 -17052
rect 934 -17076 981 -17052
rect 1331 -17071 1373 -17045
rect 1738 -17046 1742 -17043
rect 1659 -17072 1687 -17064
rect 1708 -17072 1880 -17054
rect 1659 -17079 1899 -17072
rect 1685 -17088 1899 -17079
rect 1931 -17088 1976 -17054
rect 1986 -17069 2007 -17054
rect 2020 -17062 2041 -17020
rect 2086 -17035 2131 -17001
rect 2138 -17003 2220 -16995
rect 2306 -17001 2337 -16995
rect 2158 -17035 2203 -17003
rect 2230 -17035 2275 -17001
rect 2302 -17035 2347 -17001
rect 2362 -17003 2472 -16995
rect 2477 -17003 2573 -16995
rect 2614 -16950 5784 -16940
rect 2614 -16961 5792 -16950
rect 6097 -16956 6106 -16762
rect 6137 -16778 6148 -16767
rect 6133 -16809 6148 -16778
rect 6459 -16796 6504 -16762
rect 2448 -17005 2531 -17003
rect 2477 -17038 2531 -17005
rect 2614 -17038 5784 -16961
rect 5792 -16995 5837 -16961
rect 6037 -16991 6048 -16980
rect 5792 -17011 5842 -17003
rect 5992 -17025 6048 -16991
rect 6133 -16992 6142 -16809
rect 6167 -16995 6176 -16812
rect 2616 -17046 2636 -17038
rect 2640 -17050 2693 -17038
rect 2813 -17046 2846 -17038
rect 2746 -17050 2846 -17046
rect 2400 -17051 2434 -17050
rect 2239 -17067 2311 -17063
rect 2390 -17067 2450 -17063
rect 1979 -17088 2007 -17069
rect 1685 -17114 1727 -17088
rect 2062 -17101 2522 -17097
rect 2013 -17122 2041 -17103
rect 2062 -17111 2234 -17101
rect 2270 -17111 2370 -17101
rect 2381 -17111 2426 -17101
rect 2062 -17131 2427 -17111
rect 2477 -17131 2522 -17101
rect 2534 -17131 2553 -17097
rect 2568 -17164 2587 -17063
rect 2828 -17067 2846 -17050
rect 2947 -17078 2992 -17044
rect 3013 -17050 5784 -17038
rect 3019 -17078 3064 -17050
rect 3028 -17132 3032 -17129
rect 3067 -17140 5784 -17050
rect 6179 -17076 6190 -16809
rect 6516 -16812 6520 -16752
rect 6550 -16819 6554 -16744
rect 6835 -16753 7242 -16727
rect 6809 -16761 7242 -16753
rect 7261 -16761 7657 -16727
rect 7694 -16746 7840 -16720
rect 7894 -16740 7904 -16729
rect 7955 -16740 7966 -16628
rect 7977 -16651 10053 -16608
rect 10073 -16567 10087 -16565
rect 10073 -16578 10092 -16567
rect 10134 -16578 10148 -16567
rect 10218 -16571 10302 -16565
rect 10073 -16628 10087 -16578
rect 10089 -16612 10148 -16578
rect 10234 -16581 10302 -16571
rect 10236 -16621 10302 -16581
rect 10119 -16646 10302 -16621
rect 10313 -16632 10316 -16565
rect 10347 -16637 10350 -16541
rect 7989 -16657 8003 -16651
rect 8167 -16657 8220 -16651
rect 7989 -16668 8000 -16657
rect 8160 -16662 8220 -16657
rect 8160 -16668 8204 -16662
rect 7989 -16702 8037 -16668
rect 8061 -16702 8109 -16668
rect 8133 -16691 8204 -16668
rect 8133 -16702 8181 -16691
rect 7989 -16712 8000 -16702
rect 8212 -16718 8220 -16662
rect 6809 -16819 7205 -16761
rect 7331 -16795 7448 -16786
rect 6195 -16860 6240 -16826
rect 6544 -16830 6565 -16819
rect 6544 -16832 6554 -16830
rect 6195 -16928 6240 -16894
rect 6247 -16995 6256 -16860
rect 6478 -16874 6554 -16832
rect 6607 -16874 7205 -16819
rect 7335 -16819 7345 -16795
rect 7335 -16835 7387 -16819
rect 7343 -16853 7387 -16835
rect 7388 -16853 7398 -16808
rect 7484 -16820 7492 -16761
rect 7518 -16794 7526 -16761
rect 7530 -16794 7540 -16761
rect 7498 -16835 7540 -16794
rect 7598 -16823 7606 -16761
rect 7632 -16808 7640 -16761
rect 7698 -16770 7700 -16761
rect 7749 -16770 7793 -16746
rect 7794 -16770 7804 -16746
rect 7905 -16770 7949 -16740
rect 8246 -16752 8254 -16651
rect 8262 -16672 8296 -16651
rect 8331 -16662 10053 -16651
rect 8331 -16668 10047 -16662
rect 8301 -16694 10053 -16668
rect 10182 -16681 10230 -16668
rect 10179 -16687 10246 -16681
rect 8301 -16702 8349 -16694
rect 8373 -16702 8421 -16694
rect 8445 -16702 8493 -16694
rect 8514 -16734 8558 -16700
rect 8566 -16736 8574 -16694
rect 8422 -16761 8574 -16736
rect 8600 -16770 8608 -16694
rect 8613 -16702 8661 -16694
rect 8685 -16702 10053 -16694
rect 10182 -16689 10230 -16687
rect 10182 -16702 10235 -16689
rect 8685 -16737 10047 -16702
rect 10191 -16714 10235 -16702
rect 10236 -16714 10246 -16687
rect 10254 -16702 10302 -16668
rect 10378 -16673 10388 -16525
rect 10401 -16541 10407 -16491
rect 10435 -16207 10441 -16191
rect 10492 -16207 10502 -16199
rect 10513 -16207 10590 -16178
rect 10649 -16169 11300 -16154
rect 10649 -16188 11215 -16169
rect 11256 -16188 11300 -16169
rect 11322 -16163 11442 -16144
rect 11494 -16163 11557 -16138
rect 11577 -16144 11591 -16122
rect 11639 -16138 11653 -16130
rect 11695 -16138 11709 -16130
rect 11650 -16144 11709 -16138
rect 11755 -16144 11769 -16122
rect 11577 -16163 11625 -16144
rect 11649 -16163 11709 -16144
rect 11322 -16178 11713 -16163
rect 11721 -16178 11769 -16144
rect 11330 -16188 11331 -16178
rect 11359 -16184 11713 -16178
rect 10435 -16241 10485 -16207
rect 10503 -16212 10590 -16207
rect 10687 -16212 10751 -16188
rect 10503 -16241 10557 -16212
rect 10435 -16507 10441 -16241
rect 10739 -16244 10751 -16212
rect 10773 -16244 10785 -16188
rect 10843 -16210 10902 -16188
rect 10965 -16234 10977 -16188
rect 10999 -16212 11063 -16188
rect 10999 -16234 11011 -16212
rect 11053 -16234 11063 -16212
rect 11087 -16234 11097 -16188
rect 11155 -16201 11203 -16188
rect 11330 -16200 11361 -16188
rect 11543 -16191 11557 -16184
rect 11577 -16191 11591 -16184
rect 11387 -16199 11685 -16191
rect 11155 -16210 11215 -16201
rect 11322 -16210 11361 -16200
rect 11383 -16206 11685 -16199
rect 11695 -16206 11709 -16195
rect 11383 -16210 11709 -16206
rect 11200 -16216 11219 -16210
rect 10832 -16250 10846 -16248
rect 10576 -16262 10590 -16251
rect 10492 -16290 10502 -16279
rect 10513 -16290 10590 -16262
rect 10671 -16262 10715 -16250
rect 10743 -16251 10787 -16250
rect 10732 -16262 10787 -16251
rect 10671 -16284 10787 -16262
rect 10815 -16259 10859 -16250
rect 10888 -16259 10902 -16248
rect 11057 -16250 11123 -16239
rect 11144 -16242 11219 -16216
rect 11322 -16231 11709 -16210
rect 11211 -16248 11219 -16242
rect 11144 -16250 11219 -16248
rect 11234 -16250 11244 -16242
rect 11245 -16250 11253 -16234
rect 11288 -16250 11310 -16234
rect 10815 -16284 10902 -16259
rect 10959 -16262 11003 -16250
rect 11031 -16259 11219 -16250
rect 11031 -16262 11147 -16259
rect 10959 -16284 11147 -16262
rect 10503 -16296 10590 -16290
rect 10687 -16296 10746 -16284
rect 10843 -16293 10902 -16284
rect 10999 -16296 11058 -16284
rect 11155 -16293 11219 -16259
rect 10503 -16324 10547 -16296
rect 10576 -16345 10590 -16334
rect 10676 -16345 10690 -16334
rect 10732 -16345 10746 -16334
rect 10832 -16340 10846 -16329
rect 10888 -16340 10902 -16329
rect 11057 -16333 11123 -16322
rect 11211 -16329 11219 -16293
rect 11245 -16284 11310 -16250
rect 10492 -16374 10502 -16363
rect 10513 -16374 10590 -16345
rect 10503 -16379 10590 -16374
rect 10687 -16379 10746 -16345
rect 10843 -16374 10902 -16340
rect 10988 -16345 11002 -16334
rect 11044 -16345 11058 -16334
rect 10999 -16379 11058 -16345
rect 11068 -16367 11123 -16333
rect 11144 -16340 11219 -16329
rect 11234 -16333 11244 -16322
rect 11245 -16333 11253 -16284
rect 11288 -16333 11310 -16284
rect 11155 -16374 11219 -16340
rect 10503 -16408 10547 -16379
rect 10492 -16456 10502 -16446
rect 10525 -16456 10559 -16433
rect 10492 -16457 10559 -16456
rect 10502 -16499 10559 -16457
rect 10855 -16444 10967 -16416
rect 10855 -16458 10863 -16444
rect 10889 -16458 10933 -16450
rect 10959 -16458 10967 -16444
rect 11056 -16458 11134 -16387
rect 10721 -16480 11134 -16458
rect 10502 -16506 10552 -16499
rect 10504 -16514 10552 -16506
rect 10572 -16505 10620 -16480
rect 10640 -16505 10688 -16480
rect 10708 -16505 11134 -16480
rect 11211 -16410 11219 -16374
rect 11245 -16367 11310 -16333
rect 11245 -16376 11253 -16367
rect 10572 -16516 10689 -16505
rect 10708 -16514 11144 -16505
rect 10721 -16516 10832 -16514
rect 10855 -16516 10863 -16514
rect 10572 -16534 10863 -16516
rect 10888 -16516 10988 -16514
rect 11044 -16516 11144 -16514
rect 10888 -16531 11144 -16516
rect 11211 -16520 11220 -16410
rect 11234 -16417 11244 -16406
rect 11245 -16417 11254 -16376
rect 11288 -16417 11310 -16367
rect 11245 -16451 11310 -16417
rect 11322 -16244 11397 -16231
rect 11494 -16240 11557 -16231
rect 11322 -16316 11361 -16244
rect 11484 -16282 11539 -16259
rect 11428 -16285 11539 -16282
rect 11428 -16293 11494 -16285
rect 11383 -16316 11397 -16305
rect 11322 -16350 11397 -16316
rect 11411 -16309 11527 -16293
rect 11543 -16309 11557 -16240
rect 11411 -16327 11557 -16309
rect 11322 -16384 11361 -16350
rect 11494 -16354 11557 -16327
rect 11383 -16384 11397 -16373
rect 11428 -16375 11494 -16365
rect 11428 -16376 11542 -16375
rect 11322 -16418 11397 -16384
rect 11439 -16377 11542 -16376
rect 11543 -16377 11557 -16354
rect 11439 -16410 11557 -16377
rect 11322 -16430 11361 -16418
rect 11494 -16422 11557 -16410
rect 11322 -16438 11344 -16430
rect 11234 -16500 11244 -16489
rect 11245 -16500 11254 -16451
rect 11288 -16472 11310 -16451
rect 11427 -16449 11484 -16430
rect 11427 -16494 11494 -16449
rect 11543 -16463 11557 -16422
rect 11577 -16282 11591 -16231
rect 11650 -16240 11709 -16231
rect 11755 -16240 11769 -16178
rect 11789 -16130 11803 -16122
rect 11855 -16130 11869 -16122
rect 11789 -16138 11809 -16130
rect 11851 -16138 11869 -16130
rect 11789 -16195 11803 -16138
rect 11806 -16172 11869 -16138
rect 11855 -16195 11869 -16172
rect 11789 -16206 11809 -16195
rect 11851 -16206 11869 -16195
rect 11789 -16240 11803 -16206
rect 11806 -16240 11869 -16206
rect 11889 -16144 11903 -16122
rect 11951 -16138 11965 -16130
rect 12007 -16138 12021 -16130
rect 11962 -16144 12021 -16138
rect 12067 -16144 12081 -16122
rect 11889 -16178 11937 -16144
rect 11961 -16172 12021 -16144
rect 11961 -16178 12009 -16172
rect 12033 -16178 12081 -16144
rect 11889 -16240 11903 -16178
rect 11951 -16206 11965 -16195
rect 12007 -16206 12021 -16195
rect 11962 -16240 12021 -16206
rect 11741 -16274 12039 -16240
rect 12067 -16249 12081 -16178
rect 11577 -16293 11650 -16282
rect 11577 -16365 11591 -16293
rect 11595 -16309 11650 -16293
rect 11595 -16320 11653 -16309
rect 11695 -16320 11709 -16309
rect 11755 -16320 11769 -16274
rect 11789 -16309 11803 -16274
rect 11838 -16309 11851 -16302
rect 11855 -16309 11869 -16274
rect 11789 -16320 11809 -16309
rect 11838 -16320 11869 -16309
rect 11889 -16286 11903 -16274
rect 11595 -16327 11709 -16320
rect 11806 -16325 11887 -16320
rect 11650 -16354 11709 -16327
rect 11782 -16336 11887 -16325
rect 11577 -16376 11650 -16365
rect 11765 -16370 11887 -16336
rect 11838 -16375 11851 -16370
rect 11577 -16438 11591 -16376
rect 11595 -16377 11650 -16376
rect 11806 -16377 11854 -16375
rect 11855 -16377 11887 -16370
rect 11595 -16388 11653 -16377
rect 11695 -16388 11709 -16377
rect 11795 -16388 11887 -16377
rect 11595 -16410 11709 -16388
rect 11803 -16408 11887 -16388
rect 11650 -16422 11709 -16410
rect 11782 -16419 11887 -16408
rect 11793 -16422 11887 -16419
rect 11793 -16430 11837 -16422
rect 11579 -16449 11591 -16438
rect 11594 -16449 11651 -16430
rect 11579 -16460 11651 -16449
rect 11579 -16463 11591 -16460
rect 11594 -16463 11651 -16460
rect 11245 -16514 11289 -16500
rect 11427 -16514 11484 -16494
rect 11211 -16531 11219 -16520
rect 10888 -16534 11219 -16531
rect 11245 -16532 11484 -16514
rect 11543 -16510 11651 -16463
rect 11781 -16453 11837 -16430
rect 11838 -16453 11848 -16422
rect 11781 -16472 11809 -16453
rect 11855 -16463 11887 -16422
rect 11889 -16438 11921 -16286
rect 11951 -16320 11965 -16309
rect 12007 -16320 12021 -16309
rect 11962 -16325 12021 -16320
rect 11938 -16336 12021 -16325
rect 11949 -16354 12021 -16336
rect 12061 -16351 12081 -16249
rect 12101 -16130 12115 -16122
rect 12167 -16130 12181 -16122
rect 12101 -16138 12121 -16130
rect 12163 -16138 12181 -16130
rect 12101 -16195 12115 -16138
rect 12118 -16172 12181 -16138
rect 12167 -16195 12181 -16172
rect 12101 -16206 12121 -16195
rect 12163 -16206 12181 -16195
rect 12101 -16283 12115 -16206
rect 12118 -16240 12181 -16206
rect 12167 -16283 12181 -16240
rect 12201 -16144 12215 -16122
rect 12263 -16138 12277 -16130
rect 12319 -16138 12333 -16130
rect 12274 -16144 12333 -16138
rect 12379 -16144 12393 -16122
rect 12201 -16178 12249 -16144
rect 12273 -16172 12333 -16144
rect 12273 -16178 12321 -16172
rect 12345 -16178 12393 -16144
rect 12201 -16283 12215 -16178
rect 12263 -16206 12277 -16195
rect 12319 -16206 12333 -16195
rect 12274 -16240 12333 -16206
rect 12379 -16283 12393 -16178
rect 12413 -16130 12427 -16122
rect 12479 -16130 12493 -16122
rect 12413 -16138 12433 -16130
rect 12475 -16138 12493 -16130
rect 12413 -16195 12427 -16138
rect 12430 -16172 12493 -16138
rect 12479 -16195 12493 -16172
rect 12413 -16206 12433 -16195
rect 12475 -16206 12493 -16195
rect 12413 -16283 12427 -16206
rect 12430 -16240 12493 -16206
rect 12479 -16283 12493 -16240
rect 12513 -16144 12527 -16122
rect 12575 -16138 12589 -16130
rect 12631 -16138 12645 -16130
rect 12586 -16144 12645 -16138
rect 12691 -16144 12705 -16122
rect 12513 -16178 12561 -16144
rect 12585 -16172 12645 -16144
rect 12585 -16178 12633 -16172
rect 12657 -16178 12705 -16144
rect 12513 -16283 12527 -16178
rect 12575 -16206 12589 -16195
rect 12631 -16206 12645 -16195
rect 12586 -16240 12645 -16206
rect 12095 -16309 12585 -16283
rect 12095 -16317 12589 -16309
rect 11949 -16370 11993 -16354
rect 11951 -16388 11965 -16377
rect 12007 -16388 12021 -16377
rect 11959 -16408 12021 -16388
rect 11938 -16419 12021 -16408
rect 11949 -16422 12021 -16419
rect 11949 -16430 11993 -16422
rect 11948 -16453 12005 -16430
rect 12067 -16438 12081 -16351
rect 12101 -16320 12121 -16317
rect 12163 -16320 12181 -16317
rect 12101 -16377 12115 -16320
rect 12118 -16354 12181 -16320
rect 12167 -16363 12181 -16354
rect 12201 -16363 12215 -16317
rect 12263 -16320 12277 -16317
rect 12319 -16320 12333 -16317
rect 12274 -16345 12333 -16320
rect 12263 -16354 12333 -16345
rect 12118 -16377 12166 -16375
rect 12172 -16377 12238 -16368
rect 12263 -16371 12319 -16354
rect 12379 -16363 12393 -16317
rect 12413 -16320 12433 -16317
rect 12475 -16320 12493 -16317
rect 12413 -16329 12427 -16320
rect 12430 -16329 12493 -16320
rect 12413 -16354 12493 -16329
rect 12379 -16368 12399 -16363
rect 12328 -16377 12399 -16368
rect 12101 -16379 12238 -16377
rect 12101 -16388 12177 -16379
rect 11948 -16463 11965 -16453
rect 11992 -16457 12005 -16453
rect 11990 -16463 12005 -16457
rect 11855 -16472 11965 -16463
rect 11971 -16472 12005 -16463
rect 11781 -16492 11838 -16472
rect 11245 -16534 11494 -16532
rect 10572 -16547 10689 -16534
rect 10690 -16547 10832 -16534
rect 10888 -16545 10988 -16534
rect 10838 -16547 10988 -16545
rect 11044 -16547 11144 -16534
rect 10493 -16565 11241 -16547
rect 10075 -16736 10341 -16714
rect 8776 -16746 8839 -16737
rect 8891 -16743 8974 -16737
rect 8904 -16770 8974 -16743
rect 8995 -16770 8998 -16737
rect 9026 -16770 9036 -16737
rect 9146 -16770 9200 -16737
rect 9233 -16753 10047 -16737
rect 10378 -16741 10393 -16673
rect 10419 -16707 10427 -16639
rect 10447 -16673 10472 -16603
rect 10481 -16665 10506 -16569
rect 10576 -16573 11241 -16565
rect 10519 -16587 11241 -16573
rect 10508 -16608 11241 -16587
rect 11245 -16554 11254 -16534
rect 10508 -16621 10590 -16608
rect 10519 -16655 10572 -16621
rect 10671 -16632 10791 -16608
rect 10792 -16620 10800 -16608
rect 10832 -16620 10842 -16608
rect 10983 -16615 11058 -16608
rect 10891 -16620 10972 -16616
rect 10519 -16665 10534 -16655
rect 10481 -16670 10534 -16665
rect 10689 -16666 10791 -16632
rect 10689 -16670 10732 -16666
rect 10735 -16670 10791 -16666
rect 10481 -16673 10519 -16670
rect 10488 -16681 10519 -16673
rect 10576 -16681 10590 -16670
rect 10676 -16681 10791 -16670
rect 10478 -16689 10488 -16681
rect 10499 -16689 10590 -16681
rect 10489 -16715 10590 -16689
rect 10687 -16715 10791 -16681
rect 10489 -16717 10533 -16715
rect 10689 -16717 10791 -16715
rect 10832 -16638 10972 -16620
rect 10832 -16640 10842 -16638
rect 10874 -16640 10888 -16638
rect 10891 -16640 10972 -16638
rect 10832 -16651 10846 -16640
rect 10874 -16651 10972 -16640
rect 10832 -16717 10842 -16651
rect 10843 -16685 10972 -16651
rect 10852 -16717 10972 -16685
rect 10103 -16753 10313 -16742
rect 10378 -16753 10388 -16741
rect 10487 -16751 10535 -16717
rect 10559 -16751 10607 -16717
rect 10689 -16723 10811 -16717
rect 10832 -16722 10972 -16717
rect 10983 -16670 11044 -16615
rect 10983 -16715 11058 -16670
rect 11104 -16674 11114 -16608
rect 11138 -16640 11219 -16608
rect 11139 -16668 11219 -16640
rect 10983 -16720 11044 -16715
rect 11105 -16720 11114 -16674
rect 10832 -16723 10888 -16722
rect 10709 -16734 10753 -16723
rect 10763 -16751 10811 -16723
rect 10835 -16749 10888 -16723
rect 10890 -16723 10972 -16722
rect 10976 -16723 11044 -16720
rect 11138 -16723 11219 -16668
rect 10835 -16751 10884 -16749
rect 7709 -16804 7980 -16770
rect 8028 -16804 8076 -16770
rect 8124 -16771 8268 -16770
rect 8087 -16804 8311 -16771
rect 8316 -16804 8364 -16770
rect 8367 -16804 8748 -16770
rect 8796 -16779 8844 -16770
rect 8884 -16779 9228 -16770
rect 9233 -16779 10549 -16753
rect 10757 -16757 10792 -16752
rect 8753 -16780 10549 -16779
rect 8753 -16804 9267 -16780
rect 9276 -16804 9708 -16780
rect 9756 -16804 10549 -16780
rect 10723 -16791 10792 -16786
rect 7630 -16819 7640 -16808
rect 8099 -16813 8143 -16804
rect 8144 -16813 8154 -16804
rect 8255 -16813 8299 -16804
rect 6478 -16877 7205 -16874
rect 6281 -16980 6290 -16892
rect 6393 -16900 6443 -16892
rect 6443 -16908 6454 -16900
rect 6398 -16942 6454 -16908
rect 6279 -16991 6290 -16980
rect 6281 -17025 6335 -16991
rect 6443 -17008 6454 -16997
rect 6398 -17042 6454 -17008
rect 6478 -17044 6633 -16877
rect 6809 -16899 7205 -16877
rect 6733 -16925 7205 -16899
rect 7530 -16904 7540 -16835
rect 7632 -16853 7640 -16819
rect 7641 -16853 7685 -16819
rect 7749 -16870 7793 -16836
rect 7794 -16870 7804 -16825
rect 7894 -16832 7904 -16821
rect 7905 -16866 7949 -16832
rect 8415 -16838 8543 -16806
rect 8598 -16822 8665 -16814
rect 8441 -16856 8508 -16838
rect 7642 -16906 7686 -16872
rect 7714 -16906 7758 -16872
rect 7786 -16906 7830 -16872
rect 8099 -16913 8143 -16879
rect 8144 -16913 8154 -16868
rect 8244 -16879 8254 -16868
rect 8441 -16878 8498 -16856
rect 8608 -16878 8665 -16822
rect 9026 -16845 9036 -16804
rect 9026 -16853 9041 -16845
rect 8827 -16878 8894 -16853
rect 8994 -16878 9041 -16853
rect 8255 -16913 8299 -16879
rect 8839 -16895 8883 -16878
rect 8884 -16895 8894 -16878
rect 6733 -16959 7218 -16925
rect 8067 -16949 8111 -16915
rect 8139 -16949 8183 -16915
rect 8453 -16956 8497 -16922
rect 8498 -16956 8508 -16911
rect 8598 -16922 8608 -16911
rect 9026 -16913 9041 -16878
rect 9067 -16879 9075 -16811
rect 9112 -16843 9120 -16804
rect 9146 -16809 9154 -16804
rect 9359 -16838 9403 -16804
rect 9126 -16861 9136 -16853
rect 9137 -16895 9181 -16861
rect 9359 -16906 9403 -16872
rect 8609 -16956 8653 -16922
rect 6733 -16985 7205 -16959
rect 6736 -16993 6947 -16985
rect 6752 -17003 6931 -16993
rect 6291 -17078 6336 -17044
rect 6363 -17050 6408 -17044
rect 6435 -17050 6633 -17044
rect 6363 -17058 6633 -17050
rect 6363 -17078 6408 -17058
rect 6435 -17078 6633 -17058
rect 5821 -17131 5866 -17097
rect 6478 -17114 6633 -17078
rect 6478 -17140 6663 -17114
rect 2610 -17150 2726 -17140
rect 2737 -17150 2928 -17140
rect 2929 -17150 2974 -17140
rect 2610 -17158 2975 -17150
rect 3025 -17157 5784 -17140
rect 3025 -17158 5718 -17157
rect 2610 -17174 5718 -17158
rect 5985 -17174 6030 -17140
rect 6081 -17174 6126 -17140
rect 6177 -17174 6222 -17140
rect 6273 -17174 6318 -17140
rect 6369 -17174 6414 -17140
rect 6465 -17174 6663 -17140
rect 2726 -17248 2768 -17224
rect 2928 -17248 2975 -17224
rect 3067 -17458 5718 -17174
rect 6478 -17200 6663 -17174
rect 6678 -17174 6789 -17050
rect 6937 -17062 6947 -17051
rect 2687 -17970 3066 -17936
rect 3145 -17971 3191 -17458
rect 3200 -17604 5718 -17458
rect 3200 -17858 5784 -17604
rect 3200 -17971 5718 -17858
rect 3135 -18032 5718 -17971
rect 2591 -18194 2636 -18032
rect 2787 -18108 2966 -18074
rect 3117 -18128 5718 -18032
rect 2725 -18182 2770 -18151
rect 2771 -18182 2781 -18156
rect 2952 -18182 3040 -18155
rect 2713 -18194 3096 -18182
rect 2591 -18228 3096 -18194
rect 2557 -18240 2558 -18228
rect 2591 -18240 2636 -18228
rect 2713 -18229 3096 -18228
rect 3105 -18229 5718 -18128
rect 2713 -18240 5718 -18229
rect 2525 -18506 2570 -18240
rect 2579 -18506 2636 -18240
rect 2725 -18301 2770 -18240
rect 2713 -18316 2770 -18301
rect 2771 -18316 2781 -18240
rect 2952 -18265 5718 -18240
rect 2713 -18332 2772 -18316
rect 2888 -18332 2935 -18285
rect 2713 -18366 2935 -18332
rect 2646 -18506 2648 -18413
rect 2658 -18506 2670 -18409
rect 2691 -18413 2692 -18409
rect 2713 -18413 2771 -18366
rect 2983 -18385 3028 -18265
rect 2949 -18413 2950 -18409
rect 2691 -18415 2698 -18413
rect 2719 -18415 2770 -18413
rect 2949 -18414 2956 -18413
rect 2691 -18425 2692 -18415
rect 2687 -18506 2692 -18425
rect 2725 -18506 2770 -18415
rect 2905 -18425 2956 -18414
rect 2916 -18506 2956 -18425
rect 2977 -18506 3028 -18385
rect 3038 -18506 3040 -18265
rect 3050 -18506 5718 -18265
rect 2525 -18764 5718 -18506
rect 2477 -19282 5718 -18764
rect 5857 -17936 6038 -17858
rect 6556 -17870 6601 -17200
rect 6678 -17228 6735 -17174
rect 5857 -17970 6410 -17936
rect 5857 -18506 6038 -17970
rect 6490 -17971 6518 -17924
rect 6544 -17971 6601 -17870
rect 6690 -17971 6735 -17228
rect 6736 -17971 6746 -17174
rect 6948 -17971 6993 -17062
rect 7082 -17971 7127 -16985
rect 7336 -17002 7380 -16968
rect 7432 -17002 7476 -16968
rect 7528 -17002 7572 -16968
rect 7624 -17002 7668 -16968
rect 7720 -17002 7764 -16968
rect 7816 -17002 7860 -16968
rect 7912 -17002 7956 -16968
rect 8421 -16992 8465 -16958
rect 8493 -16992 8537 -16958
rect 8839 -16995 8883 -16961
rect 8884 -16995 8894 -16950
rect 9026 -17001 9036 -16913
rect 9408 -16922 9416 -16804
rect 9126 -16961 9136 -16950
rect 9442 -16956 9450 -16804
rect 9478 -16809 9492 -16804
rect 9137 -16995 9181 -16961
rect 8074 -17045 8118 -17011
rect 8170 -17045 8214 -17011
rect 8266 -17045 8310 -17011
rect 8775 -17035 8819 -17001
rect 8847 -17035 8891 -17001
rect 8919 -17035 8963 -17001
rect 8991 -17029 9036 -17001
rect 9337 -17025 9381 -16991
rect 9382 -17025 9392 -16980
rect 9478 -16992 9486 -16809
rect 9524 -16812 9534 -16809
rect 9512 -16838 9600 -16812
rect 9823 -16830 10549 -16804
rect 10828 -16813 10836 -16757
rect 10862 -16813 10870 -16757
rect 10874 -16813 10884 -16751
rect 10890 -16751 10961 -16723
rect 10890 -16756 10934 -16751
rect 10942 -16757 10961 -16751
rect 10942 -16813 10950 -16757
rect 10976 -16785 10995 -16723
rect 11088 -16728 11138 -16723
rect 11145 -16728 11193 -16723
rect 11081 -16749 11193 -16728
rect 11081 -16764 11137 -16749
rect 11093 -16770 11137 -16764
rect 11138 -16751 11193 -16749
rect 11138 -16770 11148 -16751
rect 11211 -16757 11219 -16723
rect 11245 -16729 11253 -16554
rect 11261 -16556 11494 -16534
rect 11543 -16556 11557 -16510
rect 11577 -16556 11591 -16510
rect 11593 -16514 11651 -16510
rect 11706 -16514 11754 -16510
rect 11781 -16514 11848 -16492
rect 11593 -16537 11848 -16514
rect 11855 -16510 12005 -16472
rect 11593 -16544 11838 -16537
rect 11594 -16556 11838 -16544
rect 11855 -16556 11887 -16510
rect 11889 -16514 12005 -16510
rect 12018 -16514 12066 -16510
rect 12067 -16514 12081 -16494
rect 12101 -16514 12115 -16388
rect 12118 -16422 12177 -16388
rect 12183 -16413 12238 -16379
rect 12263 -16379 12399 -16377
rect 12263 -16413 12333 -16379
rect 12339 -16413 12399 -16379
rect 12274 -16422 12333 -16413
rect 12379 -16430 12399 -16413
rect 12171 -16451 12228 -16430
rect 12171 -16463 12238 -16451
rect 12305 -16463 12313 -16438
rect 12338 -16451 12399 -16430
rect 12328 -16462 12399 -16451
rect 12338 -16463 12399 -16462
rect 12413 -16371 12475 -16354
rect 12479 -16363 12493 -16354
rect 12513 -16363 12527 -16317
rect 12575 -16320 12589 -16317
rect 12631 -16320 12645 -16309
rect 12586 -16326 12645 -16320
rect 12691 -16326 12705 -16178
rect 12725 -16130 12739 -16122
rect 12791 -16130 12805 -16122
rect 12725 -16138 12745 -16130
rect 12787 -16138 12805 -16130
rect 12725 -16195 12739 -16138
rect 12742 -16172 12805 -16138
rect 12791 -16195 12805 -16172
rect 12725 -16206 12745 -16195
rect 12787 -16206 12805 -16195
rect 12725 -16309 12739 -16206
rect 12742 -16240 12805 -16206
rect 12791 -16309 12805 -16240
rect 12725 -16320 12745 -16309
rect 12787 -16320 12805 -16309
rect 12725 -16326 12739 -16320
rect 12742 -16326 12805 -16320
rect 12825 -16144 12839 -16122
rect 12887 -16138 12901 -16130
rect 12943 -16138 12957 -16130
rect 12898 -16144 12957 -16138
rect 13003 -16144 13017 -16122
rect 12825 -16178 12873 -16144
rect 12897 -16172 12957 -16144
rect 12897 -16178 12945 -16172
rect 12969 -16178 13017 -16144
rect 12825 -16326 12839 -16178
rect 12887 -16206 12901 -16195
rect 12943 -16206 12957 -16195
rect 12898 -16240 12957 -16206
rect 12887 -16320 12901 -16309
rect 12943 -16320 12957 -16309
rect 12898 -16326 12957 -16320
rect 13003 -16326 13017 -16178
rect 13037 -16130 13051 -16122
rect 13103 -16130 13117 -16122
rect 13037 -16138 13057 -16130
rect 13099 -16138 13117 -16130
rect 13037 -16195 13051 -16138
rect 13054 -16172 13117 -16138
rect 13103 -16195 13117 -16172
rect 13037 -16206 13057 -16195
rect 13099 -16206 13117 -16195
rect 13037 -16309 13051 -16206
rect 13054 -16240 13117 -16206
rect 13103 -16309 13117 -16240
rect 13037 -16320 13057 -16309
rect 13099 -16320 13117 -16309
rect 13037 -16326 13051 -16320
rect 13054 -16326 13117 -16320
rect 13137 -16144 13151 -16122
rect 13199 -16138 13213 -16130
rect 13255 -16138 13269 -16130
rect 13210 -16144 13269 -16138
rect 13315 -16144 13329 -16122
rect 13137 -16178 13185 -16144
rect 13209 -16172 13269 -16144
rect 13209 -16178 13257 -16172
rect 13281 -16178 13329 -16144
rect 13137 -16326 13151 -16178
rect 13199 -16206 13213 -16195
rect 13255 -16206 13269 -16195
rect 13210 -16240 13269 -16206
rect 13199 -16320 13213 -16309
rect 13255 -16320 13269 -16309
rect 13210 -16326 13269 -16320
rect 13315 -16326 13329 -16178
rect 12586 -16354 13329 -16326
rect 12643 -16366 13329 -16354
rect 12413 -16375 12433 -16371
rect 12413 -16377 12478 -16375
rect 12484 -16377 12550 -16368
rect 12691 -16375 12705 -16366
rect 12725 -16369 12739 -16366
rect 12791 -16369 12805 -16366
rect 12725 -16375 12805 -16369
rect 12825 -16375 12839 -16366
rect 13003 -16375 13017 -16366
rect 13037 -16369 13051 -16366
rect 13103 -16369 13117 -16366
rect 13037 -16375 13117 -16369
rect 13137 -16375 13151 -16366
rect 13315 -16375 13329 -16366
rect 13349 -16130 13363 -16122
rect 13414 -16130 13429 -16122
rect 13349 -16138 13369 -16130
rect 13411 -16138 13429 -16130
rect 13349 -16172 13363 -16138
rect 13366 -16172 13429 -16138
rect 13448 -16130 13937 -16111
rect 14051 -16119 14164 -16100
rect 14178 -16119 14226 -16085
rect 14274 -16119 14322 -16085
rect 14370 -16119 14418 -16085
rect 14466 -16100 14514 -16085
rect 14434 -16119 14514 -16100
rect 14562 -16100 14610 -16085
rect 14562 -16119 14632 -16100
rect 14658 -16119 14706 -16085
rect 14754 -16119 14802 -16085
rect 14831 -16119 14833 -16085
rect 14051 -16125 14703 -16120
rect 16823 -16128 16866 -16111
rect 16919 -16128 16962 -16111
rect 17015 -16128 17058 -16111
rect 17111 -16128 17154 -16111
rect 17207 -16128 17250 -16111
rect 13448 -16144 13906 -16130
rect 14885 -16143 14887 -16128
rect 14916 -16143 14964 -16128
rect 13448 -16145 13916 -16144
rect 13349 -16184 13448 -16172
rect 13449 -16178 13497 -16145
rect 13521 -16172 13581 -16145
rect 13521 -16178 13569 -16172
rect 13593 -16178 13641 -16145
rect 13349 -16195 13363 -16184
rect 13415 -16195 13429 -16184
rect 13349 -16206 13369 -16195
rect 13411 -16200 13429 -16195
rect 13382 -16206 13448 -16200
rect 13349 -16309 13363 -16206
rect 13366 -16212 13448 -16206
rect 13366 -16240 13429 -16212
rect 13415 -16309 13429 -16240
rect 13349 -16320 13369 -16309
rect 13411 -16320 13429 -16309
rect 13349 -16375 13363 -16320
rect 13366 -16354 13429 -16320
rect 12615 -16377 13363 -16375
rect 13366 -16377 13414 -16375
rect 13415 -16377 13429 -16354
rect 12413 -16379 12550 -16377
rect 12413 -16422 12489 -16379
rect 12495 -16413 12550 -16379
rect 12575 -16388 12589 -16377
rect 12615 -16388 13429 -16377
rect 12586 -16394 13363 -16388
rect 12586 -16422 12645 -16394
rect 12691 -16416 12705 -16394
rect 12725 -16416 12739 -16394
rect 12742 -16416 12805 -16394
rect 12825 -16416 12839 -16394
rect 12742 -16422 12801 -16416
rect 12898 -16422 12957 -16394
rect 13003 -16406 13017 -16394
rect 13037 -16406 13051 -16394
rect 13054 -16406 13117 -16394
rect 13137 -16406 13151 -16394
rect 13054 -16411 13113 -16406
rect 13199 -16411 13273 -16394
rect 13054 -16422 13117 -16411
rect 13199 -16414 13294 -16411
rect 13210 -16422 13294 -16414
rect 12413 -16463 12433 -16422
rect 12494 -16451 12551 -16430
rect 12484 -16462 12551 -16451
rect 12665 -16456 12709 -16422
rect 12737 -16456 12781 -16422
rect 12809 -16456 12853 -16422
rect 12953 -16456 12997 -16422
rect 13025 -16456 13141 -16422
rect 13169 -16456 13213 -16422
rect 12494 -16463 12551 -16462
rect 12171 -16510 12433 -16463
rect 12482 -16510 12551 -16463
rect 13050 -16472 13057 -16456
rect 13099 -16463 13128 -16456
rect 13205 -16463 13213 -16456
rect 13239 -16430 13294 -16422
rect 13239 -16456 13295 -16430
rect 13315 -16438 13329 -16394
rect 13099 -16472 13238 -16463
rect 13239 -16472 13247 -16456
rect 13255 -16472 13295 -16456
rect 13050 -16510 13295 -16472
rect 12171 -16514 12312 -16510
rect 11889 -16523 12312 -16514
rect 12330 -16523 12433 -16510
rect 11889 -16544 12433 -16523
rect 12494 -16514 12577 -16510
rect 12642 -16514 12690 -16510
rect 12841 -16514 12889 -16510
rect 12954 -16514 13002 -16510
rect 13050 -16514 13128 -16510
rect 12494 -16535 13128 -16514
rect 11889 -16556 11921 -16544
rect 11926 -16556 12286 -16544
rect 12310 -16556 12399 -16544
rect 12413 -16556 12433 -16544
rect 12484 -16546 13128 -16535
rect 13153 -16514 13314 -16510
rect 13315 -16514 13329 -16494
rect 13349 -16514 13363 -16394
rect 13366 -16422 13429 -16388
rect 13449 -16409 13463 -16178
rect 13627 -16191 13641 -16178
rect 13661 -16173 13675 -16145
rect 13678 -16172 13741 -16145
rect 13661 -16191 13690 -16173
rect 13511 -16206 13525 -16195
rect 13567 -16196 13581 -16195
rect 13567 -16206 13590 -16196
rect 13667 -16206 13690 -16191
rect 13727 -16191 13741 -16172
rect 13761 -16178 13818 -16145
rect 13834 -16173 13890 -16145
rect 14147 -16148 14164 -16147
rect 14439 -16148 14452 -16147
rect 14023 -16153 14675 -16148
rect 14147 -16154 14164 -16153
rect 14439 -16154 14452 -16153
rect 13997 -16165 14709 -16154
rect 14885 -16162 14971 -16143
rect 15012 -16162 15060 -16128
rect 15108 -16162 15156 -16128
rect 15204 -16162 15252 -16128
rect 15300 -16162 15348 -16128
rect 15396 -16162 15444 -16128
rect 15492 -16162 15540 -16128
rect 15588 -16162 15636 -16128
rect 15684 -16162 15732 -16128
rect 15780 -16162 15828 -16128
rect 15876 -16162 15924 -16128
rect 15972 -16162 16020 -16128
rect 16068 -16162 16116 -16128
rect 16164 -16162 16212 -16128
rect 16260 -16162 16308 -16128
rect 16356 -16162 16404 -16128
rect 16452 -16162 16500 -16128
rect 16548 -16162 16596 -16128
rect 16644 -16162 16692 -16128
rect 16740 -16151 16788 -16128
rect 16823 -16145 16884 -16128
rect 16919 -16145 16980 -16128
rect 17015 -16145 17076 -16128
rect 17111 -16145 17172 -16128
rect 17207 -16145 17268 -16128
rect 16836 -16151 16884 -16145
rect 16925 -16151 17076 -16145
rect 17081 -16151 17190 -16145
rect 17220 -16151 17268 -16145
rect 16740 -16162 17309 -16151
rect 17316 -16162 17364 -16128
rect 17378 -16154 17460 -16128
rect 17474 -16154 17556 -16128
rect 20167 -16145 20210 -16111
rect 20263 -16145 20306 -16111
rect 20359 -16145 20402 -16111
rect 20455 -16145 20498 -16111
rect 20551 -16145 20594 -16111
rect 23511 -16145 23554 -16111
rect 23607 -16145 23650 -16111
rect 23703 -16145 23746 -16111
rect 23799 -16145 23842 -16111
rect 23895 -16145 23938 -16111
rect 26856 -16145 26898 -16111
rect 26952 -16145 26994 -16111
rect 27048 -16145 27090 -16111
rect 27144 -16145 27186 -16111
rect 27240 -16145 27282 -16111
rect 30200 -16145 30242 -16111
rect 30296 -16145 30338 -16111
rect 30392 -16145 30434 -16111
rect 30488 -16145 30530 -16111
rect 30584 -16145 30626 -16111
rect 33544 -16145 33586 -16111
rect 33640 -16145 33682 -16111
rect 33736 -16145 33778 -16111
rect 33832 -16145 33874 -16111
rect 33928 -16145 33970 -16111
rect 36888 -16145 36930 -16111
rect 36984 -16145 37026 -16111
rect 37080 -16145 37122 -16111
rect 37176 -16145 37218 -16111
rect 37272 -16145 37314 -16111
rect 17369 -16162 17460 -16154
rect 17465 -16162 17556 -16154
rect 13997 -16173 14675 -16165
rect 13823 -16178 13890 -16173
rect 13727 -16195 13751 -16191
rect 13723 -16206 13751 -16195
rect 13472 -16241 13515 -16207
rect 13522 -16240 13590 -16206
rect 13536 -16241 13590 -16240
rect 13616 -16241 13659 -16207
rect 13678 -16240 13751 -16206
rect 13692 -16241 13751 -16240
rect 13567 -16290 13590 -16279
rect 13681 -16290 13690 -16279
rect 13723 -16290 13751 -16241
rect 13511 -16320 13525 -16309
rect 13536 -16320 13590 -16290
rect 13667 -16320 13690 -16309
rect 13692 -16320 13751 -16290
rect 13522 -16324 13590 -16320
rect 13522 -16354 13581 -16324
rect 13567 -16374 13590 -16363
rect 13511 -16388 13525 -16377
rect 13536 -16388 13590 -16374
rect 13638 -16375 13657 -16342
rect 13678 -16354 13751 -16320
rect 13681 -16369 13690 -16363
rect 13666 -16374 13690 -16369
rect 13723 -16374 13751 -16354
rect 13666 -16375 13685 -16374
rect 13692 -16375 13751 -16374
rect 13678 -16377 13751 -16375
rect 13667 -16388 13751 -16377
rect 13415 -16514 13429 -16422
rect 13448 -16438 13463 -16409
rect 13522 -16408 13590 -16388
rect 13522 -16422 13581 -16408
rect 13678 -16409 13751 -16388
rect 13448 -16443 13454 -16438
rect 13524 -16456 13550 -16430
rect 13567 -16446 13581 -16430
rect 13638 -16443 13657 -16409
rect 13666 -16415 13751 -16409
rect 13678 -16422 13751 -16415
rect 13524 -16463 13525 -16456
rect 13567 -16457 13590 -16446
rect 13681 -16457 13690 -16446
rect 13723 -16457 13751 -16422
rect 13761 -16438 13785 -16178
rect 13823 -16207 13846 -16178
rect 14025 -16188 14068 -16173
rect 14089 -16181 14675 -16173
rect 14732 -16181 14746 -16173
rect 14756 -16181 14791 -16163
rect 14885 -16168 15057 -16163
rect 16764 -16168 17309 -16162
rect 17338 -16168 17532 -16162
rect 17561 -16168 17604 -16154
rect 14075 -16188 14675 -16181
rect 14681 -16188 14729 -16181
rect 13786 -16210 13846 -16207
rect 13848 -16210 13901 -16207
rect 13786 -16241 13829 -16210
rect 13834 -16241 13901 -16210
rect 14075 -16215 14195 -16188
rect 14275 -16215 14339 -16188
rect 14327 -16234 14339 -16215
rect 14361 -16215 14415 -16188
rect 14431 -16215 14490 -16188
rect 14511 -16215 14565 -16188
rect 14361 -16234 14373 -16215
rect 13834 -16244 13882 -16241
rect 14402 -16250 14434 -16239
rect 14553 -16250 14565 -16215
rect 14587 -16215 14651 -16188
rect 14587 -16216 14599 -16215
rect 14576 -16242 14599 -16216
rect 14641 -16234 14651 -16215
rect 14675 -16215 14729 -16188
rect 14743 -16197 14801 -16181
rect 14857 -16196 15029 -16191
rect 16792 -16196 17281 -16179
rect 17338 -16194 17615 -16168
rect 17657 -16188 17700 -16154
rect 17753 -16188 17796 -16154
rect 17849 -16188 17892 -16154
rect 17945 -16188 17988 -16154
rect 20713 -16188 20756 -16154
rect 20809 -16188 20852 -16154
rect 20905 -16188 20948 -16154
rect 21001 -16188 21044 -16154
rect 21097 -16188 21140 -16154
rect 21193 -16188 21236 -16154
rect 21289 -16188 21332 -16154
rect 24057 -16188 24100 -16154
rect 24153 -16188 24196 -16154
rect 24249 -16188 24292 -16154
rect 24345 -16188 24388 -16154
rect 24441 -16188 24484 -16154
rect 24537 -16188 24580 -16154
rect 24633 -16188 24676 -16154
rect 27402 -16188 27444 -16154
rect 27498 -16188 27540 -16154
rect 27594 -16188 27636 -16154
rect 27690 -16188 27732 -16154
rect 27786 -16188 27828 -16154
rect 27882 -16188 27924 -16154
rect 27978 -16188 28020 -16154
rect 30746 -16188 30788 -16154
rect 30842 -16188 30884 -16154
rect 30938 -16188 30980 -16154
rect 31034 -16188 31076 -16154
rect 31130 -16188 31172 -16154
rect 31226 -16188 31268 -16154
rect 31322 -16188 31364 -16154
rect 34090 -16188 34132 -16154
rect 34186 -16188 34228 -16154
rect 34282 -16188 34324 -16154
rect 34378 -16188 34420 -16154
rect 34474 -16188 34516 -16154
rect 34570 -16188 34612 -16154
rect 34666 -16188 34708 -16154
rect 37434 -16188 37476 -16154
rect 37530 -16188 37572 -16154
rect 37626 -16188 37668 -16154
rect 37722 -16188 37764 -16154
rect 37818 -16188 37860 -16154
rect 37914 -16188 37956 -16154
rect 38010 -16188 38052 -16154
rect 14732 -16215 14825 -16197
rect 14641 -16239 14654 -16234
rect 14579 -16250 14599 -16242
rect 14632 -16250 14654 -16239
rect 13837 -16290 13846 -16279
rect 14016 -16284 14059 -16250
rect 14088 -16264 14131 -16250
rect 14160 -16264 14203 -16250
rect 14264 -16264 14278 -16253
rect 14304 -16264 14347 -16250
rect 14088 -16284 14203 -16264
rect 14275 -16284 14347 -16264
rect 14376 -16284 14491 -16250
rect 14520 -16284 14565 -16250
rect 14587 -16253 14654 -16250
rect 14576 -16264 14654 -16253
rect 13823 -16316 13846 -16305
rect 13848 -16316 13891 -16290
rect 14119 -16298 14178 -16284
rect 14275 -16298 14334 -16284
rect 14431 -16296 14490 -16284
rect 13834 -16324 13891 -16316
rect 13834 -16350 13882 -16324
rect 14402 -16333 14434 -16322
rect 14164 -16348 14178 -16337
rect 14264 -16348 14278 -16337
rect 14320 -16348 14334 -16337
rect 13837 -16373 13846 -16363
rect 13823 -16384 13846 -16373
rect 13848 -16384 13891 -16374
rect 14119 -16382 14178 -16348
rect 14275 -16382 14334 -16348
rect 14413 -16345 14465 -16333
rect 14476 -16345 14490 -16334
rect 14413 -16367 14490 -16345
rect 14431 -16379 14490 -16367
rect 13834 -16408 13891 -16384
rect 13834 -16418 13882 -16408
rect 14164 -16431 14178 -16420
rect 13536 -16463 13590 -16457
rect 13449 -16514 13463 -16494
rect 13524 -16499 13673 -16463
rect 13692 -16472 13751 -16457
rect 13690 -16491 13751 -16472
rect 13690 -16499 13737 -16491
rect 13465 -16514 13513 -16510
rect 13578 -16514 13626 -16510
rect 13153 -16544 13626 -16514
rect 12494 -16556 13128 -16546
rect 13174 -16556 13222 -16544
rect 13238 -16556 13606 -16544
rect 13627 -16555 13641 -16507
rect 13661 -16514 13675 -16507
rect 13644 -16521 13675 -16514
rect 13690 -16514 13740 -16499
rect 13746 -16514 13751 -16491
rect 13780 -16507 13785 -16438
rect 13837 -16457 13846 -16446
rect 13848 -16491 13891 -16457
rect 14119 -16465 14178 -16431
rect 13690 -16521 13822 -16514
rect 14078 -16517 14121 -16483
rect 14123 -16517 14132 -16472
rect 14200 -16519 14207 -16416
rect 14402 -16417 14434 -16406
rect 14264 -16431 14278 -16420
rect 14320 -16431 14334 -16420
rect 14234 -16472 14241 -16450
rect 14275 -16465 14334 -16431
rect 14413 -16426 14456 -16417
rect 14476 -16426 14490 -16415
rect 14413 -16451 14490 -16426
rect 14431 -16460 14490 -16451
rect 14553 -16460 14565 -16284
rect 14587 -16298 14654 -16264
rect 14587 -16322 14599 -16298
rect 14641 -16322 14654 -16298
rect 14579 -16333 14599 -16322
rect 14632 -16333 14654 -16322
rect 14587 -16337 14654 -16333
rect 14576 -16348 14654 -16337
rect 14587 -16382 14654 -16348
rect 14587 -16406 14599 -16382
rect 14641 -16406 14654 -16382
rect 14579 -16417 14599 -16406
rect 14632 -16417 14654 -16406
rect 14587 -16420 14654 -16417
rect 14576 -16431 14654 -16420
rect 14223 -16483 14278 -16472
rect 14232 -16499 14278 -16483
rect 14279 -16473 14320 -16465
rect 14279 -16499 14288 -16473
rect 14232 -16517 14288 -16499
rect 14388 -16499 14434 -16473
rect 14476 -16499 14479 -16473
rect 14553 -16496 14563 -16460
rect 14587 -16465 14654 -16431
rect 14675 -16460 14688 -16215
rect 14732 -16231 14806 -16215
rect 14831 -16216 15029 -16197
rect 17002 -16199 17009 -16196
rect 17036 -16199 17051 -16196
rect 17090 -16199 17095 -16196
rect 17124 -16199 17129 -16196
rect 15131 -16216 15145 -16208
rect 14859 -16231 14902 -16216
rect 14918 -16230 15029 -16216
rect 15071 -16224 15085 -16216
rect 15127 -16224 15145 -16216
rect 14732 -16262 14746 -16251
rect 14910 -16262 15030 -16230
rect 15082 -16240 15145 -16224
rect 15165 -16230 15179 -16208
rect 15238 -16216 15273 -16206
rect 15227 -16224 15273 -16216
rect 15283 -16224 15297 -16216
rect 15238 -16230 15297 -16224
rect 15343 -16230 15357 -16208
rect 15165 -16240 15297 -16230
rect 15309 -16240 15357 -16230
rect 15377 -16216 15391 -16208
rect 15443 -16216 15457 -16208
rect 15377 -16224 15397 -16216
rect 15439 -16224 15457 -16216
rect 15377 -16240 15391 -16224
rect 15082 -16258 15383 -16240
rect 15394 -16249 15457 -16224
rect 15477 -16230 15491 -16208
rect 15539 -16224 15553 -16216
rect 15595 -16224 15609 -16216
rect 15550 -16230 15609 -16224
rect 15655 -16230 15669 -16208
rect 15477 -16249 15525 -16230
rect 15549 -16249 15609 -16230
rect 15621 -16249 15669 -16230
rect 15689 -16216 15703 -16208
rect 15755 -16216 15769 -16208
rect 15689 -16224 15709 -16216
rect 15751 -16224 15769 -16216
rect 15689 -16249 15703 -16224
rect 15706 -16249 15769 -16224
rect 15789 -16230 15803 -16208
rect 15851 -16224 15865 -16216
rect 15907 -16224 15921 -16216
rect 15862 -16230 15921 -16224
rect 15967 -16230 15981 -16208
rect 15789 -16249 15837 -16230
rect 15861 -16249 15921 -16230
rect 15933 -16249 15981 -16230
rect 15394 -16258 15981 -16249
rect 14743 -16293 14818 -16262
rect 14910 -16264 14958 -16262
rect 14982 -16264 15030 -16262
rect 14829 -16293 14838 -16285
rect 14743 -16296 14827 -16293
rect 14756 -16327 14827 -16296
rect 14828 -16327 14871 -16293
rect 14732 -16345 14746 -16334
rect 14743 -16376 14818 -16345
rect 14743 -16379 14827 -16376
rect 14784 -16410 14827 -16379
rect 14829 -16410 14838 -16365
rect 14732 -16426 14746 -16415
rect 14743 -16460 14818 -16426
rect 14587 -16489 14599 -16465
rect 14641 -16473 14654 -16465
rect 14579 -16494 14599 -16489
rect 14619 -16494 14654 -16473
rect 14784 -16494 14827 -16460
rect 14829 -16494 14838 -16449
rect 14579 -16496 14597 -16494
rect 14232 -16519 14279 -16517
rect 14388 -16519 14479 -16499
rect 14579 -16499 14590 -16496
rect 14619 -16499 14645 -16494
rect 14579 -16500 14645 -16499
rect 14588 -16519 14645 -16500
rect 13644 -16555 13822 -16521
rect 14066 -16532 14645 -16519
rect 14042 -16534 14645 -16532
rect 14066 -16542 14645 -16534
rect 14229 -16549 14279 -16542
rect 13627 -16556 13822 -16555
rect 11261 -16565 13916 -16556
rect 11261 -16582 13391 -16565
rect 13415 -16582 13429 -16565
rect 13627 -16571 13660 -16565
rect 11238 -16740 11253 -16729
rect 11282 -16590 13391 -16582
rect 13410 -16590 13429 -16582
rect 13601 -16582 13660 -16571
rect 13661 -16582 13694 -16565
rect 11282 -16608 13429 -16590
rect 13510 -16594 13524 -16583
rect 13566 -16594 13580 -16583
rect 11282 -16740 11310 -16608
rect 11245 -16774 11310 -16740
rect 10976 -16791 11022 -16785
rect 11245 -16791 11253 -16774
rect 10976 -16813 10984 -16791
rect 10987 -16813 11022 -16791
rect 11083 -16813 11118 -16802
rect 9889 -16832 10549 -16830
rect 9512 -16995 9520 -16838
rect 8991 -17035 9035 -17029
rect 8428 -17088 8472 -17054
rect 8524 -17088 8568 -17054
rect 8620 -17088 8664 -17054
rect 9524 -17076 9534 -16838
rect 9540 -16860 9584 -16838
rect 9823 -16858 10549 -16832
rect 10590 -16832 10638 -16813
rect 10679 -16821 11245 -16813
rect 10679 -16832 11248 -16821
rect 11282 -16832 11310 -16774
rect 11316 -16624 13429 -16608
rect 11316 -16651 13391 -16624
rect 11316 -16667 11344 -16651
rect 11382 -16667 11396 -16656
rect 11466 -16657 11598 -16651
rect 11482 -16664 11598 -16657
rect 11316 -16701 11396 -16667
rect 11484 -16691 11598 -16664
rect 11638 -16667 11652 -16656
rect 11675 -16664 13391 -16651
rect 13415 -16653 13429 -16624
rect 13410 -16664 13429 -16653
rect 11675 -16667 13429 -16664
rect 11484 -16698 11564 -16691
rect 11316 -16732 11361 -16701
rect 11484 -16711 11538 -16698
rect 11543 -16711 11564 -16698
rect 11577 -16711 11598 -16691
rect 11649 -16694 13429 -16667
rect 11649 -16701 11708 -16694
rect 11805 -16698 11940 -16694
rect 11820 -16700 11940 -16698
rect 11382 -16732 11715 -16711
rect 11838 -16717 11850 -16700
rect 11823 -16732 11850 -16717
rect 11316 -16754 11344 -16732
rect 11577 -16752 11598 -16732
rect 11316 -16788 11364 -16754
rect 11388 -16771 11436 -16754
rect 11577 -16771 11625 -16754
rect 11649 -16771 11697 -16754
rect 11388 -16773 11498 -16771
rect 11388 -16788 11436 -16773
rect 11316 -16798 11344 -16788
rect 11443 -16813 11487 -16779
rect 11488 -16813 11498 -16773
rect 11577 -16773 11697 -16771
rect 11577 -16779 11625 -16773
rect 11577 -16788 11643 -16779
rect 11649 -16788 11697 -16773
rect 11721 -16788 11769 -16754
rect 11838 -16758 11850 -16732
rect 11858 -16732 11940 -16700
rect 11950 -16732 11952 -16694
rect 11961 -16701 12020 -16694
rect 12029 -16698 13429 -16694
rect 11858 -16734 11902 -16732
rect 12029 -16737 13391 -16698
rect 13415 -16714 13429 -16698
rect 12067 -16748 12081 -16737
rect 12120 -16748 12215 -16737
rect 12248 -16754 12292 -16743
rect 12379 -16748 12399 -16737
rect 12513 -16743 12527 -16737
rect 12490 -16748 12527 -16743
rect 11599 -16813 11643 -16788
rect 11725 -16798 11769 -16788
rect 11889 -16788 11937 -16754
rect 11961 -16788 12009 -16754
rect 12033 -16788 12081 -16754
rect 12201 -16777 12321 -16754
rect 12201 -16788 12249 -16777
rect 12273 -16788 12321 -16777
rect 12345 -16788 12393 -16754
rect 11889 -16798 11921 -16788
rect 12305 -16804 12308 -16798
rect 11759 -16822 11803 -16806
rect 11759 -16832 11841 -16822
rect 10590 -16847 11245 -16832
rect 10621 -16853 11245 -16847
rect 9540 -16928 9584 -16894
rect 9592 -16995 9600 -16860
rect 9823 -16874 9898 -16858
rect 9951 -16874 10549 -16858
rect 10874 -16860 10884 -16853
rect 11093 -16860 11137 -16853
rect 11138 -16860 11148 -16853
rect 11249 -16860 11293 -16832
rect 11310 -16856 11331 -16852
rect 11437 -16856 11472 -16845
rect 11616 -16856 11651 -16845
rect 11797 -16856 11841 -16832
rect 11842 -16856 11852 -16814
rect 11855 -16832 11887 -16806
rect 12339 -16809 12342 -16798
rect 11942 -16822 11952 -16814
rect 11953 -16856 11997 -16822
rect 12192 -16856 12227 -16827
rect 12370 -16845 12380 -16788
rect 12370 -16856 12385 -16845
rect 12411 -16856 12419 -16811
rect 12456 -16843 12464 -16775
rect 12490 -16809 12498 -16748
rect 12577 -16753 13391 -16737
rect 13449 -16748 13463 -16594
rect 13521 -16628 13580 -16594
rect 13601 -16590 13705 -16582
rect 13722 -16590 13751 -16565
rect 14234 -16566 14241 -16549
rect 14270 -16566 14277 -16549
rect 14590 -16566 14597 -16542
rect 14076 -16568 14616 -16566
rect 14092 -16582 14140 -16568
rect 13815 -16587 13890 -16582
rect 13601 -16603 13751 -16590
rect 13761 -16603 13785 -16594
rect 13601 -16605 13736 -16603
rect 13627 -16632 13660 -16605
rect 13661 -16624 13736 -16605
rect 13822 -16621 13896 -16587
rect 14076 -16600 14140 -16582
rect 14160 -16591 14208 -16568
rect 14228 -16591 14276 -16568
rect 14160 -16600 14276 -16591
rect 14296 -16591 14344 -16568
rect 14364 -16591 14412 -16568
rect 14432 -16591 14480 -16568
rect 14500 -16590 14548 -16568
rect 14499 -16591 14548 -16590
rect 14568 -16591 14616 -16568
rect 14784 -16577 14827 -16543
rect 14829 -16577 14838 -16532
rect 14876 -16534 14877 -16277
rect 14910 -16524 14911 -16264
rect 14918 -16285 14944 -16264
rect 15086 -16274 15383 -16258
rect 15412 -16264 15981 -16258
rect 15412 -16270 15957 -16264
rect 15131 -16281 15145 -16274
rect 14915 -16296 14938 -16285
rect 14971 -16293 14994 -16282
rect 15071 -16292 15085 -16281
rect 15127 -16292 15145 -16281
rect 14940 -16296 14994 -16293
rect 14926 -16327 14994 -16296
rect 15082 -16320 15145 -16292
rect 15165 -16320 15179 -16274
rect 15227 -16292 15241 -16281
rect 15283 -16292 15297 -16281
rect 15238 -16302 15297 -16292
rect 15082 -16325 15141 -16320
rect 15227 -16325 15297 -16302
rect 15343 -16320 15357 -16274
rect 15377 -16281 15391 -16274
rect 15443 -16277 15457 -16270
rect 15477 -16277 15491 -16270
rect 15655 -16277 15669 -16270
rect 15689 -16277 15703 -16270
rect 15755 -16277 15769 -16270
rect 15789 -16277 15803 -16270
rect 15440 -16281 15929 -16277
rect 15377 -16286 15397 -16281
rect 15377 -16292 15398 -16286
rect 15439 -16292 15929 -16281
rect 15967 -16292 15981 -16264
rect 15377 -16317 15929 -16292
rect 15343 -16325 15364 -16320
rect 15082 -16326 15192 -16325
rect 14926 -16330 14985 -16327
rect 14971 -16365 14980 -16330
rect 15127 -16336 15192 -16326
rect 15227 -16328 15364 -16325
rect 15283 -16336 15364 -16328
rect 14929 -16376 14938 -16365
rect 14971 -16376 14994 -16365
rect 15110 -16370 15225 -16336
rect 15294 -16370 15364 -16336
rect 14915 -16402 14938 -16391
rect 14940 -16402 14994 -16376
rect 14926 -16410 14994 -16402
rect 15071 -16406 15085 -16395
rect 15127 -16406 15141 -16395
rect 15227 -16406 15297 -16395
rect 15082 -16408 15141 -16406
rect 15238 -16408 15297 -16406
rect 15343 -16408 15364 -16370
rect 14926 -16436 14985 -16410
rect 14971 -16449 14980 -16436
rect 15082 -16440 15192 -16408
rect 15238 -16440 15364 -16408
rect 14929 -16459 14938 -16449
rect 14915 -16470 14938 -16459
rect 14971 -16460 14994 -16449
rect 15138 -16453 15192 -16440
rect 15294 -16453 15364 -16440
rect 14940 -16470 14994 -16460
rect 15082 -16463 15130 -16461
rect 14926 -16494 14994 -16470
rect 15071 -16474 15141 -16463
rect 15227 -16474 15297 -16463
rect 15082 -16492 15141 -16474
rect 15238 -16492 15297 -16474
rect 15343 -16492 15364 -16453
rect 14926 -16504 14985 -16494
rect 14971 -16516 14980 -16504
rect 15082 -16508 15192 -16492
rect 15238 -16508 15364 -16492
rect 15138 -16516 15192 -16508
rect 15294 -16516 15364 -16508
rect 14929 -16543 14938 -16532
rect 14969 -16542 14995 -16516
rect 14971 -16543 14995 -16542
rect 15127 -16537 15192 -16516
rect 15127 -16543 15183 -16537
rect 14940 -16577 14995 -16543
rect 14955 -16585 14995 -16577
rect 15126 -16549 15183 -16543
rect 15126 -16573 15276 -16549
rect 15292 -16573 15364 -16516
rect 13510 -16667 13524 -16656
rect 13566 -16667 13580 -16656
rect 13521 -16678 13580 -16667
rect 13627 -16673 13641 -16632
rect 13661 -16664 13694 -16624
rect 13727 -16653 13741 -16637
rect 13722 -16664 13741 -16653
rect 13661 -16673 13741 -16664
rect 13521 -16701 13590 -16678
rect 13666 -16681 13741 -16673
rect 13677 -16698 13741 -16681
rect 13536 -16723 13590 -16701
rect 13722 -16714 13741 -16698
rect 13524 -16753 13539 -16732
rect 13566 -16753 13581 -16732
rect 13722 -16753 13737 -16714
rect 13761 -16748 13775 -16637
rect 13822 -16655 13890 -16621
rect 14042 -16632 14110 -16616
rect 13822 -16656 13832 -16655
rect 13822 -16667 13836 -16656
rect 13875 -16667 13890 -16655
rect 14054 -16634 14110 -16632
rect 14054 -16666 14097 -16634
rect 14103 -16651 14110 -16634
rect 14137 -16651 14144 -16600
rect 14164 -16602 14235 -16600
rect 14278 -16602 14279 -16595
rect 14296 -16600 14871 -16591
rect 14970 -16600 14984 -16585
rect 15126 -16600 15364 -16573
rect 15377 -16326 15457 -16317
rect 15377 -16406 15398 -16326
rect 15443 -16329 15457 -16326
rect 15424 -16406 15457 -16329
rect 15477 -16363 15491 -16317
rect 15550 -16326 15609 -16317
rect 15655 -16329 15669 -16317
rect 15377 -16440 15457 -16406
rect 15377 -16461 15398 -16440
rect 15424 -16461 15457 -16440
rect 15377 -16508 15457 -16461
rect 15377 -16600 15398 -16508
rect 15424 -16600 15457 -16508
rect 15458 -16379 15491 -16363
rect 15517 -16379 15553 -16368
rect 15573 -16379 15595 -16345
rect 15650 -16379 15669 -16329
rect 15689 -16363 15703 -16317
rect 15706 -16326 15769 -16317
rect 15755 -16329 15769 -16326
rect 15738 -16345 15769 -16329
rect 15684 -16368 15703 -16363
rect 15673 -16379 15709 -16368
rect 15729 -16379 15769 -16345
rect 15789 -16363 15803 -16317
rect 15862 -16326 15921 -16317
rect 15458 -16413 15507 -16379
rect 15528 -16395 15584 -16379
rect 15608 -16395 15669 -16379
rect 15528 -16413 15669 -16395
rect 15458 -16600 15491 -16413
rect 15550 -16440 15609 -16413
rect 15517 -16462 15553 -16451
rect 15573 -16462 15595 -16440
rect 15528 -16463 15584 -16462
rect 15528 -16496 15609 -16463
rect 15550 -16508 15609 -16496
rect 15573 -16516 15595 -16508
rect 15516 -16546 15553 -16516
rect 15650 -16524 15669 -16413
rect 15684 -16413 15769 -16379
rect 15684 -16451 15703 -16413
rect 15706 -16440 15769 -16413
rect 15673 -16461 15709 -16451
rect 15729 -16461 15769 -16440
rect 15673 -16462 15769 -16461
rect 15684 -16496 15769 -16462
rect 15684 -16516 15703 -16496
rect 15706 -16508 15769 -16496
rect 15729 -16516 15769 -16508
rect 15516 -16558 15571 -16546
rect 15573 -16549 15582 -16535
rect 15650 -16549 15657 -16524
rect 15682 -16535 15709 -16516
rect 15738 -16535 15769 -16516
rect 15673 -16546 15709 -16535
rect 15682 -16549 15727 -16546
rect 15573 -16558 15727 -16549
rect 15729 -16549 15769 -16535
rect 15772 -16379 15803 -16363
rect 15829 -16379 15865 -16368
rect 15772 -16413 15821 -16379
rect 15840 -16406 15896 -16379
rect 15954 -16394 15981 -16292
rect 16001 -16216 16015 -16208
rect 16067 -16216 16081 -16208
rect 16001 -16224 16021 -16216
rect 16063 -16224 16081 -16216
rect 16001 -16281 16015 -16224
rect 16018 -16258 16081 -16224
rect 16067 -16281 16081 -16258
rect 16001 -16292 16021 -16281
rect 16063 -16292 16081 -16281
rect 16001 -16326 16015 -16292
rect 16018 -16326 16081 -16292
rect 16101 -16230 16115 -16208
rect 16163 -16224 16177 -16216
rect 16219 -16224 16233 -16216
rect 16174 -16230 16233 -16224
rect 16279 -16230 16293 -16208
rect 16101 -16264 16149 -16230
rect 16173 -16258 16233 -16230
rect 16173 -16264 16221 -16258
rect 16245 -16264 16293 -16230
rect 16101 -16326 16115 -16264
rect 16163 -16292 16177 -16281
rect 16219 -16292 16233 -16281
rect 16174 -16326 16233 -16292
rect 16279 -16326 16293 -16264
rect 16313 -16216 16327 -16208
rect 16379 -16216 16393 -16208
rect 16313 -16224 16333 -16216
rect 16375 -16224 16393 -16216
rect 16313 -16281 16327 -16224
rect 16330 -16258 16393 -16224
rect 16379 -16281 16393 -16258
rect 16313 -16292 16333 -16281
rect 16375 -16292 16393 -16281
rect 16313 -16326 16327 -16292
rect 16330 -16326 16393 -16292
rect 16413 -16230 16427 -16208
rect 16475 -16224 16489 -16216
rect 16531 -16224 16545 -16216
rect 16486 -16230 16545 -16224
rect 16591 -16230 16605 -16208
rect 16413 -16264 16461 -16230
rect 16485 -16258 16545 -16230
rect 16485 -16264 16533 -16258
rect 16557 -16264 16605 -16230
rect 16413 -16326 16427 -16264
rect 16475 -16292 16489 -16281
rect 16531 -16292 16545 -16281
rect 16486 -16326 16545 -16292
rect 16591 -16326 16605 -16264
rect 16625 -16216 16639 -16208
rect 16691 -16216 16705 -16208
rect 16625 -16224 16645 -16216
rect 16687 -16224 16705 -16216
rect 16625 -16281 16639 -16224
rect 16642 -16258 16705 -16224
rect 16691 -16281 16705 -16258
rect 16625 -16292 16645 -16281
rect 16687 -16292 16705 -16281
rect 16625 -16326 16639 -16292
rect 16642 -16326 16705 -16292
rect 15988 -16360 16669 -16326
rect 15907 -16406 15921 -16395
rect 15840 -16413 15921 -16406
rect 15772 -16549 15803 -16413
rect 15862 -16440 15921 -16413
rect 15829 -16462 15865 -16451
rect 15840 -16474 15896 -16462
rect 15907 -16474 15921 -16463
rect 15840 -16496 15921 -16474
rect 15862 -16508 15921 -16496
rect 15838 -16535 15865 -16516
rect 15829 -16546 15865 -16535
rect 15892 -16543 15895 -16516
rect 15967 -16524 15981 -16394
rect 16001 -16395 16015 -16360
rect 16067 -16395 16081 -16360
rect 16001 -16406 16021 -16395
rect 16063 -16406 16081 -16395
rect 16001 -16422 16015 -16406
rect 16018 -16416 16081 -16406
rect 16101 -16416 16115 -16360
rect 16279 -16372 16293 -16360
rect 16163 -16406 16177 -16395
rect 16219 -16406 16233 -16395
rect 16018 -16422 16077 -16416
rect 16174 -16422 16233 -16406
rect 16001 -16440 16077 -16422
rect 16001 -16456 16053 -16440
rect 16082 -16456 16125 -16422
rect 16154 -16440 16233 -16422
rect 16154 -16456 16197 -16440
rect 16001 -16463 16015 -16456
rect 16018 -16463 16066 -16461
rect 16001 -16474 16077 -16463
rect 16163 -16474 16177 -16463
rect 16219 -16474 16233 -16463
rect 15880 -16546 15895 -16543
rect 15838 -16549 15895 -16546
rect 15729 -16558 15895 -16549
rect 15516 -16580 15895 -16558
rect 15516 -16595 15729 -16580
rect 15506 -16596 15729 -16595
rect 15493 -16600 15588 -16596
rect 14320 -16602 14576 -16600
rect 14164 -16604 14576 -16602
rect 14164 -16608 14235 -16604
rect 14173 -16651 14180 -16608
rect 14278 -16633 14279 -16604
rect 14320 -16608 14576 -16604
rect 14590 -16608 14871 -16600
rect 14942 -16607 15588 -16600
rect 14499 -16624 14542 -16608
rect 14279 -16636 14320 -16633
rect 14556 -16636 14558 -16608
rect 14590 -16636 14592 -16608
rect 14259 -16638 14483 -16636
rect 14173 -16659 14201 -16651
rect 13822 -16681 13832 -16667
rect 13833 -16670 13890 -16667
rect 13833 -16701 13881 -16670
rect 14107 -16684 14201 -16659
rect 14207 -16654 14235 -16640
rect 14207 -16659 14278 -16654
rect 14632 -16659 14634 -16633
rect 14666 -16651 14871 -16608
rect 14935 -16609 15588 -16607
rect 15606 -16609 15729 -16596
rect 14935 -16618 15729 -16609
rect 15738 -16596 15895 -16580
rect 15738 -16618 15769 -16596
rect 14935 -16628 15769 -16618
rect 14901 -16642 14908 -16641
rect 14935 -16642 15252 -16628
rect 15276 -16630 15769 -16628
rect 15276 -16642 15582 -16630
rect 15586 -16642 15634 -16630
rect 15650 -16642 15669 -16630
rect 15682 -16642 15769 -16630
rect 15772 -16642 15803 -16596
rect 15805 -16600 15895 -16596
rect 15918 -16600 15966 -16596
rect 15967 -16600 15981 -16580
rect 16001 -16600 16015 -16474
rect 16018 -16508 16077 -16474
rect 16174 -16508 16233 -16474
rect 16264 -16524 16293 -16372
rect 16313 -16395 16327 -16360
rect 16379 -16395 16393 -16360
rect 16313 -16406 16333 -16395
rect 16375 -16406 16393 -16395
rect 16413 -16406 16427 -16360
rect 16475 -16395 16531 -16388
rect 16298 -16422 16327 -16406
rect 16330 -16422 16389 -16406
rect 16396 -16422 16461 -16411
rect 16475 -16414 16545 -16395
rect 16591 -16406 16605 -16360
rect 16625 -16395 16639 -16360
rect 16691 -16395 16705 -16326
rect 16625 -16406 16645 -16395
rect 16687 -16406 16705 -16395
rect 16486 -16422 16545 -16414
rect 16573 -16422 16638 -16411
rect 16298 -16440 16485 -16422
rect 16486 -16440 16557 -16422
rect 16298 -16456 16341 -16440
rect 16370 -16456 16485 -16440
rect 16514 -16456 16557 -16440
rect 16584 -16456 16638 -16422
rect 16642 -16440 16705 -16406
rect 16298 -16463 16327 -16456
rect 16330 -16463 16378 -16461
rect 16642 -16463 16690 -16461
rect 16691 -16463 16705 -16440
rect 16298 -16474 16389 -16463
rect 16475 -16474 16545 -16463
rect 16631 -16474 16705 -16463
rect 16264 -16596 16293 -16580
rect 15805 -16630 16060 -16600
rect 16117 -16609 16165 -16596
rect 16230 -16609 16293 -16596
rect 16117 -16630 16186 -16609
rect 15826 -16640 16186 -16630
rect 15826 -16642 16117 -16640
rect 16138 -16642 16186 -16640
rect 16210 -16642 16293 -16609
rect 16298 -16642 16327 -16474
rect 16330 -16508 16389 -16474
rect 16396 -16505 16461 -16494
rect 16407 -16516 16461 -16505
rect 16486 -16508 16545 -16474
rect 16573 -16505 16638 -16494
rect 16584 -16516 16638 -16505
rect 16642 -16508 16705 -16474
rect 16395 -16549 16473 -16516
rect 16550 -16549 16557 -16524
rect 16582 -16549 16639 -16516
rect 16395 -16596 16639 -16549
rect 16395 -16609 16524 -16596
rect 16542 -16600 16639 -16596
rect 16691 -16600 16705 -16508
rect 16725 -16230 16739 -16208
rect 16787 -16224 16801 -16216
rect 16811 -16224 16859 -16207
rect 16868 -16216 17247 -16199
rect 17310 -16208 17587 -16196
rect 17304 -16216 17587 -16208
rect 16798 -16230 16859 -16224
rect 16880 -16230 16934 -16216
rect 16943 -16224 17017 -16216
rect 16725 -16264 16773 -16230
rect 16797 -16241 16859 -16230
rect 16869 -16241 16934 -16230
rect 16797 -16258 16857 -16241
rect 16797 -16264 16845 -16258
rect 16869 -16264 16917 -16241
rect 16954 -16258 17017 -16224
rect 16725 -16524 16739 -16264
rect 16787 -16292 16801 -16281
rect 16843 -16292 16857 -16281
rect 16869 -16290 16934 -16279
rect 17002 -16281 17017 -16258
rect 17036 -16241 17090 -16216
rect 17099 -16224 17173 -16216
rect 17110 -16230 17173 -16224
rect 17192 -16230 17246 -16216
rect 17255 -16224 17269 -16216
rect 17284 -16222 17587 -16216
rect 17284 -16224 17478 -16222
rect 17109 -16241 17173 -16230
rect 17181 -16241 17246 -16230
rect 17036 -16264 17085 -16241
rect 17109 -16258 17169 -16241
rect 17109 -16264 17157 -16258
rect 17181 -16264 17229 -16241
rect 17266 -16242 17478 -16224
rect 18107 -16231 18150 -16197
rect 18203 -16231 18246 -16197
rect 18299 -16231 18342 -16197
rect 20269 -16207 20278 -16199
rect 20346 -16207 20353 -16191
rect 20369 -16207 20378 -16199
rect 20380 -16207 20387 -16191
rect 20434 -16199 20439 -16191
rect 17266 -16258 17329 -16242
rect 17036 -16279 17051 -16264
rect 16798 -16326 16857 -16292
rect 16880 -16324 16934 -16290
rect 16943 -16292 17017 -16281
rect 17025 -16290 17090 -16279
rect 16954 -16326 17017 -16292
rect 16869 -16374 16934 -16363
rect 16787 -16406 16801 -16395
rect 16843 -16406 16857 -16395
rect 16798 -16440 16857 -16406
rect 16880 -16408 16934 -16374
rect 17002 -16395 17017 -16326
rect 17036 -16324 17090 -16290
rect 17099 -16292 17169 -16281
rect 17181 -16290 17246 -16279
rect 17315 -16281 17329 -16258
rect 17036 -16363 17051 -16324
rect 17110 -16326 17169 -16292
rect 17192 -16324 17246 -16290
rect 17255 -16292 17269 -16281
rect 17311 -16292 17329 -16281
rect 17266 -16326 17329 -16292
rect 17025 -16374 17090 -16363
rect 17181 -16374 17246 -16363
rect 16943 -16406 17017 -16395
rect 16954 -16440 17017 -16406
rect 16869 -16457 16934 -16446
rect 16787 -16474 16801 -16463
rect 16843 -16474 16857 -16463
rect 16798 -16508 16857 -16474
rect 16880 -16491 16934 -16457
rect 17002 -16461 17017 -16440
rect 17036 -16408 17090 -16374
rect 17099 -16406 17169 -16395
rect 17036 -16446 17051 -16408
rect 17110 -16440 17169 -16406
rect 17192 -16408 17246 -16374
rect 17315 -16395 17329 -16326
rect 17255 -16406 17269 -16395
rect 17311 -16406 17329 -16395
rect 17266 -16440 17329 -16406
rect 17025 -16457 17090 -16446
rect 17181 -16457 17246 -16446
rect 16954 -16463 17017 -16461
rect 16943 -16474 17017 -16463
rect 16954 -16499 17017 -16474
rect 16943 -16507 17017 -16499
rect 16903 -16521 16917 -16507
rect 16783 -16524 16917 -16521
rect 16937 -16508 17017 -16507
rect 16937 -16516 16999 -16508
rect 16937 -16555 16951 -16516
rect 16817 -16558 16951 -16555
rect 16725 -16600 16739 -16580
rect 16542 -16609 16739 -16600
rect 16395 -16630 16739 -16609
rect 16741 -16609 16789 -16596
rect 16854 -16609 16902 -16596
rect 16945 -16605 16988 -16571
rect 16741 -16630 16810 -16609
rect 16382 -16642 16498 -16630
rect 16522 -16642 16570 -16630
rect 16582 -16642 16739 -16630
rect 14891 -16646 16739 -16642
rect 16762 -16639 16810 -16630
rect 16834 -16630 16902 -16609
rect 16834 -16639 16882 -16630
rect 16903 -16639 16917 -16632
rect 16762 -16643 16917 -16639
rect 16776 -16646 16917 -16643
rect 14891 -16651 16735 -16646
rect 14207 -16670 14334 -16659
rect 14576 -16667 14607 -16659
rect 14632 -16667 14646 -16659
rect 14207 -16684 14323 -16670
rect 14576 -16672 14646 -16667
rect 13834 -16723 13877 -16701
rect 13761 -16753 13771 -16748
rect 13832 -16753 13836 -16732
rect 14054 -16734 14097 -16700
rect 14107 -16701 14323 -16684
rect 12513 -16759 12561 -16754
rect 12500 -16788 12561 -16759
rect 12577 -16780 13893 -16753
rect 12585 -16788 12633 -16780
rect 12657 -16788 12705 -16780
rect 12500 -16793 12544 -16788
rect 12703 -16838 12747 -16804
rect 12685 -16856 12720 -16838
rect 12752 -16856 12760 -16788
rect 12786 -16856 12794 -16780
rect 12825 -16788 13017 -16780
rect 13137 -16788 13893 -16780
rect 12822 -16798 12978 -16788
rect 13148 -16796 13893 -16788
rect 14107 -16756 14164 -16701
rect 14173 -16720 14323 -16701
rect 14571 -16701 14646 -16672
rect 14345 -16720 14357 -16706
rect 14173 -16722 14320 -16720
rect 14173 -16756 14201 -16722
rect 14107 -16794 14201 -16756
rect 12822 -16809 12836 -16798
rect 12822 -16856 12830 -16809
rect 12868 -16812 12878 -16809
rect 12856 -16822 12944 -16812
rect 12856 -16832 12946 -16822
rect 12856 -16856 12864 -16832
rect 12868 -16856 12878 -16832
rect 12884 -16856 12946 -16832
rect 13167 -16856 13893 -16796
rect 14024 -16819 14073 -16794
rect 14119 -16801 14201 -16794
rect 14173 -16803 14201 -16801
rect 14075 -16819 14123 -16803
rect 14024 -16822 14123 -16819
rect 14020 -16837 14123 -16822
rect 14147 -16809 14201 -16803
rect 14207 -16756 14320 -16722
rect 14427 -16726 14434 -16725
rect 14420 -16737 14434 -16726
rect 14476 -16736 14492 -16725
rect 14438 -16737 14492 -16736
rect 14207 -16809 14235 -16756
rect 14264 -16794 14334 -16756
rect 14431 -16770 14492 -16737
rect 14431 -16771 14490 -16770
rect 14275 -16801 14334 -16794
rect 14537 -16803 14549 -16706
rect 14351 -16808 14399 -16803
rect 14147 -16823 14235 -16809
rect 14319 -16809 14399 -16808
rect 14423 -16809 14471 -16803
rect 14287 -16823 14294 -16817
rect 14319 -16819 14471 -16809
rect 14147 -16835 14219 -16823
rect 14321 -16825 14471 -16819
rect 14476 -16825 14483 -16809
rect 14147 -16837 14228 -16835
rect 14020 -16853 14086 -16837
rect 14173 -16843 14228 -16837
rect 9823 -16877 10549 -16874
rect 9626 -16980 9634 -16892
rect 9743 -16942 9787 -16908
rect 9788 -16942 9798 -16900
rect 9624 -16991 9634 -16980
rect 9626 -17025 9634 -16991
rect 9635 -17025 9679 -16991
rect 9743 -17042 9787 -17008
rect 9788 -17042 9798 -16997
rect 9823 -17044 9977 -16877
rect 10153 -16899 10549 -16877
rect 10649 -16866 11293 -16860
rect 10649 -16881 11273 -16866
rect 11297 -16878 11302 -16856
rect 11328 -16875 11376 -16856
rect 11424 -16875 11664 -16856
rect 11712 -16875 11760 -16856
rect 10077 -16925 10549 -16899
rect 10874 -16904 10884 -16881
rect 10986 -16906 11030 -16881
rect 11058 -16906 11102 -16881
rect 11130 -16906 11174 -16881
rect 11328 -16890 11760 -16875
rect 11785 -16890 12048 -16856
rect 12096 -16890 12144 -16856
rect 12171 -16890 12537 -16856
rect 12576 -16890 12624 -16856
rect 12672 -16890 12836 -16856
rect 12837 -16890 13999 -16856
rect 14020 -16865 14077 -16853
rect 14020 -16886 14079 -16865
rect 14186 -16878 14228 -16843
rect 14321 -16853 14492 -16825
rect 14495 -16837 14549 -16803
rect 14571 -16728 14592 -16701
rect 14571 -16729 14583 -16728
rect 14632 -16729 14634 -16728
rect 14571 -16740 14592 -16729
rect 14632 -16740 14648 -16729
rect 14571 -16756 14583 -16740
rect 14571 -16767 14592 -16756
rect 14594 -16767 14648 -16740
rect 14571 -16817 14583 -16767
rect 14587 -16774 14648 -16767
rect 14587 -16801 14646 -16774
rect 14632 -16809 14634 -16801
rect 14583 -16825 14592 -16821
rect 14619 -16825 14645 -16809
rect 14693 -16817 14702 -16651
rect 14727 -16659 14736 -16651
rect 14727 -16667 14746 -16659
rect 14727 -16756 14736 -16667
rect 14743 -16701 14791 -16667
rect 14849 -16691 14892 -16657
rect 14901 -16664 14908 -16651
rect 14935 -16664 14942 -16651
rect 14970 -16668 14984 -16651
rect 14917 -16680 14957 -16668
rect 14970 -16680 14984 -16669
rect 14917 -16714 14984 -16680
rect 15020 -16680 16735 -16651
rect 16937 -16668 16951 -16632
rect 17002 -16668 17017 -16508
rect 17036 -16491 17090 -16457
rect 17099 -16474 17169 -16463
rect 17036 -16637 17051 -16491
rect 17110 -16499 17169 -16474
rect 17192 -16491 17246 -16457
rect 17266 -16463 17314 -16461
rect 17315 -16463 17329 -16440
rect 17255 -16474 17329 -16463
rect 17099 -16508 17169 -16499
rect 17099 -16516 17155 -16508
rect 17215 -16524 17229 -16507
rect 17249 -16558 17263 -16507
rect 17266 -16508 17329 -16474
rect 17315 -16558 17329 -16508
rect 17349 -16264 17406 -16242
rect 17422 -16262 17478 -16242
rect 17900 -16250 17907 -16234
rect 17923 -16250 17932 -16242
rect 17934 -16250 17941 -16234
rect 17430 -16264 17478 -16262
rect 17349 -16284 17403 -16264
rect 17432 -16284 17475 -16264
rect 17504 -16284 17547 -16250
rect 17648 -16284 17691 -16250
rect 17720 -16284 17835 -16250
rect 17864 -16284 17907 -16250
rect 17349 -16524 17363 -16284
rect 17411 -16296 17425 -16285
rect 17422 -16330 17470 -16296
rect 17757 -16367 17800 -16333
rect 17411 -16402 17425 -16391
rect 17422 -16417 17470 -16402
rect 17422 -16436 17478 -16417
rect 17452 -16458 17478 -16436
rect 17411 -16470 17425 -16459
rect 17467 -16470 17481 -16459
rect 17422 -16504 17481 -16470
rect 17422 -16516 17465 -16504
rect 17356 -16534 17363 -16524
rect 17410 -16517 17465 -16516
rect 17467 -16517 17476 -16504
rect 17410 -16527 17436 -16517
rect 17410 -16542 17440 -16527
rect 17544 -16534 17551 -16416
rect 17567 -16483 17576 -16472
rect 17578 -16483 17585 -16450
rect 17614 -16483 17621 -16450
rect 17578 -16517 17621 -16483
rect 17623 -16517 17632 -16472
rect 17322 -16568 17329 -16558
rect 17424 -16559 17425 -16542
rect 17578 -16568 17585 -16517
rect 17614 -16568 17621 -16517
rect 17648 -16534 17655 -16417
rect 17745 -16458 17747 -16417
rect 17757 -16451 17800 -16417
rect 17757 -16534 17800 -16500
rect 17900 -16534 17907 -16284
rect 17934 -16284 17977 -16250
rect 18461 -16274 18504 -16240
rect 18557 -16274 18600 -16240
rect 18653 -16274 18696 -16240
rect 20160 -16241 20203 -16207
rect 20224 -16241 20278 -16207
rect 20304 -16241 20353 -16207
rect 17923 -16333 17932 -16322
rect 17934 -16333 17941 -16284
rect 18173 -16293 18182 -16285
rect 18273 -16293 18282 -16285
rect 18100 -16327 18171 -16293
rect 18172 -16327 18215 -16293
rect 18284 -16327 18327 -16293
rect 18815 -16317 18858 -16283
rect 18911 -16317 18954 -16283
rect 19007 -16317 19050 -16283
rect 19103 -16317 19146 -16283
rect 19199 -16317 19242 -16283
rect 20224 -16324 20267 -16290
rect 20269 -16324 20278 -16279
rect 17934 -16367 17977 -16333
rect 18527 -16336 18536 -16328
rect 18627 -16336 18636 -16328
rect 17923 -16417 17932 -16406
rect 17934 -16417 17941 -16367
rect 18128 -16410 18171 -16376
rect 18173 -16410 18182 -16365
rect 18273 -16376 18282 -16365
rect 18454 -16370 18525 -16336
rect 18526 -16370 18569 -16336
rect 18638 -16370 18681 -16336
rect 19363 -16360 19406 -16326
rect 19459 -16360 19502 -16326
rect 19555 -16360 19598 -16326
rect 19651 -16360 19694 -16326
rect 19747 -16360 19790 -16326
rect 19843 -16360 19886 -16326
rect 19939 -16360 19982 -16326
rect 18284 -16410 18327 -16376
rect 18917 -16379 18926 -16371
rect 18994 -16379 19001 -16363
rect 19017 -16379 19026 -16371
rect 19028 -16379 19035 -16363
rect 19082 -16371 19087 -16363
rect 17934 -16451 17977 -16417
rect 17923 -16500 17932 -16489
rect 17934 -16500 17941 -16451
rect 18128 -16494 18171 -16460
rect 18173 -16494 18182 -16449
rect 18273 -16460 18282 -16449
rect 18482 -16453 18525 -16419
rect 18527 -16453 18536 -16408
rect 18627 -16419 18636 -16408
rect 18808 -16413 18851 -16379
rect 18872 -16413 18926 -16379
rect 18952 -16413 19001 -16379
rect 18638 -16453 18681 -16419
rect 18284 -16494 18327 -16460
rect 17934 -16534 17977 -16500
rect 17934 -16568 17941 -16534
rect 17180 -16596 17240 -16587
rect 17053 -16609 17101 -16596
rect 17166 -16609 17240 -16596
rect 17272 -16608 17410 -16600
rect 17053 -16630 17122 -16609
rect 17037 -16639 17051 -16637
rect 17074 -16639 17122 -16630
rect 17037 -16643 17122 -16639
rect 17146 -16621 17240 -16609
rect 17146 -16630 17214 -16621
rect 17146 -16639 17194 -16630
rect 17215 -16639 17229 -16637
rect 17146 -16643 17229 -16639
rect 17037 -16646 17115 -16643
rect 17160 -16646 17229 -16643
rect 17249 -16639 17263 -16637
rect 17108 -16668 17115 -16646
rect 16842 -16673 16856 -16669
rect 16937 -16673 17017 -16668
rect 17098 -16669 17154 -16668
rect 17098 -16673 17168 -16669
rect 16810 -16680 17081 -16673
rect 15020 -16694 16739 -16680
rect 15081 -16710 15140 -16694
rect 15165 -16700 15296 -16694
rect 15203 -16714 15296 -16700
rect 14727 -16767 14746 -16756
rect 14803 -16767 14833 -16751
rect 14727 -16803 14736 -16767
rect 14743 -16771 14833 -16767
rect 14743 -16779 14822 -16771
rect 14743 -16801 14831 -16779
rect 14583 -16832 14645 -16825
rect 14537 -16843 14549 -16837
rect 14328 -16870 14492 -16853
rect 14592 -16865 14645 -16832
rect 14727 -16837 14781 -16803
rect 14788 -16813 14831 -16801
rect 14833 -16813 14842 -16771
rect 14727 -16843 14736 -16837
rect 14328 -16872 14483 -16870
rect 14328 -16878 14518 -16872
rect 11359 -16896 11713 -16890
rect 12183 -16895 12227 -16890
rect 12228 -16895 12238 -16890
rect 11443 -16903 11487 -16896
rect 11488 -16903 11498 -16896
rect 11599 -16903 11643 -16896
rect 11387 -16924 11685 -16903
rect 10077 -16959 10562 -16925
rect 11411 -16949 11455 -16924
rect 11483 -16949 11527 -16924
rect 11797 -16956 11841 -16922
rect 11842 -16956 11852 -16911
rect 11942 -16922 11952 -16911
rect 11953 -16956 11997 -16922
rect 10077 -16985 10549 -16959
rect 10081 -16993 10291 -16985
rect 10097 -17003 10275 -16993
rect 9636 -17078 9680 -17044
rect 9708 -17078 9752 -17044
rect 9780 -17078 9977 -17044
rect 8782 -17131 8826 -17097
rect 8878 -17131 8922 -17097
rect 8974 -17131 9018 -17097
rect 9070 -17131 9114 -17097
rect 9166 -17131 9210 -17097
rect 9823 -17114 9977 -17078
rect 9823 -17140 10007 -17114
rect 9330 -17174 9374 -17140
rect 9426 -17174 9470 -17140
rect 9522 -17174 9566 -17140
rect 9618 -17174 9662 -17140
rect 9714 -17174 9758 -17140
rect 9810 -17174 10007 -17140
rect 9823 -17200 10007 -17174
rect 10023 -17174 10133 -17050
rect 10282 -17062 10291 -17051
rect 9901 -17870 9945 -17200
rect 10023 -17228 10079 -17174
rect 9376 -17970 9754 -17936
rect 9835 -17971 9862 -17924
rect 9889 -17971 9945 -17870
rect 10035 -17971 10079 -17228
rect 10081 -17971 10090 -17174
rect 10293 -17971 10337 -17062
rect 10427 -17971 10471 -16985
rect 10680 -17002 10724 -16968
rect 10776 -17002 10820 -16968
rect 10872 -17002 10916 -16968
rect 10968 -17002 11012 -16968
rect 11064 -17002 11108 -16968
rect 11160 -17002 11204 -16968
rect 11256 -17002 11300 -16968
rect 11765 -16992 11809 -16958
rect 11837 -16992 11881 -16958
rect 12183 -16995 12227 -16961
rect 12228 -16995 12238 -16950
rect 12370 -17001 12380 -16890
rect 12481 -16895 12525 -16890
rect 12703 -16906 12747 -16890
rect 12752 -16922 12760 -16890
rect 12470 -16961 12480 -16950
rect 12786 -16956 12794 -16890
rect 12481 -16995 12525 -16961
rect 11418 -17045 11462 -17011
rect 11514 -17045 11558 -17011
rect 11610 -17045 11654 -17011
rect 12119 -17035 12163 -17001
rect 12191 -17035 12235 -17001
rect 12263 -17035 12307 -17001
rect 12335 -17029 12380 -17001
rect 12681 -17025 12725 -16991
rect 12726 -17025 12736 -16980
rect 12822 -16992 12830 -16890
rect 12856 -16995 12864 -16890
rect 12335 -17035 12379 -17029
rect 11772 -17088 11816 -17054
rect 11868 -17088 11912 -17054
rect 11964 -17088 12008 -17054
rect 12868 -17076 12878 -16890
rect 12884 -16928 12928 -16894
rect 12936 -16995 12944 -16890
rect 13167 -16891 13893 -16890
rect 13167 -16892 13965 -16891
rect 12970 -16896 13965 -16892
rect 12970 -16916 13893 -16896
rect 14219 -16899 14228 -16878
rect 14331 -16899 14446 -16878
rect 14475 -16899 14518 -16878
rect 14590 -16886 14654 -16865
rect 14788 -16868 14836 -16865
rect 14788 -16899 14842 -16868
rect 12970 -16924 13321 -16916
rect 12970 -16980 12978 -16924
rect 13075 -16942 13142 -16924
rect 13075 -16964 13132 -16942
rect 12968 -16991 12978 -16980
rect 12970 -17025 12978 -16991
rect 12979 -17025 13023 -16991
rect 13087 -17042 13131 -17008
rect 13132 -17042 13142 -16997
rect 13167 -17044 13321 -16924
rect 13422 -16919 13893 -16916
rect 14051 -16914 14719 -16899
rect 14754 -16913 14842 -16899
rect 14870 -16908 14877 -16763
rect 14904 -16840 14911 -16729
rect 14917 -16753 14942 -16714
rect 15203 -16734 15284 -16714
rect 14970 -16753 14984 -16742
rect 15070 -16750 15084 -16739
rect 15126 -16750 15140 -16739
rect 14917 -16768 14984 -16753
rect 15081 -16761 15140 -16750
rect 15226 -16742 15282 -16734
rect 14917 -16771 14998 -16768
rect 14925 -16787 14998 -16771
rect 15081 -16772 15145 -16761
rect 14944 -16813 14998 -16787
rect 15070 -16800 15145 -16772
rect 15165 -16806 15179 -16761
rect 15104 -16811 15179 -16806
rect 15226 -16787 15296 -16742
rect 14970 -16818 14984 -16813
rect 14970 -16840 14999 -16818
rect 15104 -16834 15196 -16811
rect 15226 -16814 15282 -16787
rect 15343 -16811 15364 -16694
rect 15374 -16737 16739 -16694
rect 16797 -16714 16856 -16680
rect 16869 -16689 16934 -16680
rect 16942 -16681 17012 -16680
rect 17098 -16681 17237 -16673
rect 16880 -16723 16934 -16689
rect 16953 -16710 17012 -16681
rect 17109 -16689 17237 -16681
rect 17109 -16714 17168 -16689
rect 17178 -16723 17237 -16689
rect 15377 -16750 15398 -16737
rect 15431 -16750 15457 -16737
rect 15377 -16784 15457 -16750
rect 15377 -16800 15398 -16784
rect 15431 -16793 15457 -16784
rect 15465 -16793 15491 -16737
rect 15538 -16753 15552 -16742
rect 15555 -16743 15674 -16737
rect 15573 -16753 15674 -16743
rect 15549 -16777 15674 -16753
rect 15684 -16739 15703 -16737
rect 15715 -16739 15750 -16737
rect 15755 -16739 15769 -16737
rect 15684 -16750 15708 -16739
rect 15715 -16750 15769 -16739
rect 15549 -16787 15608 -16777
rect 15573 -16793 15594 -16787
rect 15650 -16793 15669 -16777
rect 15684 -16793 15703 -16750
rect 15705 -16775 15769 -16750
rect 15789 -16775 15803 -16737
rect 15807 -16742 15906 -16737
rect 15807 -16759 15920 -16742
rect 15705 -16784 15764 -16775
rect 15715 -16793 15750 -16784
rect 15845 -16787 15920 -16759
rect 15922 -16753 16739 -16737
rect 16786 -16753 16800 -16742
rect 16842 -16753 16856 -16742
rect 16942 -16750 17012 -16739
rect 16953 -16753 17012 -16750
rect 17098 -16753 17168 -16742
rect 17215 -16753 17237 -16723
rect 15922 -16780 17237 -16753
rect 15845 -16793 15926 -16787
rect 15431 -16800 15941 -16793
rect 15287 -16822 15364 -16811
rect 15456 -16818 15941 -16800
rect 15130 -16840 15196 -16834
rect 15296 -16834 15364 -16822
rect 15477 -16834 15491 -16818
rect 15296 -16840 15353 -16834
rect 15573 -16840 15594 -16818
rect 15650 -16840 15669 -16818
rect 14904 -16868 14952 -16840
rect 14970 -16844 15024 -16840
rect 14976 -16868 15024 -16844
rect 15130 -16856 15213 -16840
rect 15130 -16859 15145 -16856
rect 14904 -16874 15024 -16868
rect 15165 -16874 15213 -16856
rect 15237 -16874 15285 -16840
rect 15296 -16844 15357 -16840
rect 15298 -16856 15357 -16844
rect 15309 -16874 15357 -16856
rect 15477 -16853 15525 -16840
rect 15549 -16853 15597 -16840
rect 15477 -16859 15597 -16853
rect 15477 -16874 15525 -16859
rect 15549 -16861 15597 -16859
rect 15528 -16874 15597 -16861
rect 15621 -16874 15669 -16840
rect 15715 -16844 15750 -16818
rect 15715 -16845 15724 -16844
rect 15715 -16853 15729 -16845
rect 15682 -16859 15729 -16853
rect 14904 -16884 14911 -16874
rect 14933 -16879 14999 -16874
rect 14942 -16908 14999 -16879
rect 15528 -16895 15571 -16874
rect 15573 -16895 15582 -16874
rect 13422 -16924 13937 -16919
rect 13422 -16925 13893 -16924
rect 13422 -16944 13937 -16925
rect 14051 -16933 14729 -16914
rect 14754 -16915 14833 -16913
rect 14851 -16915 14877 -16908
rect 14754 -16933 14877 -16915
rect 14935 -16929 15010 -16908
rect 15142 -16911 15190 -16908
rect 14051 -16939 14703 -16934
rect 13422 -16959 13906 -16944
rect 14756 -16949 14877 -16933
rect 15142 -16942 15196 -16911
rect 15266 -16942 15341 -16908
rect 15715 -16913 15729 -16859
rect 15756 -16879 15763 -16818
rect 15967 -16834 15981 -16780
rect 16001 -16800 16129 -16780
rect 16010 -16804 16129 -16800
rect 15979 -16840 15981 -16834
rect 15789 -16853 15837 -16840
rect 15861 -16853 15909 -16840
rect 15789 -16859 15909 -16853
rect 15789 -16861 15837 -16859
rect 15861 -16861 15909 -16859
rect 15789 -16874 15909 -16861
rect 15933 -16874 15981 -16840
rect 15826 -16895 15869 -16874
rect 15979 -16884 15981 -16874
rect 16013 -16906 16015 -16804
rect 16020 -16818 16129 -16804
rect 16162 -16787 16232 -16780
rect 16162 -16803 16180 -16787
rect 16279 -16788 16293 -16780
rect 16313 -16784 16393 -16780
rect 16191 -16803 16310 -16788
rect 16313 -16800 16374 -16784
rect 16379 -16800 16393 -16784
rect 16162 -16818 16310 -16803
rect 16318 -16818 16374 -16800
rect 16028 -16838 16091 -16818
rect 16028 -16844 16062 -16838
rect 16048 -16906 16091 -16872
rect 16101 -16874 16149 -16840
rect 16168 -16859 16222 -16818
rect 16173 -16874 16222 -16859
rect 16229 -16840 16272 -16826
rect 16279 -16834 16293 -16818
rect 16413 -16831 16427 -16780
rect 16474 -16818 17237 -16780
rect 17249 -16676 17271 -16639
rect 17315 -16668 17329 -16646
rect 17398 -16666 17441 -16632
rect 17447 -16668 17454 -16616
rect 17310 -16676 17329 -16668
rect 17249 -16710 17329 -16676
rect 17360 -16680 17478 -16668
rect 17481 -16680 17488 -16590
rect 17521 -16606 17530 -16595
rect 17517 -16637 17530 -16606
rect 17843 -16624 17886 -16590
rect 17249 -16750 17271 -16710
rect 17315 -16739 17329 -16710
rect 17310 -16750 17329 -16739
rect 17249 -16784 17329 -16750
rect 17249 -16800 17271 -16784
rect 17315 -16800 17329 -16784
rect 17349 -16700 17478 -16680
rect 16512 -16840 17237 -16818
rect 17349 -16834 17363 -16700
rect 17398 -16734 17478 -16700
rect 17410 -16768 17478 -16734
rect 17421 -16794 17478 -16768
rect 17365 -16818 17430 -16808
rect 17368 -16840 17430 -16818
rect 17517 -16820 17524 -16637
rect 17551 -16823 17558 -16640
rect 16229 -16860 16293 -16840
rect 16245 -16874 16293 -16860
rect 16097 -16908 16104 -16884
rect 15505 -16942 15540 -16927
rect 15715 -16942 15724 -16913
rect 16013 -16922 16104 -16908
rect 15793 -16942 15828 -16927
rect 16028 -16940 16071 -16931
rect 16131 -16942 16138 -16884
rect 16167 -16942 16174 -16884
rect 16201 -16942 16208 -16884
rect 16213 -16942 16222 -16874
rect 16281 -16884 16293 -16874
rect 16413 -16858 16461 -16840
rect 16485 -16858 17237 -16840
rect 16413 -16884 17237 -16858
rect 17358 -16844 17478 -16840
rect 17358 -16853 17419 -16844
rect 17421 -16853 17478 -16844
rect 17358 -16868 17406 -16853
rect 17430 -16868 17478 -16853
rect 17563 -16868 17572 -16637
rect 17900 -16640 17902 -16570
rect 17579 -16688 17622 -16654
rect 17934 -16674 17936 -16568
rect 18128 -16577 18171 -16543
rect 18173 -16577 18182 -16532
rect 18273 -16543 18282 -16532
rect 18482 -16537 18525 -16503
rect 18527 -16537 18536 -16492
rect 18627 -16503 18636 -16492
rect 18872 -16496 18915 -16462
rect 18917 -16496 18926 -16451
rect 18638 -16537 18681 -16503
rect 18284 -16577 18327 -16543
rect 17579 -16756 17622 -16722
rect 17631 -16823 17638 -16688
rect 18193 -16691 18236 -16657
rect 18245 -16718 18252 -16641
rect 17665 -16808 17672 -16720
rect 17782 -16770 17825 -16736
rect 17827 -16770 17836 -16728
rect 17927 -16740 17936 -16729
rect 17938 -16774 17981 -16740
rect 18279 -16752 18286 -16607
rect 18482 -16620 18525 -16586
rect 18527 -16620 18536 -16575
rect 18627 -16586 18636 -16575
rect 18872 -16580 18915 -16546
rect 18917 -16580 18926 -16535
rect 18638 -16620 18681 -16586
rect 18547 -16734 18590 -16700
rect 18599 -16761 18606 -16684
rect 17663 -16819 17672 -16808
rect 18132 -16813 18175 -16779
rect 18177 -16813 18186 -16771
rect 18277 -16779 18286 -16771
rect 18288 -16813 18331 -16779
rect 18633 -16795 18640 -16650
rect 18872 -16663 18915 -16629
rect 18917 -16663 18926 -16618
rect 18994 -16679 19001 -16413
rect 19028 -16413 19071 -16379
rect 19073 -16413 19087 -16371
rect 19017 -16462 19026 -16451
rect 19028 -16462 19035 -16413
rect 19082 -16451 19087 -16413
rect 19028 -16496 19071 -16462
rect 19073 -16496 19087 -16451
rect 19017 -16546 19026 -16535
rect 19028 -16546 19035 -16496
rect 19082 -16535 19087 -16496
rect 19028 -16580 19071 -16546
rect 19073 -16580 19087 -16535
rect 19017 -16629 19026 -16618
rect 19028 -16629 19035 -16580
rect 19082 -16618 19087 -16580
rect 19028 -16663 19071 -16629
rect 19073 -16663 19087 -16618
rect 19017 -16697 19026 -16671
rect 19028 -16713 19035 -16663
rect 18937 -16777 18980 -16743
rect 18994 -16804 18996 -16727
rect 19028 -16809 19030 -16713
rect 17665 -16853 17672 -16819
rect 17674 -16853 17717 -16819
rect 17358 -16874 17661 -16868
rect 17782 -16870 17825 -16836
rect 17827 -16870 17836 -16825
rect 17927 -16832 17936 -16821
rect 17938 -16866 17981 -16832
rect 18486 -16856 18529 -16822
rect 18531 -16856 18540 -16814
rect 18631 -16822 18640 -16814
rect 18642 -16856 18685 -16822
rect 19059 -16845 19068 -16697
rect 19082 -16713 19087 -16663
rect 19116 -16679 19121 -16363
rect 19173 -16379 19182 -16371
rect 19122 -16413 19165 -16379
rect 19184 -16413 19237 -16379
rect 19894 -16422 19901 -16406
rect 19917 -16422 19926 -16414
rect 19928 -16422 19935 -16406
rect 20224 -16408 20267 -16374
rect 20269 -16408 20278 -16363
rect 19173 -16462 19182 -16451
rect 19354 -16456 19397 -16422
rect 19426 -16456 19469 -16422
rect 19498 -16456 19541 -16422
rect 19642 -16456 19685 -16422
rect 19714 -16456 19829 -16422
rect 19858 -16456 19901 -16422
rect 19184 -16496 19227 -16462
rect 19173 -16546 19182 -16535
rect 19751 -16539 19794 -16505
rect 19184 -16580 19227 -16546
rect 19173 -16629 19182 -16618
rect 19184 -16663 19227 -16629
rect 19416 -16689 19459 -16655
rect 19461 -16689 19470 -16644
rect 19538 -16706 19545 -16588
rect 19561 -16655 19570 -16644
rect 19572 -16655 19579 -16622
rect 19608 -16655 19615 -16622
rect 19572 -16689 19615 -16655
rect 19617 -16689 19626 -16644
rect 19572 -16740 19579 -16689
rect 19608 -16740 19615 -16689
rect 19642 -16706 19649 -16589
rect 19739 -16630 19741 -16589
rect 19751 -16623 19794 -16589
rect 19751 -16706 19794 -16672
rect 19894 -16706 19901 -16456
rect 19928 -16456 19971 -16422
rect 19917 -16505 19926 -16494
rect 19928 -16505 19935 -16456
rect 20224 -16491 20267 -16457
rect 20269 -16491 20278 -16446
rect 19928 -16539 19971 -16505
rect 19917 -16589 19926 -16578
rect 19928 -16589 19935 -16539
rect 20079 -16565 20186 -16499
rect 20346 -16507 20353 -16241
rect 20380 -16241 20423 -16207
rect 20425 -16241 20439 -16199
rect 20369 -16290 20378 -16279
rect 20380 -16290 20387 -16241
rect 20434 -16279 20439 -16241
rect 20380 -16324 20423 -16290
rect 20425 -16324 20439 -16279
rect 20369 -16374 20378 -16363
rect 20380 -16374 20387 -16324
rect 20434 -16363 20439 -16324
rect 20380 -16408 20423 -16374
rect 20425 -16408 20439 -16363
rect 20369 -16457 20378 -16446
rect 20380 -16457 20387 -16408
rect 20434 -16446 20439 -16408
rect 20380 -16491 20423 -16457
rect 20425 -16491 20439 -16446
rect 20369 -16525 20378 -16499
rect 20380 -16541 20387 -16491
rect 19928 -16623 19971 -16589
rect 20289 -16605 20332 -16571
rect 19917 -16672 19926 -16661
rect 19928 -16672 19935 -16623
rect 20346 -16632 20348 -16555
rect 20380 -16637 20382 -16541
rect 19928 -16706 19971 -16672
rect 20411 -16673 20420 -16525
rect 20434 -16541 20439 -16491
rect 20468 -16507 20473 -16191
rect 20525 -16207 20534 -16199
rect 20474 -16241 20517 -16207
rect 20536 -16241 20589 -16207
rect 21451 -16231 21494 -16197
rect 21547 -16231 21590 -16197
rect 21643 -16231 21686 -16197
rect 23613 -16207 23622 -16199
rect 23690 -16207 23697 -16191
rect 23713 -16207 23722 -16199
rect 23724 -16207 23731 -16191
rect 23778 -16199 23783 -16191
rect 21244 -16250 21251 -16234
rect 21267 -16250 21276 -16242
rect 21278 -16250 21285 -16234
rect 20525 -16290 20534 -16279
rect 20704 -16284 20747 -16250
rect 20776 -16284 20819 -16250
rect 20848 -16284 20891 -16250
rect 20992 -16284 21035 -16250
rect 21064 -16284 21179 -16250
rect 21208 -16284 21251 -16250
rect 20536 -16324 20579 -16290
rect 20525 -16374 20534 -16363
rect 21101 -16367 21144 -16333
rect 20536 -16408 20579 -16374
rect 20525 -16457 20534 -16446
rect 20536 -16491 20579 -16457
rect 20766 -16517 20809 -16483
rect 20811 -16517 20820 -16472
rect 20888 -16534 20895 -16416
rect 20911 -16483 20920 -16472
rect 20922 -16483 20929 -16450
rect 20958 -16483 20965 -16450
rect 20922 -16517 20965 -16483
rect 20967 -16517 20976 -16472
rect 20922 -16568 20929 -16517
rect 20958 -16568 20965 -16517
rect 20992 -16534 20999 -16417
rect 21089 -16458 21091 -16417
rect 21101 -16451 21144 -16417
rect 21101 -16534 21144 -16500
rect 21244 -16534 21251 -16284
rect 21278 -16284 21321 -16250
rect 21805 -16274 21848 -16240
rect 21901 -16274 21944 -16240
rect 21997 -16274 22040 -16240
rect 23504 -16241 23547 -16207
rect 23568 -16241 23622 -16207
rect 23648 -16241 23697 -16207
rect 21267 -16333 21276 -16322
rect 21278 -16333 21285 -16284
rect 21517 -16293 21526 -16285
rect 21617 -16293 21626 -16285
rect 21444 -16327 21515 -16293
rect 21516 -16327 21559 -16293
rect 21628 -16327 21671 -16293
rect 22159 -16317 22202 -16283
rect 22255 -16317 22298 -16283
rect 22351 -16317 22394 -16283
rect 22447 -16317 22490 -16283
rect 22543 -16317 22586 -16283
rect 23568 -16324 23611 -16290
rect 23613 -16324 23622 -16279
rect 21278 -16367 21321 -16333
rect 21871 -16336 21880 -16328
rect 21971 -16336 21980 -16328
rect 21267 -16417 21276 -16406
rect 21278 -16417 21285 -16367
rect 21472 -16410 21515 -16376
rect 21517 -16410 21526 -16365
rect 21617 -16376 21626 -16365
rect 21798 -16370 21869 -16336
rect 21870 -16370 21913 -16336
rect 21982 -16370 22025 -16336
rect 22707 -16360 22750 -16326
rect 22803 -16360 22846 -16326
rect 22899 -16360 22942 -16326
rect 22995 -16360 23038 -16326
rect 23091 -16360 23134 -16326
rect 23187 -16360 23230 -16326
rect 23283 -16360 23326 -16326
rect 21628 -16410 21671 -16376
rect 22261 -16379 22270 -16371
rect 22338 -16379 22345 -16363
rect 22361 -16379 22370 -16371
rect 22372 -16379 22379 -16363
rect 22426 -16371 22431 -16363
rect 21278 -16451 21321 -16417
rect 21267 -16500 21276 -16489
rect 21278 -16500 21285 -16451
rect 21472 -16494 21515 -16460
rect 21517 -16494 21526 -16449
rect 21617 -16460 21626 -16449
rect 21826 -16453 21869 -16419
rect 21871 -16453 21880 -16408
rect 21971 -16419 21980 -16408
rect 22152 -16413 22195 -16379
rect 22216 -16413 22270 -16379
rect 22296 -16413 22345 -16379
rect 21982 -16453 22025 -16419
rect 21628 -16494 21671 -16460
rect 21278 -16534 21321 -16500
rect 21278 -16568 21285 -16534
rect 19928 -16740 19935 -16706
rect 20224 -16723 20267 -16689
rect 20269 -16723 20278 -16681
rect 17368 -16878 17661 -16874
rect 16229 -16928 16272 -16894
rect 16281 -16942 16288 -16884
rect 16512 -16891 17237 -16884
rect 16512 -16892 17309 -16891
rect 16315 -16918 16327 -16892
rect 16379 -16908 17309 -16892
rect 17563 -16904 17572 -16878
rect 17675 -16906 17718 -16872
rect 17747 -16906 17790 -16872
rect 17819 -16906 17862 -16872
rect 16379 -16918 17237 -16908
rect 16315 -16942 16322 -16918
rect 16432 -16942 16475 -16918
rect 16477 -16942 16486 -16918
rect 16512 -16919 17237 -16918
rect 16512 -16936 17281 -16919
rect 17338 -16934 17615 -16908
rect 18132 -16913 18175 -16879
rect 18177 -16913 18186 -16868
rect 18277 -16879 18286 -16868
rect 18288 -16913 18331 -16879
rect 18872 -16895 18915 -16861
rect 18917 -16895 18926 -16853
rect 16512 -16942 17250 -16936
rect 14851 -16955 14877 -16949
rect 14885 -16957 15073 -16942
rect 13422 -16985 13893 -16959
rect 14023 -16967 14675 -16962
rect 13425 -16993 13635 -16985
rect 13441 -17003 13619 -16993
rect 12980 -17078 13024 -17044
rect 13052 -17078 13096 -17044
rect 13124 -17078 13321 -17044
rect 12126 -17131 12170 -17097
rect 12222 -17131 12266 -17097
rect 12318 -17131 12362 -17097
rect 12414 -17131 12458 -17097
rect 12510 -17131 12554 -17097
rect 13167 -17114 13321 -17078
rect 13167 -17140 13351 -17114
rect 12674 -17174 12718 -17140
rect 12770 -17174 12814 -17140
rect 12866 -17174 12910 -17140
rect 12962 -17174 13006 -17140
rect 13058 -17174 13102 -17140
rect 13154 -17174 13351 -17140
rect 13167 -17200 13351 -17174
rect 13367 -17174 13477 -17050
rect 13626 -17062 13635 -17051
rect 13245 -17870 13289 -17200
rect 13367 -17228 13423 -17174
rect 12720 -17970 13098 -17936
rect 13179 -17971 13206 -17924
rect 13233 -17971 13289 -17870
rect 13379 -17971 13423 -17228
rect 13425 -17971 13434 -17174
rect 13637 -17971 13681 -17062
rect 13771 -17971 13815 -16985
rect 13997 -16987 14675 -16968
rect 14885 -16976 15083 -16957
rect 15108 -16964 15353 -16942
rect 15396 -16961 15444 -16942
rect 15492 -16961 15924 -16942
rect 15972 -16956 16212 -16942
rect 15108 -16976 15156 -16964
rect 15182 -16976 15296 -16964
rect 15300 -16976 15348 -16964
rect 15396 -16976 15957 -16961
rect 15972 -16966 16020 -16956
rect 16068 -16966 16212 -16956
rect 16213 -16944 16404 -16942
rect 16213 -16966 16322 -16944
rect 16356 -16966 16404 -16944
rect 16420 -16966 17268 -16942
rect 17310 -16962 17587 -16936
rect 18100 -16949 18143 -16915
rect 18172 -16949 18215 -16915
rect 18486 -16956 18529 -16922
rect 18531 -16956 18540 -16911
rect 18631 -16922 18640 -16911
rect 19059 -16913 19073 -16845
rect 19100 -16879 19107 -16811
rect 19145 -16843 19152 -16775
rect 19179 -16809 19186 -16743
rect 19189 -16793 19232 -16759
rect 19392 -16838 19435 -16804
rect 19159 -16861 19168 -16853
rect 19170 -16895 19213 -16861
rect 19392 -16906 19435 -16872
rect 18642 -16956 18685 -16922
rect 15972 -16976 17268 -16966
rect 17316 -16976 17364 -16962
rect 17378 -16968 17460 -16962
rect 17474 -16968 17556 -16962
rect 17369 -16976 17460 -16968
rect 17465 -16976 17556 -16968
rect 14885 -16982 15057 -16977
rect 14025 -17002 14068 -16987
rect 14121 -17002 14164 -16987
rect 14217 -17002 14260 -16987
rect 14313 -17002 14356 -16987
rect 14409 -17002 14452 -16987
rect 14505 -17002 14548 -16987
rect 14601 -17002 14644 -16987
rect 15110 -16992 15153 -16976
rect 15182 -16992 15225 -16976
rect 15412 -16982 15957 -16976
rect 15528 -16989 15571 -16982
rect 15573 -16989 15582 -16982
rect 15715 -16989 15724 -16982
rect 15826 -16989 15869 -16982
rect 14857 -17010 15029 -17005
rect 15440 -17010 15929 -16989
rect 14763 -17045 14806 -17011
rect 14831 -17030 15029 -17011
rect 14859 -17045 14902 -17030
rect 14955 -17045 14998 -17030
rect 15464 -17035 15507 -17010
rect 15536 -17035 15579 -17010
rect 15608 -17035 15651 -17010
rect 15680 -17029 15724 -17010
rect 16026 -17025 16069 -16991
rect 16071 -17025 16080 -16980
rect 16167 -16992 16174 -16976
rect 16201 -16995 16208 -16976
rect 15680 -17035 15723 -17029
rect 15117 -17088 15160 -17054
rect 15213 -17088 15256 -17054
rect 15309 -17088 15352 -17054
rect 16213 -17076 16222 -16976
rect 16281 -16995 16288 -16976
rect 16315 -16980 16322 -16976
rect 16313 -16991 16322 -16980
rect 16315 -17025 16322 -16991
rect 16324 -17025 16367 -16991
rect 16432 -17042 16475 -17008
rect 16477 -17042 16486 -16997
rect 16512 -17002 17237 -16976
rect 17369 -17002 17412 -16976
rect 17465 -17002 17508 -16976
rect 17561 -17002 17604 -16968
rect 17657 -17002 17700 -16968
rect 17753 -17002 17796 -16968
rect 17849 -17002 17892 -16968
rect 17945 -17002 17988 -16968
rect 18454 -16992 18497 -16958
rect 18526 -16992 18569 -16958
rect 18872 -16995 18915 -16961
rect 18917 -16995 18926 -16950
rect 19059 -17001 19068 -16913
rect 19441 -16922 19448 -16788
rect 19159 -16961 19168 -16950
rect 19475 -16956 19482 -16762
rect 19515 -16778 19524 -16767
rect 19511 -16809 19524 -16778
rect 19837 -16796 19880 -16762
rect 19170 -16995 19213 -16961
rect 16512 -17044 16665 -17002
rect 16786 -17003 16963 -17002
rect 16325 -17078 16368 -17044
rect 16397 -17078 16440 -17044
rect 16469 -17078 16665 -17044
rect 15471 -17131 15514 -17097
rect 15567 -17131 15610 -17097
rect 15663 -17131 15706 -17097
rect 15759 -17131 15802 -17097
rect 15855 -17131 15898 -17097
rect 16512 -17114 16665 -17078
rect 16512 -17140 16695 -17114
rect 16019 -17174 16062 -17140
rect 16115 -17174 16158 -17140
rect 16211 -17174 16254 -17140
rect 16307 -17174 16350 -17140
rect 16403 -17174 16446 -17140
rect 16499 -17174 16695 -17140
rect 16512 -17200 16695 -17174
rect 16712 -17174 16821 -17050
rect 16971 -17062 16979 -17051
rect 16590 -17870 16633 -17200
rect 16712 -17228 16723 -17174
rect 16065 -17970 16442 -17936
rect 16524 -17971 16550 -17924
rect 16578 -17971 16633 -17870
rect 16724 -17971 16767 -17174
rect 16770 -17971 16778 -17174
rect 16982 -17971 17025 -17062
rect 17116 -17971 17159 -17002
rect 18107 -17045 18150 -17011
rect 18203 -17045 18246 -17011
rect 18299 -17045 18342 -17011
rect 18808 -17035 18851 -17001
rect 18880 -17035 18923 -17001
rect 18952 -17035 18995 -17001
rect 19024 -17029 19068 -17001
rect 19370 -17025 19413 -16991
rect 19415 -17025 19424 -16980
rect 19511 -16992 19518 -16809
rect 19545 -16995 19552 -16812
rect 19024 -17035 19067 -17029
rect 18461 -17088 18504 -17054
rect 18557 -17088 18600 -17054
rect 18653 -17088 18696 -17054
rect 19557 -17076 19566 -16809
rect 19894 -16812 19896 -16742
rect 19928 -16819 19930 -16740
rect 20411 -16741 20425 -16673
rect 20452 -16707 20459 -16639
rect 20497 -16671 20504 -16603
rect 20531 -16637 20538 -16571
rect 20541 -16621 20584 -16587
rect 20742 -16666 20785 -16632
rect 20511 -16689 20520 -16681
rect 20522 -16723 20565 -16689
rect 20742 -16734 20785 -16700
rect 20411 -16753 20420 -16741
rect 20791 -16750 20798 -16616
rect 20186 -16819 20581 -16753
rect 20825 -16784 20832 -16590
rect 20865 -16606 20874 -16595
rect 20861 -16637 20874 -16606
rect 21187 -16624 21230 -16590
rect 19573 -16860 19616 -16826
rect 19922 -16830 19941 -16819
rect 19922 -16832 19930 -16830
rect 19573 -16928 19616 -16894
rect 19625 -16995 19632 -16860
rect 19856 -16874 19930 -16832
rect 19984 -16874 20581 -16819
rect 20720 -16853 20763 -16819
rect 20765 -16853 20774 -16808
rect 20861 -16820 20868 -16637
rect 20895 -16823 20902 -16640
rect 19856 -16877 20581 -16874
rect 19659 -16980 19666 -16892
rect 19776 -16942 19819 -16908
rect 19821 -16942 19830 -16900
rect 19657 -16991 19666 -16980
rect 19659 -17025 19666 -16991
rect 19668 -17025 19711 -16991
rect 19776 -17042 19819 -17008
rect 19821 -17042 19830 -16997
rect 19856 -17044 20009 -16877
rect 20186 -16899 20581 -16877
rect 20110 -16925 20581 -16899
rect 20907 -16904 20916 -16637
rect 21244 -16640 21246 -16570
rect 20923 -16688 20966 -16654
rect 21278 -16674 21280 -16568
rect 21472 -16577 21515 -16543
rect 21517 -16577 21526 -16532
rect 21617 -16543 21626 -16532
rect 21826 -16537 21869 -16503
rect 21871 -16537 21880 -16492
rect 21971 -16503 21980 -16492
rect 22216 -16496 22259 -16462
rect 22261 -16496 22270 -16451
rect 21982 -16537 22025 -16503
rect 21628 -16577 21671 -16543
rect 20923 -16756 20966 -16722
rect 20975 -16823 20982 -16688
rect 21537 -16691 21580 -16657
rect 21589 -16718 21596 -16641
rect 21009 -16808 21016 -16720
rect 21126 -16770 21169 -16736
rect 21171 -16770 21180 -16728
rect 21271 -16740 21280 -16729
rect 21282 -16774 21325 -16740
rect 21623 -16752 21630 -16607
rect 21826 -16620 21869 -16586
rect 21871 -16620 21880 -16575
rect 21971 -16586 21980 -16575
rect 22216 -16580 22259 -16546
rect 22261 -16580 22270 -16535
rect 21982 -16620 22025 -16586
rect 21891 -16734 21934 -16700
rect 21943 -16761 21950 -16684
rect 21007 -16819 21016 -16808
rect 21476 -16813 21519 -16779
rect 21521 -16813 21530 -16771
rect 21621 -16779 21630 -16771
rect 21632 -16813 21675 -16779
rect 21977 -16795 21984 -16650
rect 22216 -16663 22259 -16629
rect 22261 -16663 22270 -16618
rect 22338 -16679 22345 -16413
rect 22372 -16413 22415 -16379
rect 22417 -16413 22431 -16371
rect 22361 -16462 22370 -16451
rect 22372 -16462 22379 -16413
rect 22426 -16451 22431 -16413
rect 22372 -16496 22415 -16462
rect 22417 -16496 22431 -16451
rect 22361 -16546 22370 -16535
rect 22372 -16546 22379 -16496
rect 22426 -16535 22431 -16496
rect 22372 -16580 22415 -16546
rect 22417 -16580 22431 -16535
rect 22361 -16629 22370 -16618
rect 22372 -16629 22379 -16580
rect 22426 -16618 22431 -16580
rect 22372 -16663 22415 -16629
rect 22417 -16663 22431 -16618
rect 22361 -16697 22370 -16671
rect 22372 -16713 22379 -16663
rect 22281 -16777 22324 -16743
rect 22338 -16804 22340 -16727
rect 22372 -16809 22374 -16713
rect 21009 -16853 21016 -16819
rect 21018 -16853 21061 -16819
rect 21126 -16870 21169 -16836
rect 21171 -16870 21180 -16825
rect 21271 -16832 21280 -16821
rect 21282 -16866 21325 -16832
rect 21830 -16856 21873 -16822
rect 21875 -16856 21884 -16814
rect 21975 -16822 21984 -16814
rect 21986 -16856 22029 -16822
rect 22403 -16845 22412 -16697
rect 22426 -16713 22431 -16663
rect 22460 -16679 22465 -16363
rect 22517 -16379 22526 -16371
rect 22466 -16413 22509 -16379
rect 22528 -16413 22581 -16379
rect 23238 -16422 23245 -16406
rect 23261 -16422 23270 -16414
rect 23272 -16422 23279 -16406
rect 23568 -16408 23611 -16374
rect 23613 -16408 23622 -16363
rect 22517 -16462 22526 -16451
rect 22698 -16456 22741 -16422
rect 22770 -16456 22813 -16422
rect 22842 -16456 22885 -16422
rect 22986 -16456 23029 -16422
rect 23058 -16456 23173 -16422
rect 23202 -16456 23245 -16422
rect 22528 -16496 22571 -16462
rect 22517 -16546 22526 -16535
rect 23095 -16539 23138 -16505
rect 22528 -16580 22571 -16546
rect 22517 -16629 22526 -16618
rect 22528 -16663 22571 -16629
rect 22760 -16689 22803 -16655
rect 22805 -16689 22814 -16644
rect 22882 -16706 22889 -16588
rect 22905 -16655 22914 -16644
rect 22916 -16655 22923 -16622
rect 22952 -16655 22959 -16622
rect 22916 -16689 22959 -16655
rect 22961 -16689 22970 -16644
rect 22916 -16740 22923 -16689
rect 22952 -16740 22959 -16689
rect 22986 -16706 22993 -16589
rect 23083 -16630 23085 -16589
rect 23095 -16623 23138 -16589
rect 23095 -16706 23138 -16672
rect 23238 -16706 23245 -16456
rect 23272 -16456 23315 -16422
rect 23261 -16505 23270 -16494
rect 23272 -16505 23279 -16456
rect 23568 -16491 23611 -16457
rect 23613 -16491 23622 -16446
rect 23272 -16539 23315 -16505
rect 23261 -16589 23270 -16578
rect 23272 -16589 23279 -16539
rect 23423 -16565 23530 -16499
rect 23690 -16507 23697 -16241
rect 23724 -16241 23767 -16207
rect 23769 -16241 23783 -16199
rect 23713 -16290 23722 -16279
rect 23724 -16290 23731 -16241
rect 23778 -16279 23783 -16241
rect 23724 -16324 23767 -16290
rect 23769 -16324 23783 -16279
rect 23713 -16374 23722 -16363
rect 23724 -16374 23731 -16324
rect 23778 -16363 23783 -16324
rect 23724 -16408 23767 -16374
rect 23769 -16408 23783 -16363
rect 23713 -16457 23722 -16446
rect 23724 -16457 23731 -16408
rect 23778 -16446 23783 -16408
rect 23724 -16491 23767 -16457
rect 23769 -16491 23783 -16446
rect 23713 -16525 23722 -16499
rect 23724 -16541 23731 -16491
rect 23272 -16623 23315 -16589
rect 23633 -16605 23676 -16571
rect 23261 -16672 23270 -16661
rect 23272 -16672 23279 -16623
rect 23690 -16632 23692 -16555
rect 23724 -16637 23726 -16541
rect 23272 -16706 23315 -16672
rect 23755 -16673 23764 -16525
rect 23778 -16541 23783 -16491
rect 23812 -16507 23817 -16191
rect 23869 -16207 23878 -16199
rect 23818 -16241 23861 -16207
rect 23880 -16241 23933 -16207
rect 24795 -16231 24838 -16197
rect 24891 -16231 24934 -16197
rect 24987 -16231 25030 -16197
rect 26958 -16207 26966 -16199
rect 27035 -16207 27041 -16191
rect 27058 -16207 27066 -16199
rect 27069 -16207 27075 -16191
rect 24588 -16250 24595 -16234
rect 24611 -16250 24620 -16242
rect 24622 -16250 24629 -16234
rect 23869 -16290 23878 -16279
rect 24048 -16284 24091 -16250
rect 24120 -16284 24163 -16250
rect 24192 -16284 24235 -16250
rect 24336 -16284 24379 -16250
rect 24408 -16284 24523 -16250
rect 24552 -16284 24595 -16250
rect 23880 -16324 23923 -16290
rect 23869 -16374 23878 -16363
rect 24445 -16367 24488 -16333
rect 23880 -16408 23923 -16374
rect 23869 -16457 23878 -16446
rect 23880 -16491 23923 -16457
rect 24110 -16517 24153 -16483
rect 24155 -16517 24164 -16472
rect 24232 -16534 24239 -16416
rect 24255 -16483 24264 -16472
rect 24266 -16483 24273 -16450
rect 24302 -16483 24309 -16450
rect 24266 -16517 24309 -16483
rect 24311 -16517 24320 -16472
rect 24266 -16568 24273 -16517
rect 24302 -16568 24309 -16517
rect 24336 -16534 24343 -16417
rect 24433 -16458 24435 -16417
rect 24445 -16451 24488 -16417
rect 24445 -16534 24488 -16500
rect 24588 -16534 24595 -16284
rect 24622 -16284 24665 -16250
rect 25149 -16274 25192 -16240
rect 25245 -16274 25288 -16240
rect 25341 -16274 25384 -16240
rect 26849 -16241 26891 -16207
rect 26913 -16241 26966 -16207
rect 26993 -16241 27041 -16207
rect 24611 -16333 24620 -16322
rect 24622 -16333 24629 -16284
rect 24861 -16293 24870 -16285
rect 24961 -16293 24970 -16285
rect 24788 -16327 24859 -16293
rect 24860 -16327 24903 -16293
rect 24972 -16327 25015 -16293
rect 25503 -16317 25546 -16283
rect 25599 -16317 25642 -16283
rect 25695 -16317 25738 -16283
rect 25791 -16317 25834 -16283
rect 25887 -16317 25930 -16283
rect 26913 -16324 26955 -16290
rect 26958 -16324 26966 -16279
rect 24622 -16367 24665 -16333
rect 25215 -16336 25224 -16328
rect 25315 -16336 25324 -16328
rect 24611 -16417 24620 -16406
rect 24622 -16417 24629 -16367
rect 24816 -16410 24859 -16376
rect 24861 -16410 24870 -16365
rect 24961 -16376 24970 -16365
rect 25142 -16370 25213 -16336
rect 25214 -16370 25257 -16336
rect 25326 -16370 25369 -16336
rect 26051 -16360 26094 -16326
rect 26147 -16360 26190 -16326
rect 26243 -16360 26286 -16326
rect 26339 -16360 26382 -16326
rect 26435 -16360 26478 -16326
rect 26531 -16360 26574 -16326
rect 26627 -16360 26670 -16326
rect 24972 -16410 25015 -16376
rect 25605 -16379 25614 -16371
rect 25682 -16379 25689 -16363
rect 25705 -16379 25714 -16371
rect 25716 -16379 25723 -16363
rect 25770 -16371 25775 -16363
rect 24622 -16451 24665 -16417
rect 24611 -16500 24620 -16489
rect 24622 -16500 24629 -16451
rect 24816 -16494 24859 -16460
rect 24861 -16494 24870 -16449
rect 24961 -16460 24970 -16449
rect 25170 -16453 25213 -16419
rect 25215 -16453 25224 -16408
rect 25315 -16419 25324 -16408
rect 25496 -16413 25539 -16379
rect 25560 -16413 25614 -16379
rect 25640 -16413 25689 -16379
rect 25326 -16453 25369 -16419
rect 24972 -16494 25015 -16460
rect 24622 -16534 24665 -16500
rect 24622 -16568 24629 -16534
rect 23272 -16740 23279 -16706
rect 23568 -16723 23611 -16689
rect 23613 -16723 23622 -16681
rect 21019 -16906 21062 -16872
rect 21091 -16906 21134 -16872
rect 21163 -16906 21206 -16872
rect 21476 -16913 21519 -16879
rect 21521 -16913 21530 -16868
rect 21621 -16879 21630 -16868
rect 21632 -16913 21675 -16879
rect 22216 -16895 22259 -16861
rect 22261 -16895 22270 -16853
rect 20110 -16959 20594 -16925
rect 21444 -16949 21487 -16915
rect 21516 -16949 21559 -16915
rect 21830 -16956 21873 -16922
rect 21875 -16956 21884 -16911
rect 21975 -16922 21984 -16911
rect 22403 -16913 22417 -16845
rect 22444 -16879 22451 -16811
rect 22489 -16843 22496 -16775
rect 22523 -16809 22530 -16743
rect 22533 -16793 22576 -16759
rect 22736 -16838 22779 -16804
rect 22503 -16861 22512 -16853
rect 22514 -16895 22557 -16861
rect 22736 -16906 22779 -16872
rect 21986 -16956 22029 -16922
rect 20110 -16985 20581 -16959
rect 20114 -16993 20323 -16985
rect 20130 -17003 20307 -16993
rect 19669 -17078 19712 -17044
rect 19741 -17078 19784 -17044
rect 19813 -17078 20009 -17044
rect 18815 -17131 18858 -17097
rect 18911 -17131 18954 -17097
rect 19007 -17131 19050 -17097
rect 19103 -17131 19146 -17097
rect 19199 -17131 19242 -17097
rect 19856 -17114 20009 -17078
rect 19856 -17140 20039 -17114
rect 19363 -17174 19406 -17140
rect 19459 -17174 19502 -17140
rect 19555 -17174 19598 -17140
rect 19651 -17174 19694 -17140
rect 19747 -17174 19790 -17140
rect 19843 -17174 20039 -17140
rect 19856 -17200 20039 -17174
rect 20056 -17174 20165 -17050
rect 20315 -17062 20323 -17051
rect 19934 -17870 19977 -17200
rect 20056 -17228 20067 -17174
rect 19409 -17970 19786 -17936
rect 19868 -17971 19894 -17924
rect 19922 -17971 19977 -17870
rect 20068 -17971 20111 -17174
rect 20114 -17971 20122 -17174
rect 20326 -17971 20369 -17062
rect 20460 -17971 20503 -16985
rect 20713 -17002 20756 -16968
rect 20809 -17002 20852 -16968
rect 20905 -17002 20948 -16968
rect 21001 -17002 21044 -16968
rect 21097 -17002 21140 -16968
rect 21193 -17002 21236 -16968
rect 21289 -17002 21332 -16968
rect 21798 -16992 21841 -16958
rect 21870 -16992 21913 -16958
rect 22216 -16995 22259 -16961
rect 22261 -16995 22270 -16950
rect 22403 -17001 22412 -16913
rect 22785 -16922 22792 -16788
rect 22503 -16961 22512 -16950
rect 22819 -16956 22826 -16762
rect 22859 -16778 22868 -16767
rect 22855 -16809 22868 -16778
rect 23181 -16796 23224 -16762
rect 22514 -16995 22557 -16961
rect 21451 -17045 21494 -17011
rect 21547 -17045 21590 -17011
rect 21643 -17045 21686 -17011
rect 22152 -17035 22195 -17001
rect 22224 -17035 22267 -17001
rect 22296 -17035 22339 -17001
rect 22368 -17029 22412 -17001
rect 22714 -17025 22757 -16991
rect 22759 -17025 22768 -16980
rect 22855 -16992 22862 -16809
rect 22889 -16995 22896 -16812
rect 22368 -17035 22411 -17029
rect 21805 -17088 21848 -17054
rect 21901 -17088 21944 -17054
rect 21997 -17088 22040 -17054
rect 22901 -17076 22910 -16809
rect 23238 -16812 23240 -16742
rect 23272 -16819 23274 -16740
rect 23755 -16741 23769 -16673
rect 23796 -16707 23803 -16639
rect 23841 -16671 23848 -16603
rect 23875 -16637 23882 -16571
rect 23885 -16621 23928 -16587
rect 24086 -16666 24129 -16632
rect 23855 -16689 23864 -16681
rect 23866 -16723 23909 -16689
rect 24086 -16734 24129 -16700
rect 23755 -16753 23764 -16741
rect 24135 -16750 24142 -16616
rect 23530 -16819 23925 -16753
rect 24169 -16784 24176 -16590
rect 24209 -16606 24218 -16595
rect 24205 -16637 24218 -16606
rect 24531 -16624 24574 -16590
rect 22917 -16860 22960 -16826
rect 23266 -16830 23285 -16819
rect 23266 -16832 23274 -16830
rect 22917 -16928 22960 -16894
rect 22969 -16995 22976 -16860
rect 23200 -16874 23274 -16832
rect 23328 -16874 23925 -16819
rect 24064 -16853 24107 -16819
rect 24109 -16853 24118 -16808
rect 24205 -16820 24212 -16637
rect 24239 -16823 24246 -16640
rect 23200 -16877 23925 -16874
rect 23003 -16980 23010 -16892
rect 23120 -16942 23163 -16908
rect 23165 -16942 23174 -16900
rect 23001 -16991 23010 -16980
rect 23003 -17025 23010 -16991
rect 23012 -17025 23055 -16991
rect 23120 -17042 23163 -17008
rect 23165 -17042 23174 -16997
rect 23200 -17044 23353 -16877
rect 23530 -16899 23925 -16877
rect 23454 -16925 23925 -16899
rect 24251 -16904 24260 -16637
rect 24588 -16640 24590 -16570
rect 24267 -16688 24310 -16654
rect 24622 -16674 24624 -16568
rect 24816 -16577 24859 -16543
rect 24861 -16577 24870 -16532
rect 24961 -16543 24970 -16532
rect 25170 -16537 25213 -16503
rect 25215 -16537 25224 -16492
rect 25315 -16503 25324 -16492
rect 25560 -16496 25603 -16462
rect 25605 -16496 25614 -16451
rect 25326 -16537 25369 -16503
rect 24972 -16577 25015 -16543
rect 24267 -16756 24310 -16722
rect 24319 -16823 24326 -16688
rect 24881 -16691 24924 -16657
rect 24933 -16718 24940 -16641
rect 24353 -16808 24360 -16720
rect 24470 -16770 24513 -16736
rect 24515 -16770 24524 -16728
rect 24615 -16740 24624 -16729
rect 24626 -16774 24669 -16740
rect 24967 -16752 24974 -16607
rect 25170 -16620 25213 -16586
rect 25215 -16620 25224 -16575
rect 25315 -16586 25324 -16575
rect 25560 -16580 25603 -16546
rect 25605 -16580 25614 -16535
rect 25326 -16620 25369 -16586
rect 25235 -16734 25278 -16700
rect 25287 -16761 25294 -16684
rect 24351 -16819 24360 -16808
rect 24820 -16813 24863 -16779
rect 24865 -16813 24874 -16771
rect 24965 -16779 24974 -16771
rect 24976 -16813 25019 -16779
rect 25321 -16795 25328 -16650
rect 25560 -16663 25603 -16629
rect 25605 -16663 25614 -16618
rect 25682 -16679 25689 -16413
rect 25716 -16413 25759 -16379
rect 25761 -16413 25775 -16371
rect 25705 -16462 25714 -16451
rect 25716 -16462 25723 -16413
rect 25770 -16451 25775 -16413
rect 25716 -16496 25759 -16462
rect 25761 -16496 25775 -16451
rect 25705 -16546 25714 -16535
rect 25716 -16546 25723 -16496
rect 25770 -16535 25775 -16496
rect 25716 -16580 25759 -16546
rect 25761 -16580 25775 -16535
rect 25705 -16629 25714 -16618
rect 25716 -16629 25723 -16580
rect 25770 -16618 25775 -16580
rect 25716 -16663 25759 -16629
rect 25761 -16663 25775 -16618
rect 25705 -16697 25714 -16671
rect 25716 -16713 25723 -16663
rect 25625 -16777 25668 -16743
rect 25682 -16804 25684 -16727
rect 25716 -16809 25718 -16713
rect 24353 -16853 24360 -16819
rect 24362 -16853 24405 -16819
rect 24470 -16870 24513 -16836
rect 24515 -16870 24524 -16825
rect 24615 -16832 24624 -16821
rect 24626 -16866 24669 -16832
rect 25174 -16856 25217 -16822
rect 25219 -16856 25228 -16814
rect 25319 -16822 25328 -16814
rect 25330 -16856 25373 -16822
rect 25747 -16845 25756 -16697
rect 25770 -16713 25775 -16663
rect 25804 -16679 25809 -16363
rect 25861 -16379 25870 -16371
rect 25810 -16413 25853 -16379
rect 25872 -16413 25925 -16379
rect 26582 -16422 26589 -16406
rect 26605 -16422 26614 -16414
rect 26616 -16422 26623 -16406
rect 26913 -16408 26955 -16374
rect 26958 -16408 26966 -16363
rect 25861 -16462 25870 -16451
rect 26042 -16456 26085 -16422
rect 26114 -16456 26157 -16422
rect 26186 -16456 26229 -16422
rect 26330 -16456 26373 -16422
rect 26402 -16456 26517 -16422
rect 26546 -16456 26589 -16422
rect 25872 -16496 25915 -16462
rect 25861 -16546 25870 -16535
rect 26439 -16539 26482 -16505
rect 25872 -16580 25915 -16546
rect 25861 -16629 25870 -16618
rect 25872 -16663 25915 -16629
rect 26104 -16689 26147 -16655
rect 26149 -16689 26158 -16644
rect 26226 -16706 26233 -16588
rect 26249 -16655 26258 -16644
rect 26260 -16655 26267 -16622
rect 26296 -16655 26303 -16622
rect 26260 -16689 26303 -16655
rect 26305 -16689 26314 -16644
rect 26260 -16740 26267 -16689
rect 26296 -16740 26303 -16689
rect 26330 -16706 26337 -16589
rect 26427 -16630 26429 -16589
rect 26439 -16623 26482 -16589
rect 26439 -16706 26482 -16672
rect 26582 -16706 26589 -16456
rect 26616 -16456 26659 -16422
rect 26605 -16505 26614 -16494
rect 26616 -16505 26623 -16456
rect 26913 -16491 26955 -16457
rect 26958 -16491 26966 -16446
rect 26616 -16539 26659 -16505
rect 26605 -16589 26614 -16578
rect 26616 -16589 26623 -16539
rect 26767 -16565 26875 -16499
rect 27035 -16507 27041 -16241
rect 27069 -16241 27111 -16207
rect 27114 -16241 27122 -16199
rect 27058 -16290 27066 -16279
rect 27069 -16290 27075 -16241
rect 27069 -16324 27111 -16290
rect 27114 -16324 27122 -16279
rect 27058 -16374 27066 -16363
rect 27069 -16374 27075 -16324
rect 27069 -16408 27111 -16374
rect 27114 -16408 27122 -16363
rect 27058 -16457 27066 -16446
rect 27069 -16457 27075 -16408
rect 27069 -16491 27111 -16457
rect 27114 -16491 27122 -16446
rect 27058 -16525 27066 -16499
rect 27069 -16541 27075 -16491
rect 26616 -16623 26659 -16589
rect 26978 -16605 27020 -16571
rect 26605 -16672 26614 -16661
rect 26616 -16672 26623 -16623
rect 27035 -16632 27036 -16555
rect 27069 -16637 27070 -16541
rect 26616 -16706 26659 -16672
rect 27100 -16673 27108 -16525
rect 27123 -16541 27127 -16191
rect 27157 -16507 27161 -16191
rect 27214 -16207 27222 -16199
rect 27163 -16241 27205 -16207
rect 27225 -16241 27277 -16207
rect 28140 -16231 28182 -16197
rect 28236 -16231 28278 -16197
rect 28332 -16231 28374 -16197
rect 30302 -16207 30310 -16199
rect 30379 -16207 30385 -16191
rect 30402 -16207 30410 -16199
rect 30413 -16207 30419 -16191
rect 27933 -16250 27939 -16234
rect 27956 -16250 27964 -16242
rect 27967 -16250 27973 -16234
rect 27214 -16290 27222 -16279
rect 27393 -16284 27435 -16250
rect 27465 -16284 27507 -16250
rect 27537 -16284 27579 -16250
rect 27681 -16284 27723 -16250
rect 27753 -16284 27867 -16250
rect 27897 -16284 27939 -16250
rect 27225 -16324 27267 -16290
rect 27214 -16374 27222 -16363
rect 27790 -16367 27832 -16333
rect 27225 -16408 27267 -16374
rect 27214 -16457 27222 -16446
rect 27225 -16491 27267 -16457
rect 27455 -16517 27497 -16483
rect 27500 -16517 27508 -16472
rect 27577 -16534 27583 -16416
rect 27600 -16483 27608 -16472
rect 27611 -16483 27617 -16450
rect 27647 -16483 27653 -16450
rect 27611 -16517 27653 -16483
rect 27656 -16517 27664 -16472
rect 27611 -16568 27617 -16517
rect 27647 -16568 27653 -16517
rect 27681 -16534 27687 -16417
rect 27778 -16458 27779 -16417
rect 27790 -16451 27832 -16417
rect 27790 -16534 27832 -16500
rect 27933 -16534 27939 -16284
rect 27967 -16284 28009 -16250
rect 28494 -16274 28536 -16240
rect 28590 -16274 28632 -16240
rect 28686 -16274 28728 -16240
rect 30193 -16241 30235 -16207
rect 30257 -16241 30310 -16207
rect 30337 -16241 30385 -16207
rect 27956 -16333 27964 -16322
rect 27967 -16333 27973 -16284
rect 28206 -16293 28214 -16285
rect 28306 -16293 28314 -16285
rect 28133 -16327 28203 -16293
rect 28205 -16327 28247 -16293
rect 28317 -16327 28359 -16293
rect 28848 -16317 28890 -16283
rect 28944 -16317 28986 -16283
rect 29040 -16317 29082 -16283
rect 29136 -16317 29178 -16283
rect 29232 -16317 29274 -16283
rect 30257 -16324 30299 -16290
rect 30302 -16324 30310 -16279
rect 27967 -16367 28009 -16333
rect 28560 -16336 28568 -16328
rect 28660 -16336 28668 -16328
rect 27956 -16417 27964 -16406
rect 27967 -16417 27973 -16367
rect 28161 -16410 28203 -16376
rect 28206 -16410 28214 -16365
rect 28306 -16376 28314 -16365
rect 28487 -16370 28557 -16336
rect 28559 -16370 28601 -16336
rect 28671 -16370 28713 -16336
rect 29396 -16360 29438 -16326
rect 29492 -16360 29534 -16326
rect 29588 -16360 29630 -16326
rect 29684 -16360 29726 -16326
rect 29780 -16360 29822 -16326
rect 29876 -16360 29918 -16326
rect 29972 -16360 30014 -16326
rect 28317 -16410 28359 -16376
rect 28950 -16379 28958 -16371
rect 29027 -16379 29033 -16363
rect 29050 -16379 29058 -16371
rect 29061 -16379 29067 -16363
rect 27967 -16451 28009 -16417
rect 27956 -16500 27964 -16489
rect 27967 -16500 27973 -16451
rect 28161 -16494 28203 -16460
rect 28206 -16494 28214 -16449
rect 28306 -16460 28314 -16449
rect 28515 -16453 28557 -16419
rect 28560 -16453 28568 -16408
rect 28660 -16419 28668 -16408
rect 28841 -16413 28883 -16379
rect 28905 -16413 28958 -16379
rect 28985 -16413 29033 -16379
rect 28671 -16453 28713 -16419
rect 28317 -16494 28359 -16460
rect 27967 -16534 28009 -16500
rect 27967 -16568 27973 -16534
rect 26616 -16740 26623 -16706
rect 26913 -16723 26955 -16689
rect 26958 -16723 26966 -16681
rect 24363 -16906 24406 -16872
rect 24435 -16906 24478 -16872
rect 24507 -16906 24550 -16872
rect 24820 -16913 24863 -16879
rect 24865 -16913 24874 -16868
rect 24965 -16879 24974 -16868
rect 24976 -16913 25019 -16879
rect 25560 -16895 25603 -16861
rect 25605 -16895 25614 -16853
rect 23454 -16959 23938 -16925
rect 24788 -16949 24831 -16915
rect 24860 -16949 24903 -16915
rect 25174 -16956 25217 -16922
rect 25219 -16956 25228 -16911
rect 25319 -16922 25328 -16911
rect 25747 -16913 25761 -16845
rect 25788 -16879 25795 -16811
rect 25833 -16843 25840 -16775
rect 25867 -16809 25874 -16743
rect 25877 -16793 25920 -16759
rect 26080 -16838 26123 -16804
rect 25847 -16861 25856 -16853
rect 25858 -16895 25901 -16861
rect 26080 -16906 26123 -16872
rect 25330 -16956 25373 -16922
rect 23454 -16985 23925 -16959
rect 23458 -16993 23667 -16985
rect 23474 -17003 23651 -16993
rect 23013 -17078 23056 -17044
rect 23085 -17078 23128 -17044
rect 23157 -17078 23353 -17044
rect 22159 -17131 22202 -17097
rect 22255 -17131 22298 -17097
rect 22351 -17131 22394 -17097
rect 22447 -17131 22490 -17097
rect 22543 -17131 22586 -17097
rect 23200 -17114 23353 -17078
rect 23200 -17140 23383 -17114
rect 22707 -17174 22750 -17140
rect 22803 -17174 22846 -17140
rect 22899 -17174 22942 -17140
rect 22995 -17174 23038 -17140
rect 23091 -17174 23134 -17140
rect 23187 -17174 23383 -17140
rect 23200 -17200 23383 -17174
rect 23400 -17174 23509 -17050
rect 23659 -17062 23667 -17051
rect 23278 -17870 23321 -17200
rect 23400 -17228 23411 -17174
rect 22753 -17970 23130 -17936
rect 23212 -17971 23238 -17924
rect 23266 -17971 23321 -17870
rect 23412 -17971 23455 -17174
rect 23458 -17971 23466 -17174
rect 23670 -17971 23713 -17062
rect 23804 -17971 23847 -16985
rect 24057 -17002 24100 -16968
rect 24153 -17002 24196 -16968
rect 24249 -17002 24292 -16968
rect 24345 -17002 24388 -16968
rect 24441 -17002 24484 -16968
rect 24537 -17002 24580 -16968
rect 24633 -17002 24676 -16968
rect 25142 -16992 25185 -16958
rect 25214 -16992 25257 -16958
rect 25560 -16995 25603 -16961
rect 25605 -16995 25614 -16950
rect 25747 -17001 25756 -16913
rect 26129 -16922 26136 -16788
rect 25847 -16961 25856 -16950
rect 26163 -16956 26170 -16762
rect 26203 -16778 26212 -16767
rect 26199 -16809 26212 -16778
rect 26525 -16796 26568 -16762
rect 25858 -16995 25901 -16961
rect 24795 -17045 24838 -17011
rect 24891 -17045 24934 -17011
rect 24987 -17045 25030 -17011
rect 25496 -17035 25539 -17001
rect 25568 -17035 25611 -17001
rect 25640 -17035 25683 -17001
rect 25712 -17029 25756 -17001
rect 26058 -17025 26101 -16991
rect 26103 -17025 26112 -16980
rect 26199 -16992 26206 -16809
rect 26233 -16995 26240 -16812
rect 25712 -17035 25755 -17029
rect 25149 -17088 25192 -17054
rect 25245 -17088 25288 -17054
rect 25341 -17088 25384 -17054
rect 26245 -17076 26254 -16809
rect 26582 -16812 26584 -16742
rect 26616 -16819 26618 -16740
rect 27100 -16741 27113 -16673
rect 27141 -16707 27147 -16639
rect 27186 -16671 27192 -16603
rect 27220 -16637 27226 -16571
rect 27230 -16621 27272 -16587
rect 27431 -16666 27473 -16632
rect 27200 -16689 27208 -16681
rect 27211 -16723 27253 -16689
rect 27431 -16734 27473 -16700
rect 27100 -16753 27108 -16741
rect 27480 -16750 27486 -16616
rect 26875 -16819 27269 -16753
rect 27514 -16784 27520 -16590
rect 27554 -16606 27562 -16595
rect 27550 -16637 27562 -16606
rect 27876 -16624 27918 -16590
rect 26261 -16860 26304 -16826
rect 26610 -16830 26629 -16819
rect 26610 -16832 26618 -16830
rect 26261 -16928 26304 -16894
rect 26313 -16995 26320 -16860
rect 26544 -16874 26618 -16832
rect 26673 -16874 27269 -16819
rect 27409 -16853 27451 -16819
rect 27454 -16853 27462 -16808
rect 27550 -16820 27556 -16637
rect 27584 -16823 27590 -16640
rect 26544 -16877 27269 -16874
rect 26347 -16980 26354 -16892
rect 26464 -16942 26507 -16908
rect 26509 -16942 26518 -16900
rect 26345 -16991 26354 -16980
rect 26347 -17025 26354 -16991
rect 26356 -17025 26399 -16991
rect 26464 -17042 26507 -17008
rect 26509 -17042 26518 -16997
rect 26544 -17044 26697 -16877
rect 26875 -16899 27269 -16877
rect 26799 -16925 27269 -16899
rect 27596 -16904 27604 -16637
rect 27933 -16640 27934 -16570
rect 27612 -16688 27654 -16654
rect 27967 -16674 27968 -16568
rect 28161 -16577 28203 -16543
rect 28206 -16577 28214 -16532
rect 28306 -16543 28314 -16532
rect 28515 -16537 28557 -16503
rect 28560 -16537 28568 -16492
rect 28660 -16503 28668 -16492
rect 28905 -16496 28947 -16462
rect 28950 -16496 28958 -16451
rect 28671 -16537 28713 -16503
rect 28317 -16577 28359 -16543
rect 27612 -16756 27654 -16722
rect 27664 -16823 27670 -16688
rect 28226 -16691 28268 -16657
rect 28278 -16718 28284 -16641
rect 27698 -16808 27704 -16720
rect 27815 -16770 27857 -16736
rect 27860 -16770 27868 -16728
rect 27960 -16740 27968 -16729
rect 27971 -16774 28013 -16740
rect 28312 -16752 28318 -16607
rect 28515 -16620 28557 -16586
rect 28560 -16620 28568 -16575
rect 28660 -16586 28668 -16575
rect 28905 -16580 28947 -16546
rect 28950 -16580 28958 -16535
rect 28671 -16620 28713 -16586
rect 28580 -16734 28622 -16700
rect 28632 -16761 28638 -16684
rect 27696 -16819 27704 -16808
rect 28165 -16813 28207 -16779
rect 28210 -16813 28218 -16771
rect 28310 -16779 28318 -16771
rect 28321 -16813 28363 -16779
rect 28666 -16795 28672 -16650
rect 28905 -16663 28947 -16629
rect 28950 -16663 28958 -16618
rect 29027 -16679 29033 -16413
rect 29061 -16413 29103 -16379
rect 29106 -16413 29114 -16371
rect 29050 -16462 29058 -16451
rect 29061 -16462 29067 -16413
rect 29061 -16496 29103 -16462
rect 29106 -16496 29114 -16451
rect 29050 -16546 29058 -16535
rect 29061 -16546 29067 -16496
rect 29061 -16580 29103 -16546
rect 29106 -16580 29114 -16535
rect 29050 -16629 29058 -16618
rect 29061 -16629 29067 -16580
rect 29061 -16663 29103 -16629
rect 29106 -16663 29114 -16618
rect 29050 -16697 29058 -16671
rect 29061 -16713 29067 -16663
rect 28970 -16777 29012 -16743
rect 29027 -16804 29028 -16727
rect 29061 -16809 29062 -16713
rect 27698 -16853 27704 -16819
rect 27707 -16853 27749 -16819
rect 27815 -16870 27857 -16836
rect 27860 -16870 27868 -16825
rect 27960 -16832 27968 -16821
rect 27971 -16866 28013 -16832
rect 28519 -16856 28561 -16822
rect 28564 -16856 28572 -16814
rect 28664 -16822 28672 -16814
rect 28675 -16856 28717 -16822
rect 29092 -16845 29100 -16697
rect 29115 -16713 29119 -16363
rect 29149 -16679 29153 -16363
rect 29206 -16379 29214 -16371
rect 29155 -16413 29197 -16379
rect 29217 -16413 29269 -16379
rect 29927 -16422 29933 -16406
rect 29950 -16422 29958 -16414
rect 29961 -16422 29967 -16406
rect 30257 -16408 30299 -16374
rect 30302 -16408 30310 -16363
rect 29206 -16462 29214 -16451
rect 29387 -16456 29429 -16422
rect 29459 -16456 29501 -16422
rect 29531 -16456 29573 -16422
rect 29675 -16456 29717 -16422
rect 29747 -16456 29861 -16422
rect 29891 -16456 29933 -16422
rect 29217 -16496 29259 -16462
rect 29206 -16546 29214 -16535
rect 29784 -16539 29826 -16505
rect 29217 -16580 29259 -16546
rect 29206 -16629 29214 -16618
rect 29217 -16663 29259 -16629
rect 29449 -16689 29491 -16655
rect 29494 -16689 29502 -16644
rect 29571 -16706 29577 -16588
rect 29594 -16655 29602 -16644
rect 29605 -16655 29611 -16622
rect 29641 -16655 29647 -16622
rect 29605 -16689 29647 -16655
rect 29650 -16689 29658 -16644
rect 29605 -16740 29611 -16689
rect 29641 -16740 29647 -16689
rect 29675 -16706 29681 -16589
rect 29772 -16630 29773 -16589
rect 29784 -16623 29826 -16589
rect 29784 -16706 29826 -16672
rect 29927 -16706 29933 -16456
rect 29961 -16456 30003 -16422
rect 29950 -16505 29958 -16494
rect 29961 -16505 29967 -16456
rect 30257 -16491 30299 -16457
rect 30302 -16491 30310 -16446
rect 29961 -16539 30003 -16505
rect 29950 -16589 29958 -16578
rect 29961 -16589 29967 -16539
rect 30111 -16565 30219 -16499
rect 30379 -16507 30385 -16241
rect 30413 -16241 30455 -16207
rect 30458 -16241 30466 -16199
rect 30402 -16290 30410 -16279
rect 30413 -16290 30419 -16241
rect 30413 -16324 30455 -16290
rect 30458 -16324 30466 -16279
rect 30402 -16374 30410 -16363
rect 30413 -16374 30419 -16324
rect 30413 -16408 30455 -16374
rect 30458 -16408 30466 -16363
rect 30402 -16457 30410 -16446
rect 30413 -16457 30419 -16408
rect 30413 -16491 30455 -16457
rect 30458 -16491 30466 -16446
rect 30402 -16525 30410 -16499
rect 30413 -16541 30419 -16491
rect 29961 -16623 30003 -16589
rect 30322 -16605 30364 -16571
rect 29950 -16672 29958 -16661
rect 29961 -16672 29967 -16623
rect 30379 -16632 30380 -16555
rect 30413 -16637 30414 -16541
rect 29961 -16706 30003 -16672
rect 30444 -16673 30452 -16525
rect 30467 -16541 30471 -16191
rect 30501 -16507 30505 -16191
rect 30558 -16207 30566 -16199
rect 30507 -16241 30549 -16207
rect 30569 -16241 30621 -16207
rect 31484 -16231 31526 -16197
rect 31580 -16231 31622 -16197
rect 31676 -16231 31718 -16197
rect 33646 -16207 33654 -16199
rect 33723 -16207 33729 -16191
rect 33746 -16207 33754 -16199
rect 33757 -16207 33763 -16191
rect 31277 -16250 31283 -16234
rect 31300 -16250 31308 -16242
rect 31311 -16250 31317 -16234
rect 30558 -16290 30566 -16279
rect 30737 -16284 30779 -16250
rect 30809 -16284 30851 -16250
rect 30881 -16284 30923 -16250
rect 31025 -16284 31067 -16250
rect 31097 -16284 31211 -16250
rect 31241 -16284 31283 -16250
rect 30569 -16324 30611 -16290
rect 30558 -16374 30566 -16363
rect 31134 -16367 31176 -16333
rect 30569 -16408 30611 -16374
rect 30558 -16457 30566 -16446
rect 30569 -16491 30611 -16457
rect 30799 -16517 30841 -16483
rect 30844 -16517 30852 -16472
rect 30921 -16534 30927 -16416
rect 30944 -16483 30952 -16472
rect 30955 -16483 30961 -16450
rect 30991 -16483 30997 -16450
rect 30955 -16517 30997 -16483
rect 31000 -16517 31008 -16472
rect 30955 -16568 30961 -16517
rect 30991 -16568 30997 -16517
rect 31025 -16534 31031 -16417
rect 31122 -16458 31123 -16417
rect 31134 -16451 31176 -16417
rect 31134 -16534 31176 -16500
rect 31277 -16534 31283 -16284
rect 31311 -16284 31353 -16250
rect 31838 -16274 31880 -16240
rect 31934 -16274 31976 -16240
rect 32030 -16274 32072 -16240
rect 33537 -16241 33579 -16207
rect 33601 -16241 33654 -16207
rect 33681 -16241 33729 -16207
rect 31300 -16333 31308 -16322
rect 31311 -16333 31317 -16284
rect 31550 -16293 31558 -16285
rect 31650 -16293 31658 -16285
rect 31477 -16327 31547 -16293
rect 31549 -16327 31591 -16293
rect 31661 -16327 31703 -16293
rect 32192 -16317 32234 -16283
rect 32288 -16317 32330 -16283
rect 32384 -16317 32426 -16283
rect 32480 -16317 32522 -16283
rect 32576 -16317 32618 -16283
rect 33601 -16324 33643 -16290
rect 33646 -16324 33654 -16279
rect 31311 -16367 31353 -16333
rect 31904 -16336 31912 -16328
rect 32004 -16336 32012 -16328
rect 31300 -16417 31308 -16406
rect 31311 -16417 31317 -16367
rect 31505 -16410 31547 -16376
rect 31550 -16410 31558 -16365
rect 31650 -16376 31658 -16365
rect 31831 -16370 31901 -16336
rect 31903 -16370 31945 -16336
rect 32015 -16370 32057 -16336
rect 32740 -16360 32782 -16326
rect 32836 -16360 32878 -16326
rect 32932 -16360 32974 -16326
rect 33028 -16360 33070 -16326
rect 33124 -16360 33166 -16326
rect 33220 -16360 33262 -16326
rect 33316 -16360 33358 -16326
rect 31661 -16410 31703 -16376
rect 32294 -16379 32302 -16371
rect 32371 -16379 32377 -16363
rect 32394 -16379 32402 -16371
rect 32405 -16379 32411 -16363
rect 31311 -16451 31353 -16417
rect 31300 -16500 31308 -16489
rect 31311 -16500 31317 -16451
rect 31505 -16494 31547 -16460
rect 31550 -16494 31558 -16449
rect 31650 -16460 31658 -16449
rect 31859 -16453 31901 -16419
rect 31904 -16453 31912 -16408
rect 32004 -16419 32012 -16408
rect 32185 -16413 32227 -16379
rect 32249 -16413 32302 -16379
rect 32329 -16413 32377 -16379
rect 32015 -16453 32057 -16419
rect 31661 -16494 31703 -16460
rect 31311 -16534 31353 -16500
rect 31311 -16568 31317 -16534
rect 29961 -16740 29967 -16706
rect 30257 -16723 30299 -16689
rect 30302 -16723 30310 -16681
rect 27708 -16906 27750 -16872
rect 27780 -16906 27822 -16872
rect 27852 -16906 27894 -16872
rect 28165 -16913 28207 -16879
rect 28210 -16913 28218 -16868
rect 28310 -16879 28318 -16868
rect 28321 -16913 28363 -16879
rect 28905 -16895 28947 -16861
rect 28950 -16895 28958 -16853
rect 26799 -16959 27282 -16925
rect 28133 -16949 28175 -16915
rect 28205 -16949 28247 -16915
rect 28519 -16956 28561 -16922
rect 28564 -16956 28572 -16911
rect 28664 -16922 28672 -16911
rect 29092 -16913 29105 -16845
rect 29133 -16879 29139 -16811
rect 29178 -16843 29184 -16775
rect 29212 -16809 29218 -16743
rect 29222 -16793 29264 -16759
rect 29425 -16838 29467 -16804
rect 29192 -16861 29200 -16853
rect 29203 -16895 29245 -16861
rect 29425 -16906 29467 -16872
rect 28675 -16956 28717 -16922
rect 26799 -16985 27269 -16959
rect 26802 -16993 27011 -16985
rect 26818 -17003 26995 -16993
rect 26357 -17078 26400 -17044
rect 26429 -17078 26472 -17044
rect 26501 -17078 26697 -17044
rect 25503 -17131 25546 -17097
rect 25599 -17131 25642 -17097
rect 25695 -17131 25738 -17097
rect 25791 -17131 25834 -17097
rect 25887 -17131 25930 -17097
rect 26544 -17114 26697 -17078
rect 26544 -17140 26727 -17114
rect 26051 -17174 26094 -17140
rect 26147 -17174 26190 -17140
rect 26243 -17174 26286 -17140
rect 26339 -17174 26382 -17140
rect 26435 -17174 26478 -17140
rect 26531 -17174 26727 -17140
rect 26544 -17200 26727 -17174
rect 26744 -17174 26853 -17050
rect 27003 -17062 27011 -17051
rect 26622 -17870 26665 -17200
rect 26744 -17228 26755 -17174
rect 26097 -17970 26474 -17936
rect 26556 -17971 26582 -17924
rect 26610 -17971 26665 -17870
rect 26756 -17971 26799 -17174
rect 26802 -17971 26810 -17174
rect 27014 -17971 27057 -17062
rect 27148 -17971 27191 -16985
rect 27402 -17002 27444 -16968
rect 27498 -17002 27540 -16968
rect 27594 -17002 27636 -16968
rect 27690 -17002 27732 -16968
rect 27786 -17002 27828 -16968
rect 27882 -17002 27924 -16968
rect 27978 -17002 28020 -16968
rect 28487 -16992 28529 -16958
rect 28559 -16992 28601 -16958
rect 28905 -16995 28947 -16961
rect 28950 -16995 28958 -16950
rect 29092 -17001 29100 -16913
rect 29474 -16922 29480 -16788
rect 29192 -16961 29200 -16950
rect 29508 -16956 29514 -16762
rect 29548 -16778 29556 -16767
rect 29544 -16809 29556 -16778
rect 29870 -16796 29912 -16762
rect 29203 -16995 29245 -16961
rect 28140 -17045 28182 -17011
rect 28236 -17045 28278 -17011
rect 28332 -17045 28374 -17011
rect 28841 -17035 28883 -17001
rect 28913 -17035 28955 -17001
rect 28985 -17035 29027 -17001
rect 29057 -17029 29100 -17001
rect 29403 -17025 29445 -16991
rect 29448 -17025 29456 -16980
rect 29544 -16992 29550 -16809
rect 29578 -16995 29584 -16812
rect 29057 -17035 29099 -17029
rect 28494 -17088 28536 -17054
rect 28590 -17088 28632 -17054
rect 28686 -17088 28728 -17054
rect 29590 -17076 29598 -16809
rect 29927 -16812 29928 -16742
rect 29961 -16819 29962 -16740
rect 30444 -16741 30457 -16673
rect 30485 -16707 30491 -16639
rect 30530 -16671 30536 -16603
rect 30564 -16637 30570 -16571
rect 30574 -16621 30616 -16587
rect 30775 -16666 30817 -16632
rect 30544 -16689 30552 -16681
rect 30555 -16723 30597 -16689
rect 30775 -16734 30817 -16700
rect 30444 -16753 30452 -16741
rect 30824 -16750 30830 -16616
rect 30219 -16819 30613 -16753
rect 30858 -16784 30864 -16590
rect 30898 -16606 30906 -16595
rect 30894 -16637 30906 -16606
rect 31220 -16624 31262 -16590
rect 29606 -16860 29648 -16826
rect 29955 -16830 29973 -16819
rect 29955 -16832 29962 -16830
rect 29606 -16928 29648 -16894
rect 29658 -16995 29664 -16860
rect 29889 -16874 29962 -16832
rect 30017 -16874 30613 -16819
rect 30753 -16853 30795 -16819
rect 30798 -16853 30806 -16808
rect 30894 -16820 30900 -16637
rect 30928 -16823 30934 -16640
rect 29889 -16877 30613 -16874
rect 29692 -16980 29698 -16892
rect 29809 -16942 29851 -16908
rect 29854 -16942 29862 -16900
rect 29690 -16991 29698 -16980
rect 29692 -17025 29698 -16991
rect 29701 -17025 29743 -16991
rect 29809 -17042 29851 -17008
rect 29854 -17042 29862 -16997
rect 29702 -17078 29744 -17044
rect 29774 -17078 29816 -17044
rect 29846 -17078 29888 -17044
rect 28848 -17131 28890 -17097
rect 28944 -17131 28986 -17097
rect 29040 -17131 29082 -17097
rect 29136 -17131 29178 -17097
rect 29232 -17131 29274 -17097
rect 29889 -17114 30041 -16877
rect 30219 -16899 30613 -16877
rect 30143 -16925 30613 -16899
rect 30940 -16904 30948 -16637
rect 31277 -16640 31278 -16570
rect 30956 -16688 30998 -16654
rect 31311 -16674 31312 -16568
rect 31505 -16577 31547 -16543
rect 31550 -16577 31558 -16532
rect 31650 -16543 31658 -16532
rect 31859 -16537 31901 -16503
rect 31904 -16537 31912 -16492
rect 32004 -16503 32012 -16492
rect 32249 -16496 32291 -16462
rect 32294 -16496 32302 -16451
rect 32015 -16537 32057 -16503
rect 31661 -16577 31703 -16543
rect 30956 -16756 30998 -16722
rect 31008 -16823 31014 -16688
rect 31570 -16691 31612 -16657
rect 31622 -16718 31628 -16641
rect 31042 -16808 31048 -16720
rect 31159 -16770 31201 -16736
rect 31204 -16770 31212 -16728
rect 31304 -16740 31312 -16729
rect 31315 -16774 31357 -16740
rect 31656 -16752 31662 -16607
rect 31859 -16620 31901 -16586
rect 31904 -16620 31912 -16575
rect 32004 -16586 32012 -16575
rect 32249 -16580 32291 -16546
rect 32294 -16580 32302 -16535
rect 32015 -16620 32057 -16586
rect 31924 -16734 31966 -16700
rect 31976 -16761 31982 -16684
rect 31040 -16819 31048 -16808
rect 31509 -16813 31551 -16779
rect 31554 -16813 31562 -16771
rect 31654 -16779 31662 -16771
rect 31665 -16813 31707 -16779
rect 32010 -16795 32016 -16650
rect 32249 -16663 32291 -16629
rect 32294 -16663 32302 -16618
rect 32371 -16679 32377 -16413
rect 32405 -16413 32447 -16379
rect 32450 -16413 32458 -16371
rect 32394 -16462 32402 -16451
rect 32405 -16462 32411 -16413
rect 32405 -16496 32447 -16462
rect 32450 -16496 32458 -16451
rect 32394 -16546 32402 -16535
rect 32405 -16546 32411 -16496
rect 32405 -16580 32447 -16546
rect 32450 -16580 32458 -16535
rect 32394 -16629 32402 -16618
rect 32405 -16629 32411 -16580
rect 32405 -16663 32447 -16629
rect 32450 -16663 32458 -16618
rect 32394 -16697 32402 -16671
rect 32405 -16713 32411 -16663
rect 32314 -16777 32356 -16743
rect 32371 -16804 32372 -16727
rect 32405 -16809 32406 -16713
rect 31042 -16853 31048 -16819
rect 31051 -16853 31093 -16819
rect 31159 -16870 31201 -16836
rect 31204 -16870 31212 -16825
rect 31304 -16832 31312 -16821
rect 31315 -16866 31357 -16832
rect 31863 -16856 31905 -16822
rect 31908 -16856 31916 -16814
rect 32008 -16822 32016 -16814
rect 32019 -16856 32061 -16822
rect 32436 -16845 32444 -16697
rect 32459 -16713 32463 -16363
rect 32493 -16679 32497 -16363
rect 32550 -16379 32558 -16371
rect 32499 -16413 32541 -16379
rect 32561 -16413 32613 -16379
rect 33271 -16422 33277 -16406
rect 33294 -16422 33302 -16414
rect 33305 -16422 33311 -16406
rect 33601 -16408 33643 -16374
rect 33646 -16408 33654 -16363
rect 32550 -16462 32558 -16451
rect 32731 -16456 32773 -16422
rect 32803 -16456 32845 -16422
rect 32875 -16456 32917 -16422
rect 33019 -16456 33061 -16422
rect 33091 -16456 33205 -16422
rect 33235 -16456 33277 -16422
rect 32561 -16496 32603 -16462
rect 32550 -16546 32558 -16535
rect 33128 -16539 33170 -16505
rect 32561 -16580 32603 -16546
rect 32550 -16629 32558 -16618
rect 32561 -16663 32603 -16629
rect 32793 -16689 32835 -16655
rect 32838 -16689 32846 -16644
rect 32915 -16706 32921 -16588
rect 32938 -16655 32946 -16644
rect 32949 -16655 32955 -16622
rect 32985 -16655 32991 -16622
rect 32949 -16689 32991 -16655
rect 32994 -16689 33002 -16644
rect 32949 -16740 32955 -16689
rect 32985 -16740 32991 -16689
rect 33019 -16706 33025 -16589
rect 33116 -16630 33117 -16589
rect 33128 -16623 33170 -16589
rect 33128 -16706 33170 -16672
rect 33271 -16706 33277 -16456
rect 33305 -16456 33347 -16422
rect 33294 -16505 33302 -16494
rect 33305 -16505 33311 -16456
rect 33601 -16491 33643 -16457
rect 33646 -16491 33654 -16446
rect 33305 -16539 33347 -16505
rect 33294 -16589 33302 -16578
rect 33305 -16589 33311 -16539
rect 33455 -16565 33563 -16499
rect 33723 -16507 33729 -16241
rect 33757 -16241 33799 -16207
rect 33802 -16241 33810 -16199
rect 33746 -16290 33754 -16279
rect 33757 -16290 33763 -16241
rect 33757 -16324 33799 -16290
rect 33802 -16324 33810 -16279
rect 33746 -16374 33754 -16363
rect 33757 -16374 33763 -16324
rect 33757 -16408 33799 -16374
rect 33802 -16408 33810 -16363
rect 33746 -16457 33754 -16446
rect 33757 -16457 33763 -16408
rect 33757 -16491 33799 -16457
rect 33802 -16491 33810 -16446
rect 33746 -16525 33754 -16499
rect 33757 -16541 33763 -16491
rect 33305 -16623 33347 -16589
rect 33666 -16605 33708 -16571
rect 33294 -16672 33302 -16661
rect 33305 -16672 33311 -16623
rect 33723 -16632 33724 -16555
rect 33757 -16637 33758 -16541
rect 33305 -16706 33347 -16672
rect 33788 -16673 33796 -16525
rect 33811 -16541 33815 -16191
rect 33845 -16507 33849 -16191
rect 33902 -16207 33910 -16199
rect 33851 -16241 33893 -16207
rect 33913 -16241 33965 -16207
rect 34828 -16231 34870 -16197
rect 34924 -16231 34966 -16197
rect 35020 -16231 35062 -16197
rect 36990 -16207 36998 -16199
rect 37067 -16207 37073 -16191
rect 37090 -16207 37098 -16199
rect 37101 -16207 37107 -16191
rect 34621 -16250 34627 -16234
rect 34644 -16250 34652 -16242
rect 34655 -16250 34661 -16234
rect 33902 -16290 33910 -16279
rect 34081 -16284 34123 -16250
rect 34153 -16284 34195 -16250
rect 34225 -16284 34267 -16250
rect 34369 -16284 34411 -16250
rect 34441 -16284 34555 -16250
rect 34585 -16284 34627 -16250
rect 33913 -16324 33955 -16290
rect 33902 -16374 33910 -16363
rect 34478 -16367 34520 -16333
rect 33913 -16408 33955 -16374
rect 33902 -16457 33910 -16446
rect 33913 -16491 33955 -16457
rect 34143 -16517 34185 -16483
rect 34188 -16517 34196 -16472
rect 34265 -16534 34271 -16416
rect 34288 -16483 34296 -16472
rect 34299 -16483 34305 -16450
rect 34335 -16483 34341 -16450
rect 34299 -16517 34341 -16483
rect 34344 -16517 34352 -16472
rect 34299 -16568 34305 -16517
rect 34335 -16568 34341 -16517
rect 34369 -16534 34375 -16417
rect 34466 -16458 34467 -16417
rect 34478 -16451 34520 -16417
rect 34478 -16534 34520 -16500
rect 34621 -16534 34627 -16284
rect 34655 -16284 34697 -16250
rect 35182 -16274 35224 -16240
rect 35278 -16274 35320 -16240
rect 35374 -16274 35416 -16240
rect 36881 -16241 36923 -16207
rect 36945 -16241 36998 -16207
rect 37025 -16241 37073 -16207
rect 34644 -16333 34652 -16322
rect 34655 -16333 34661 -16284
rect 34894 -16293 34902 -16285
rect 34994 -16293 35002 -16285
rect 34821 -16327 34891 -16293
rect 34893 -16327 34935 -16293
rect 35005 -16327 35047 -16293
rect 35536 -16317 35578 -16283
rect 35632 -16317 35674 -16283
rect 35728 -16317 35770 -16283
rect 35824 -16317 35866 -16283
rect 35920 -16317 35962 -16283
rect 36945 -16324 36987 -16290
rect 36990 -16324 36998 -16279
rect 34655 -16367 34697 -16333
rect 35248 -16336 35256 -16328
rect 35348 -16336 35356 -16328
rect 34644 -16417 34652 -16406
rect 34655 -16417 34661 -16367
rect 34849 -16410 34891 -16376
rect 34894 -16410 34902 -16365
rect 34994 -16376 35002 -16365
rect 35175 -16370 35245 -16336
rect 35247 -16370 35289 -16336
rect 35359 -16370 35401 -16336
rect 36084 -16360 36126 -16326
rect 36180 -16360 36222 -16326
rect 36276 -16360 36318 -16326
rect 36372 -16360 36414 -16326
rect 36468 -16360 36510 -16326
rect 36564 -16360 36606 -16326
rect 36660 -16360 36702 -16326
rect 35005 -16410 35047 -16376
rect 35638 -16379 35646 -16371
rect 35715 -16379 35721 -16363
rect 35738 -16379 35746 -16371
rect 35749 -16379 35755 -16363
rect 34655 -16451 34697 -16417
rect 34644 -16500 34652 -16489
rect 34655 -16500 34661 -16451
rect 34849 -16494 34891 -16460
rect 34894 -16494 34902 -16449
rect 34994 -16460 35002 -16449
rect 35203 -16453 35245 -16419
rect 35248 -16453 35256 -16408
rect 35348 -16419 35356 -16408
rect 35529 -16413 35571 -16379
rect 35593 -16413 35646 -16379
rect 35673 -16413 35721 -16379
rect 35359 -16453 35401 -16419
rect 35005 -16494 35047 -16460
rect 34655 -16534 34697 -16500
rect 34655 -16568 34661 -16534
rect 33305 -16740 33311 -16706
rect 33601 -16723 33643 -16689
rect 33646 -16723 33654 -16681
rect 31052 -16906 31094 -16872
rect 31124 -16906 31166 -16872
rect 31196 -16906 31238 -16872
rect 31509 -16913 31551 -16879
rect 31554 -16913 31562 -16868
rect 31654 -16879 31662 -16868
rect 31665 -16913 31707 -16879
rect 32249 -16895 32291 -16861
rect 32294 -16895 32302 -16853
rect 30143 -16959 30626 -16925
rect 31477 -16949 31519 -16915
rect 31549 -16949 31591 -16915
rect 31863 -16956 31905 -16922
rect 31908 -16956 31916 -16911
rect 32008 -16922 32016 -16911
rect 32436 -16913 32449 -16845
rect 32477 -16879 32483 -16811
rect 32522 -16843 32528 -16775
rect 32556 -16809 32562 -16743
rect 32566 -16793 32608 -16759
rect 32769 -16838 32811 -16804
rect 32536 -16861 32544 -16853
rect 32547 -16895 32589 -16861
rect 32769 -16906 32811 -16872
rect 32019 -16956 32061 -16922
rect 30143 -16985 30613 -16959
rect 30147 -16993 30355 -16985
rect 30163 -17003 30339 -16993
rect 29889 -17140 30071 -17114
rect 29396 -17174 29438 -17140
rect 29492 -17174 29534 -17140
rect 29588 -17174 29630 -17140
rect 29684 -17174 29726 -17140
rect 29780 -17174 29822 -17140
rect 29876 -17174 30071 -17140
rect 29889 -17200 30071 -17174
rect 30089 -17174 30197 -17050
rect 30348 -17062 30355 -17051
rect 29967 -17870 30009 -17200
rect 30089 -17228 30099 -17174
rect 29774 -17936 29926 -17924
rect 29442 -17970 29926 -17936
rect 29774 -17971 29926 -17970
rect 29955 -17971 30009 -17870
rect 30101 -17971 30143 -17174
rect 30147 -17971 30154 -17174
rect 30359 -17971 30401 -17062
rect 30493 -17971 30535 -16985
rect 30746 -17002 30788 -16968
rect 30842 -17002 30884 -16968
rect 30938 -17002 30980 -16968
rect 31034 -17002 31076 -16968
rect 31130 -17002 31172 -16968
rect 31226 -17002 31268 -16968
rect 31322 -17002 31364 -16968
rect 31831 -16992 31873 -16958
rect 31903 -16992 31945 -16958
rect 32249 -16995 32291 -16961
rect 32294 -16995 32302 -16950
rect 32436 -17001 32444 -16913
rect 32818 -16922 32824 -16788
rect 32536 -16961 32544 -16950
rect 32852 -16956 32858 -16762
rect 32892 -16778 32900 -16767
rect 32888 -16809 32900 -16778
rect 33214 -16796 33256 -16762
rect 32547 -16995 32589 -16961
rect 31484 -17045 31526 -17011
rect 31580 -17045 31622 -17011
rect 31676 -17045 31718 -17011
rect 32185 -17035 32227 -17001
rect 32257 -17035 32299 -17001
rect 32329 -17035 32371 -17001
rect 32401 -17029 32444 -17001
rect 32747 -17025 32789 -16991
rect 32792 -17025 32800 -16980
rect 32888 -16992 32894 -16809
rect 32922 -16995 32928 -16812
rect 32401 -17035 32443 -17029
rect 31838 -17088 31880 -17054
rect 31934 -17088 31976 -17054
rect 32030 -17088 32072 -17054
rect 32934 -17076 32942 -16809
rect 33271 -16812 33272 -16742
rect 33305 -16819 33306 -16740
rect 33788 -16741 33801 -16673
rect 33829 -16707 33835 -16639
rect 33874 -16671 33880 -16603
rect 33908 -16637 33914 -16571
rect 33918 -16621 33960 -16587
rect 34119 -16666 34161 -16632
rect 33888 -16689 33896 -16681
rect 33899 -16723 33941 -16689
rect 34119 -16734 34161 -16700
rect 33788 -16753 33796 -16741
rect 34168 -16750 34174 -16616
rect 33563 -16819 33957 -16753
rect 34202 -16784 34208 -16590
rect 34242 -16606 34250 -16595
rect 34238 -16637 34250 -16606
rect 34564 -16624 34606 -16590
rect 32950 -16860 32992 -16826
rect 33299 -16830 33317 -16819
rect 33299 -16832 33306 -16830
rect 32950 -16928 32992 -16894
rect 33002 -16995 33008 -16860
rect 33233 -16874 33306 -16832
rect 33361 -16874 33957 -16819
rect 34097 -16853 34139 -16819
rect 34142 -16853 34150 -16808
rect 34238 -16820 34244 -16637
rect 34272 -16823 34278 -16640
rect 33233 -16877 33957 -16874
rect 33036 -16980 33042 -16892
rect 33153 -16942 33195 -16908
rect 33198 -16942 33206 -16900
rect 33034 -16991 33042 -16980
rect 33036 -17025 33042 -16991
rect 33045 -17025 33087 -16991
rect 33153 -17042 33195 -17008
rect 33198 -17042 33206 -16997
rect 33046 -17078 33088 -17044
rect 33118 -17078 33160 -17044
rect 33190 -17078 33232 -17044
rect 32192 -17131 32234 -17097
rect 32288 -17131 32330 -17097
rect 32384 -17131 32426 -17097
rect 32480 -17131 32522 -17097
rect 32576 -17131 32618 -17097
rect 33233 -17114 33385 -16877
rect 33563 -16899 33957 -16877
rect 33487 -16925 33957 -16899
rect 34284 -16904 34292 -16637
rect 34621 -16640 34622 -16570
rect 34300 -16688 34342 -16654
rect 34655 -16674 34656 -16568
rect 34849 -16577 34891 -16543
rect 34894 -16577 34902 -16532
rect 34994 -16543 35002 -16532
rect 35203 -16537 35245 -16503
rect 35248 -16537 35256 -16492
rect 35348 -16503 35356 -16492
rect 35593 -16496 35635 -16462
rect 35638 -16496 35646 -16451
rect 35359 -16537 35401 -16503
rect 35005 -16577 35047 -16543
rect 34300 -16756 34342 -16722
rect 34352 -16823 34358 -16688
rect 34914 -16691 34956 -16657
rect 34966 -16718 34972 -16641
rect 34386 -16808 34392 -16720
rect 34503 -16770 34545 -16736
rect 34548 -16770 34556 -16728
rect 34648 -16740 34656 -16729
rect 34659 -16774 34701 -16740
rect 35000 -16752 35006 -16607
rect 35203 -16620 35245 -16586
rect 35248 -16620 35256 -16575
rect 35348 -16586 35356 -16575
rect 35593 -16580 35635 -16546
rect 35638 -16580 35646 -16535
rect 35359 -16620 35401 -16586
rect 35268 -16734 35310 -16700
rect 35320 -16761 35326 -16684
rect 34384 -16819 34392 -16808
rect 34853 -16813 34895 -16779
rect 34898 -16813 34906 -16771
rect 34998 -16779 35006 -16771
rect 35009 -16813 35051 -16779
rect 35354 -16795 35360 -16650
rect 35593 -16663 35635 -16629
rect 35638 -16663 35646 -16618
rect 35715 -16679 35721 -16413
rect 35749 -16413 35791 -16379
rect 35794 -16413 35802 -16371
rect 35738 -16462 35746 -16451
rect 35749 -16462 35755 -16413
rect 35749 -16496 35791 -16462
rect 35794 -16496 35802 -16451
rect 35738 -16546 35746 -16535
rect 35749 -16546 35755 -16496
rect 35749 -16580 35791 -16546
rect 35794 -16580 35802 -16535
rect 35738 -16629 35746 -16618
rect 35749 -16629 35755 -16580
rect 35749 -16663 35791 -16629
rect 35794 -16663 35802 -16618
rect 35738 -16697 35746 -16671
rect 35749 -16713 35755 -16663
rect 35658 -16777 35700 -16743
rect 35715 -16804 35716 -16727
rect 35749 -16809 35750 -16713
rect 34386 -16853 34392 -16819
rect 34395 -16853 34437 -16819
rect 34503 -16870 34545 -16836
rect 34548 -16870 34556 -16825
rect 34648 -16832 34656 -16821
rect 34659 -16866 34701 -16832
rect 35207 -16856 35249 -16822
rect 35252 -16856 35260 -16814
rect 35352 -16822 35360 -16814
rect 35363 -16856 35405 -16822
rect 35780 -16845 35788 -16697
rect 35803 -16713 35807 -16363
rect 35837 -16679 35841 -16363
rect 35894 -16379 35902 -16371
rect 35843 -16413 35885 -16379
rect 35905 -16413 35957 -16379
rect 36615 -16422 36621 -16406
rect 36638 -16422 36646 -16414
rect 36649 -16422 36655 -16406
rect 36945 -16408 36987 -16374
rect 36990 -16408 36998 -16363
rect 35894 -16462 35902 -16451
rect 36075 -16456 36117 -16422
rect 36147 -16456 36189 -16422
rect 36219 -16456 36261 -16422
rect 36363 -16456 36405 -16422
rect 36435 -16456 36549 -16422
rect 36579 -16456 36621 -16422
rect 35905 -16496 35947 -16462
rect 35894 -16546 35902 -16535
rect 36472 -16539 36514 -16505
rect 35905 -16580 35947 -16546
rect 35894 -16629 35902 -16618
rect 35905 -16663 35947 -16629
rect 36137 -16689 36179 -16655
rect 36182 -16689 36190 -16644
rect 36259 -16706 36265 -16588
rect 36282 -16655 36290 -16644
rect 36293 -16655 36299 -16622
rect 36329 -16655 36335 -16622
rect 36293 -16689 36335 -16655
rect 36338 -16689 36346 -16644
rect 36293 -16740 36299 -16689
rect 36329 -16740 36335 -16689
rect 36363 -16706 36369 -16589
rect 36460 -16630 36461 -16589
rect 36472 -16623 36514 -16589
rect 36472 -16706 36514 -16672
rect 36615 -16706 36621 -16456
rect 36649 -16456 36691 -16422
rect 36638 -16505 36646 -16494
rect 36649 -16505 36655 -16456
rect 36945 -16491 36987 -16457
rect 36990 -16491 36998 -16446
rect 36649 -16539 36691 -16505
rect 36638 -16589 36646 -16578
rect 36649 -16589 36655 -16539
rect 36799 -16565 36907 -16499
rect 37067 -16507 37073 -16241
rect 37101 -16241 37143 -16207
rect 37146 -16241 37154 -16199
rect 37090 -16290 37098 -16279
rect 37101 -16290 37107 -16241
rect 37101 -16324 37143 -16290
rect 37146 -16324 37154 -16279
rect 37090 -16374 37098 -16363
rect 37101 -16374 37107 -16324
rect 37101 -16408 37143 -16374
rect 37146 -16408 37154 -16363
rect 37090 -16457 37098 -16446
rect 37101 -16457 37107 -16408
rect 37101 -16491 37143 -16457
rect 37146 -16491 37154 -16446
rect 37090 -16525 37098 -16499
rect 37101 -16541 37107 -16491
rect 36649 -16623 36691 -16589
rect 37010 -16605 37052 -16571
rect 36638 -16672 36646 -16661
rect 36649 -16672 36655 -16623
rect 37067 -16632 37068 -16555
rect 37101 -16637 37102 -16541
rect 36649 -16706 36691 -16672
rect 37132 -16673 37140 -16525
rect 37155 -16541 37159 -16191
rect 37189 -16507 37193 -16191
rect 37246 -16207 37254 -16199
rect 37195 -16241 37237 -16207
rect 37257 -16241 37309 -16207
rect 38172 -16231 38214 -16197
rect 38268 -16231 38274 -16197
rect 37965 -16250 37971 -16234
rect 37988 -16250 37996 -16242
rect 37999 -16250 38005 -16234
rect 37246 -16290 37254 -16279
rect 37425 -16284 37467 -16250
rect 37497 -16284 37539 -16250
rect 37569 -16284 37611 -16250
rect 37713 -16284 37755 -16250
rect 37785 -16284 37899 -16250
rect 37929 -16284 37971 -16250
rect 37257 -16324 37299 -16290
rect 37246 -16374 37254 -16363
rect 37822 -16367 37864 -16333
rect 37257 -16408 37299 -16374
rect 37246 -16457 37254 -16446
rect 37257 -16491 37299 -16457
rect 37487 -16517 37529 -16483
rect 37532 -16517 37540 -16472
rect 37609 -16534 37615 -16416
rect 37632 -16483 37640 -16472
rect 37643 -16483 37649 -16450
rect 37679 -16483 37685 -16450
rect 37643 -16517 37685 -16483
rect 37688 -16517 37696 -16472
rect 37643 -16568 37649 -16517
rect 37679 -16568 37685 -16517
rect 37713 -16534 37719 -16417
rect 37810 -16458 37811 -16417
rect 37822 -16451 37864 -16417
rect 37822 -16534 37864 -16500
rect 37965 -16534 37971 -16284
rect 37999 -16284 38041 -16250
rect 37988 -16333 37996 -16322
rect 37999 -16333 38005 -16284
rect 38238 -16293 38246 -16285
rect 38165 -16327 38235 -16293
rect 38237 -16327 38274 -16293
rect 37999 -16367 38041 -16333
rect 37988 -16417 37996 -16406
rect 37999 -16417 38005 -16367
rect 38193 -16410 38235 -16376
rect 38238 -16410 38246 -16365
rect 37999 -16451 38041 -16417
rect 37988 -16500 37996 -16489
rect 37999 -16500 38005 -16451
rect 38193 -16494 38235 -16460
rect 38238 -16494 38246 -16449
rect 37999 -16534 38041 -16500
rect 37999 -16568 38005 -16534
rect 36649 -16740 36655 -16706
rect 36945 -16723 36987 -16689
rect 36990 -16723 36998 -16681
rect 34396 -16906 34438 -16872
rect 34468 -16906 34510 -16872
rect 34540 -16906 34582 -16872
rect 34853 -16913 34895 -16879
rect 34898 -16913 34906 -16868
rect 34998 -16879 35006 -16868
rect 35009 -16913 35051 -16879
rect 35593 -16895 35635 -16861
rect 35638 -16895 35646 -16853
rect 33487 -16959 33970 -16925
rect 34821 -16949 34863 -16915
rect 34893 -16949 34935 -16915
rect 35207 -16956 35249 -16922
rect 35252 -16956 35260 -16911
rect 35352 -16922 35360 -16911
rect 35780 -16913 35793 -16845
rect 35821 -16879 35827 -16811
rect 35866 -16843 35872 -16775
rect 35900 -16809 35906 -16743
rect 35910 -16793 35952 -16759
rect 36113 -16838 36155 -16804
rect 35880 -16861 35888 -16853
rect 35891 -16895 35933 -16861
rect 36113 -16906 36155 -16872
rect 35363 -16956 35405 -16922
rect 33487 -16985 33957 -16959
rect 33491 -16993 33699 -16985
rect 33507 -17003 33683 -16993
rect 33233 -17140 33415 -17114
rect 32740 -17174 32782 -17140
rect 32836 -17174 32878 -17140
rect 32932 -17174 32974 -17140
rect 33028 -17174 33070 -17140
rect 33124 -17174 33166 -17140
rect 33220 -17174 33415 -17140
rect 33233 -17200 33415 -17174
rect 33433 -17174 33541 -17050
rect 33692 -17062 33699 -17051
rect 33311 -17870 33353 -17200
rect 33433 -17228 33443 -17174
rect 33118 -17936 33270 -17924
rect 32786 -17970 33270 -17936
rect 33118 -17971 33270 -17970
rect 33299 -17971 33353 -17870
rect 33445 -17971 33487 -17174
rect 33491 -17971 33498 -17174
rect 33703 -17971 33745 -17062
rect 33837 -17971 33879 -16985
rect 34090 -17002 34132 -16968
rect 34186 -17002 34228 -16968
rect 34282 -17002 34324 -16968
rect 34378 -17002 34420 -16968
rect 34474 -17002 34516 -16968
rect 34570 -17002 34612 -16968
rect 34666 -17002 34708 -16968
rect 35175 -16992 35217 -16958
rect 35247 -16992 35289 -16958
rect 35593 -16995 35635 -16961
rect 35638 -16995 35646 -16950
rect 35780 -17001 35788 -16913
rect 36162 -16922 36168 -16788
rect 35880 -16961 35888 -16950
rect 36196 -16956 36202 -16762
rect 36236 -16778 36244 -16767
rect 36232 -16809 36244 -16778
rect 36558 -16796 36600 -16762
rect 35891 -16995 35933 -16961
rect 34828 -17045 34870 -17011
rect 34924 -17045 34966 -17011
rect 35020 -17045 35062 -17011
rect 35529 -17035 35571 -17001
rect 35601 -17035 35643 -17001
rect 35673 -17035 35715 -17001
rect 35745 -17029 35788 -17001
rect 36091 -17025 36133 -16991
rect 36136 -17025 36144 -16980
rect 36232 -16992 36238 -16809
rect 36266 -16995 36272 -16812
rect 35745 -17035 35787 -17029
rect 35182 -17088 35224 -17054
rect 35278 -17088 35320 -17054
rect 35374 -17088 35416 -17054
rect 36278 -17076 36286 -16809
rect 36615 -16812 36616 -16742
rect 36649 -16819 36650 -16740
rect 37132 -16741 37145 -16673
rect 37173 -16707 37179 -16639
rect 37218 -16671 37224 -16603
rect 37252 -16637 37258 -16571
rect 37262 -16621 37304 -16587
rect 37463 -16666 37505 -16632
rect 37232 -16689 37240 -16681
rect 37243 -16723 37285 -16689
rect 37463 -16734 37505 -16700
rect 37132 -16753 37140 -16741
rect 37512 -16750 37518 -16616
rect 36907 -16819 37301 -16753
rect 37546 -16784 37552 -16590
rect 37586 -16606 37594 -16595
rect 37582 -16637 37594 -16606
rect 37908 -16624 37950 -16590
rect 36294 -16860 36336 -16826
rect 36643 -16830 36661 -16819
rect 36643 -16832 36650 -16830
rect 36294 -16928 36336 -16894
rect 36346 -16995 36352 -16860
rect 36577 -16874 36650 -16832
rect 36705 -16874 37301 -16819
rect 37441 -16853 37483 -16819
rect 37486 -16853 37494 -16808
rect 37582 -16820 37588 -16637
rect 37616 -16823 37622 -16640
rect 36577 -16877 37301 -16874
rect 36380 -16980 36386 -16892
rect 36497 -16942 36539 -16908
rect 36542 -16942 36550 -16900
rect 36378 -16991 36386 -16980
rect 36380 -17025 36386 -16991
rect 36389 -17025 36431 -16991
rect 36497 -17042 36539 -17008
rect 36542 -17042 36550 -16997
rect 36390 -17078 36432 -17044
rect 36462 -17078 36504 -17044
rect 36534 -17078 36576 -17044
rect 35536 -17131 35578 -17097
rect 35632 -17131 35674 -17097
rect 35728 -17131 35770 -17097
rect 35824 -17131 35866 -17097
rect 35920 -17131 35962 -17097
rect 36577 -17114 36729 -16877
rect 36907 -16899 37301 -16877
rect 36831 -16925 37301 -16899
rect 37628 -16904 37636 -16637
rect 37965 -16640 37966 -16570
rect 37644 -16688 37686 -16654
rect 37999 -16674 38000 -16568
rect 38193 -16577 38235 -16543
rect 38238 -16577 38246 -16532
rect 37644 -16756 37686 -16722
rect 37696 -16823 37702 -16688
rect 38258 -16691 38274 -16657
rect 37730 -16808 37736 -16720
rect 37847 -16770 37889 -16736
rect 37892 -16770 37900 -16728
rect 37992 -16740 38000 -16729
rect 38003 -16774 38045 -16740
rect 37728 -16819 37736 -16808
rect 38197 -16813 38239 -16779
rect 38242 -16813 38250 -16771
rect 37730 -16853 37736 -16819
rect 37739 -16853 37781 -16819
rect 37847 -16870 37889 -16836
rect 37892 -16870 37900 -16825
rect 37992 -16832 38000 -16821
rect 38003 -16866 38045 -16832
rect 37740 -16906 37782 -16872
rect 37812 -16906 37854 -16872
rect 37884 -16906 37926 -16872
rect 38197 -16913 38239 -16879
rect 38242 -16913 38250 -16868
rect 36831 -16959 37314 -16925
rect 38165 -16949 38207 -16915
rect 38237 -16949 38274 -16915
rect 36831 -16985 37301 -16959
rect 36835 -16993 37043 -16985
rect 36851 -17003 37027 -16993
rect 36577 -17140 36759 -17114
rect 36084 -17174 36126 -17140
rect 36180 -17174 36222 -17140
rect 36276 -17174 36318 -17140
rect 36372 -17174 36414 -17140
rect 36468 -17174 36510 -17140
rect 36564 -17174 36759 -17140
rect 36577 -17200 36759 -17174
rect 36777 -17174 36885 -17050
rect 37036 -17062 37043 -17051
rect 36655 -17870 36697 -17200
rect 36777 -17228 36787 -17174
rect 36462 -17936 36614 -17924
rect 36130 -17970 36614 -17936
rect 36462 -17971 36614 -17970
rect 36643 -17971 36697 -17870
rect 36789 -17971 36831 -17174
rect 36835 -17971 36842 -17174
rect 37047 -17971 37089 -17062
rect 37181 -17971 37223 -16985
rect 37434 -17002 37476 -16968
rect 37530 -17002 37572 -16968
rect 37626 -17002 37668 -16968
rect 37722 -17002 37764 -16968
rect 37818 -17002 37860 -16968
rect 37914 -17002 37956 -16968
rect 38010 -17002 38052 -16968
rect 38172 -17045 38214 -17011
rect 38268 -17045 38274 -17011
rect 6479 -18032 7146 -17971
rect 9824 -18032 10490 -17971
rect 13168 -18032 13834 -17971
rect 16513 -18032 17178 -17971
rect 19857 -18032 20522 -17971
rect 23201 -18032 23866 -17971
rect 26545 -18032 27210 -17971
rect 29774 -17982 30554 -17971
rect 33118 -17982 33898 -17971
rect 36462 -17982 37242 -17971
rect 29860 -18007 30554 -17982
rect 33204 -18007 33898 -17982
rect 36548 -18007 37242 -17982
rect 29890 -18032 30554 -18007
rect 33234 -18032 33898 -18007
rect 36578 -18032 37242 -18007
rect 6461 -18036 7146 -18032
rect 6131 -18108 6310 -18074
rect 6069 -18506 6114 -18167
rect 6115 -18506 6125 -18156
rect 6316 -18167 6326 -18156
rect 6327 -18506 6372 -18167
rect 6461 -18448 7205 -18036
rect 7214 -18118 7593 -18084
rect 7675 -18180 7689 -18118
rect 7314 -18256 7493 -18222
rect 7240 -18448 7249 -18294
rect 7252 -18448 7297 -18306
rect 7298 -18448 7308 -18295
rect 7499 -18306 7509 -18295
rect 7510 -18448 7555 -18306
rect 7558 -18448 7567 -18294
rect 7632 -18448 7641 -18220
rect 7644 -18448 7689 -18180
rect 7709 -18245 7723 -18149
rect 7805 -18183 8184 -18149
rect 7709 -18448 7754 -18245
rect 7757 -18448 7766 -18285
rect 7905 -18321 8084 -18287
rect 6461 -18506 7826 -18448
rect 5857 -18543 7826 -18506
rect 7831 -18543 7840 -18359
rect 7843 -18543 7888 -18371
rect 7889 -18543 7899 -18360
rect 8090 -18371 8100 -18360
rect 8101 -18543 8146 -18371
rect 8149 -18543 8158 -18359
rect 8223 -18543 8232 -18285
rect 8235 -18543 8280 -18245
rect 9280 -18506 9324 -18032
rect 9806 -18036 10490 -18032
rect 9476 -18108 9654 -18074
rect 9414 -18506 9458 -18167
rect 9460 -18506 9469 -18156
rect 9661 -18167 9670 -18156
rect 9672 -18506 9716 -18167
rect 9806 -18448 10549 -18036
rect 10559 -18118 10937 -18084
rect 11020 -18180 11033 -18118
rect 10659 -18256 10837 -18222
rect 10585 -18448 10593 -18294
rect 10597 -18448 10641 -18306
rect 10643 -18448 10652 -18295
rect 10844 -18306 10853 -18295
rect 10855 -18448 10899 -18306
rect 10903 -18448 10911 -18294
rect 10977 -18448 10985 -18220
rect 10989 -18448 11033 -18180
rect 11054 -18245 11067 -18149
rect 11150 -18183 11528 -18149
rect 11054 -18448 11098 -18245
rect 11102 -18448 11110 -18285
rect 11250 -18321 11428 -18287
rect 9806 -18506 11170 -18448
rect 9233 -18543 11170 -18506
rect 11176 -18543 11184 -18359
rect 11188 -18543 11232 -18371
rect 11234 -18543 11243 -18360
rect 11435 -18371 11444 -18360
rect 11446 -18543 11490 -18371
rect 11494 -18543 11502 -18359
rect 11568 -18543 11576 -18285
rect 11580 -18543 11624 -18245
rect 12624 -18506 12668 -18032
rect 13150 -18036 13834 -18032
rect 12820 -18108 12998 -18074
rect 12758 -18506 12802 -18167
rect 12804 -18506 12813 -18156
rect 13005 -18167 13014 -18156
rect 13016 -18506 13060 -18167
rect 13150 -18448 13893 -18036
rect 13903 -18118 14281 -18084
rect 14364 -18180 14377 -18118
rect 14003 -18256 14181 -18222
rect 13929 -18448 13937 -18294
rect 13941 -18448 13985 -18306
rect 13987 -18448 13996 -18295
rect 14188 -18306 14197 -18295
rect 14199 -18448 14243 -18306
rect 14247 -18448 14255 -18294
rect 14321 -18448 14329 -18220
rect 14333 -18448 14377 -18180
rect 14398 -18245 14411 -18149
rect 14494 -18183 14872 -18149
rect 14398 -18448 14442 -18245
rect 14446 -18448 14454 -18285
rect 14594 -18321 14772 -18287
rect 13150 -18506 14514 -18448
rect 12577 -18543 14514 -18506
rect 14520 -18543 14528 -18359
rect 14532 -18543 14576 -18371
rect 14578 -18543 14587 -18360
rect 14779 -18371 14788 -18360
rect 14790 -18543 14834 -18371
rect 14838 -18543 14846 -18359
rect 14912 -18543 14920 -18285
rect 14924 -18543 14968 -18245
rect 15969 -18506 16012 -18032
rect 16495 -18036 17178 -18032
rect 16165 -18108 16342 -18074
rect 16103 -18506 16146 -18167
rect 16149 -18506 16157 -18156
rect 16350 -18167 16358 -18156
rect 16361 -18506 16404 -18167
rect 16495 -18448 17237 -18036
rect 17248 -18118 17625 -18084
rect 17709 -18180 17721 -18118
rect 17348 -18256 17525 -18222
rect 17274 -18448 17281 -18294
rect 17286 -18448 17329 -18306
rect 17332 -18448 17340 -18295
rect 17533 -18306 17541 -18295
rect 17544 -18448 17587 -18306
rect 17592 -18448 17599 -18294
rect 17666 -18448 17673 -18220
rect 17678 -18448 17721 -18180
rect 17743 -18245 17755 -18149
rect 17839 -18183 18216 -18149
rect 17743 -18448 17786 -18245
rect 17791 -18448 17798 -18285
rect 17939 -18321 18116 -18287
rect 16495 -18506 17858 -18448
rect 15922 -18543 17858 -18506
rect 17865 -18543 17872 -18359
rect 17877 -18543 17920 -18371
rect 17923 -18543 17931 -18360
rect 18124 -18371 18132 -18360
rect 18135 -18543 18178 -18371
rect 18183 -18543 18190 -18359
rect 18257 -18543 18264 -18285
rect 18269 -18543 18312 -18245
rect 19313 -18506 19356 -18032
rect 19839 -18036 20522 -18032
rect 19509 -18108 19686 -18074
rect 19447 -18506 19490 -18167
rect 19493 -18506 19501 -18156
rect 19694 -18167 19702 -18156
rect 19705 -18506 19748 -18167
rect 19839 -18448 20581 -18036
rect 20592 -18118 20969 -18084
rect 21053 -18180 21065 -18118
rect 20692 -18256 20869 -18222
rect 20618 -18448 20625 -18294
rect 20630 -18448 20673 -18306
rect 20676 -18448 20684 -18295
rect 20877 -18306 20885 -18295
rect 20888 -18448 20931 -18306
rect 20936 -18448 20943 -18294
rect 21010 -18448 21017 -18220
rect 21022 -18448 21065 -18180
rect 21087 -18245 21099 -18149
rect 21183 -18183 21560 -18149
rect 21087 -18448 21130 -18245
rect 21135 -18448 21142 -18285
rect 21283 -18321 21460 -18287
rect 19839 -18506 21202 -18448
rect 19266 -18543 21202 -18506
rect 21209 -18543 21216 -18359
rect 21221 -18543 21264 -18371
rect 21267 -18543 21275 -18360
rect 21468 -18371 21476 -18360
rect 21479 -18543 21522 -18371
rect 21527 -18543 21534 -18359
rect 21601 -18543 21608 -18285
rect 21613 -18543 21656 -18245
rect 22657 -18506 22700 -18032
rect 23183 -18036 23866 -18032
rect 22853 -18108 23030 -18074
rect 22791 -18506 22834 -18167
rect 22837 -18506 22845 -18156
rect 23038 -18167 23046 -18156
rect 23049 -18506 23092 -18167
rect 23183 -18448 23925 -18036
rect 23936 -18118 24313 -18084
rect 24397 -18180 24409 -18118
rect 24036 -18256 24213 -18222
rect 23962 -18448 23969 -18294
rect 23974 -18448 24017 -18306
rect 24020 -18448 24028 -18295
rect 24221 -18306 24229 -18295
rect 24232 -18448 24275 -18306
rect 24280 -18448 24287 -18294
rect 24354 -18448 24361 -18220
rect 24366 -18448 24409 -18180
rect 24431 -18245 24443 -18149
rect 24527 -18183 24904 -18149
rect 24431 -18448 24474 -18245
rect 24479 -18448 24486 -18285
rect 24627 -18321 24804 -18287
rect 23183 -18506 24546 -18448
rect 22610 -18543 24546 -18506
rect 24553 -18543 24560 -18359
rect 24565 -18543 24608 -18371
rect 24611 -18543 24619 -18360
rect 24812 -18371 24820 -18360
rect 24823 -18543 24866 -18371
rect 24871 -18543 24878 -18359
rect 24945 -18543 24952 -18285
rect 24957 -18543 25000 -18245
rect 26001 -18506 26044 -18032
rect 26527 -18036 27210 -18032
rect 26197 -18108 26374 -18074
rect 26135 -18506 26178 -18167
rect 26181 -18506 26189 -18156
rect 26382 -18167 26390 -18156
rect 26393 -18506 26436 -18167
rect 26527 -18448 27269 -18036
rect 27280 -18118 27657 -18084
rect 27741 -18180 27753 -18118
rect 27380 -18256 27557 -18222
rect 27306 -18448 27313 -18294
rect 27318 -18448 27361 -18306
rect 27364 -18448 27372 -18295
rect 27565 -18306 27573 -18295
rect 27576 -18448 27619 -18306
rect 27624 -18448 27631 -18294
rect 27698 -18448 27705 -18220
rect 27710 -18448 27753 -18180
rect 27775 -18245 27787 -18149
rect 27871 -18183 28248 -18149
rect 27775 -18448 27818 -18245
rect 27823 -18448 27830 -18285
rect 27971 -18321 28148 -18287
rect 26527 -18506 27890 -18448
rect 25954 -18543 27890 -18506
rect 27897 -18543 27904 -18359
rect 27909 -18543 27952 -18371
rect 27955 -18543 27963 -18360
rect 28156 -18371 28164 -18360
rect 28167 -18543 28210 -18371
rect 28215 -18543 28222 -18359
rect 28289 -18543 28296 -18285
rect 28301 -18543 28344 -18245
rect 29346 -18506 29388 -18032
rect 29872 -18036 30554 -18032
rect 29542 -18108 29718 -18074
rect 29480 -18506 29522 -18167
rect 29526 -18506 29533 -18156
rect 29727 -18167 29734 -18156
rect 29738 -18506 29780 -18167
rect 29872 -18448 30613 -18036
rect 30625 -18118 31001 -18084
rect 31086 -18180 31097 -18118
rect 30725 -18256 30901 -18222
rect 30651 -18448 30657 -18294
rect 30663 -18448 30705 -18306
rect 30709 -18448 30716 -18295
rect 30910 -18306 30917 -18295
rect 30921 -18448 30963 -18306
rect 30969 -18448 30975 -18294
rect 31043 -18448 31049 -18220
rect 31055 -18448 31097 -18180
rect 31120 -18245 31131 -18149
rect 31216 -18183 31592 -18149
rect 31120 -18448 31162 -18245
rect 31168 -18448 31174 -18285
rect 31316 -18321 31492 -18287
rect 29872 -18506 31234 -18448
rect 29299 -18543 31234 -18506
rect 31242 -18543 31248 -18359
rect 31254 -18543 31296 -18371
rect 31300 -18543 31307 -18360
rect 31501 -18371 31508 -18360
rect 31512 -18543 31554 -18371
rect 31560 -18543 31566 -18359
rect 31634 -18543 31640 -18285
rect 31646 -18543 31688 -18245
rect 32690 -18506 32732 -18032
rect 33216 -18036 33898 -18032
rect 32886 -18108 33062 -18074
rect 32824 -18506 32866 -18167
rect 32870 -18506 32877 -18156
rect 33071 -18167 33078 -18156
rect 33082 -18506 33124 -18167
rect 33216 -18448 33957 -18036
rect 33969 -18118 34345 -18084
rect 34430 -18180 34441 -18118
rect 34069 -18256 34245 -18222
rect 33995 -18448 34001 -18294
rect 34007 -18448 34049 -18306
rect 34053 -18448 34060 -18295
rect 34254 -18306 34261 -18295
rect 34265 -18448 34307 -18306
rect 34313 -18448 34319 -18294
rect 34387 -18448 34393 -18220
rect 34399 -18448 34441 -18180
rect 34464 -18245 34475 -18149
rect 34560 -18183 34936 -18149
rect 34464 -18448 34506 -18245
rect 34512 -18448 34518 -18285
rect 34660 -18321 34836 -18287
rect 33216 -18506 34578 -18448
rect 32643 -18543 34578 -18506
rect 34586 -18543 34592 -18359
rect 34598 -18543 34640 -18371
rect 34644 -18543 34651 -18360
rect 34845 -18371 34852 -18360
rect 34856 -18543 34898 -18371
rect 34904 -18543 34910 -18359
rect 34978 -18543 34984 -18285
rect 34990 -18543 35032 -18245
rect 36034 -18506 36076 -18032
rect 36560 -18036 37242 -18032
rect 36230 -18108 36406 -18074
rect 36168 -18506 36210 -18167
rect 36214 -18506 36221 -18156
rect 36415 -18167 36422 -18156
rect 36426 -18506 36468 -18167
rect 36560 -18448 37301 -18036
rect 37313 -18118 37689 -18084
rect 37774 -18180 37785 -18118
rect 37413 -18256 37589 -18222
rect 37339 -18448 37345 -18294
rect 37351 -18448 37393 -18306
rect 37397 -18448 37404 -18295
rect 37598 -18306 37605 -18295
rect 37609 -18448 37651 -18306
rect 37657 -18448 37663 -18294
rect 37731 -18448 37737 -18220
rect 37743 -18448 37785 -18180
rect 37808 -18245 37819 -18149
rect 37904 -18183 38274 -18149
rect 37808 -18448 37850 -18245
rect 37856 -18448 37862 -18285
rect 38004 -18321 38180 -18287
rect 36560 -18506 37922 -18448
rect 35987 -18543 37922 -18506
rect 37930 -18543 37936 -18359
rect 37942 -18543 37984 -18371
rect 37988 -18543 37995 -18360
rect 38189 -18371 38196 -18360
rect 38200 -18543 38242 -18371
rect 38248 -18543 38254 -18359
rect 5857 -18667 8328 -18543
rect 9233 -18667 11672 -18543
rect 12577 -18667 15016 -18543
rect 15922 -18667 18360 -18543
rect 19266 -18667 21704 -18543
rect 22610 -18667 25048 -18543
rect 25954 -18667 28392 -18543
rect 29299 -18667 31736 -18543
rect 32643 -18667 35080 -18543
rect 2477 -19318 5681 -19282
rect 2477 -19763 5025 -19318
rect 5192 -19336 5681 -19318
rect 5228 -19360 5610 -19336
rect 5857 -19438 8381 -18667
rect 5888 -19622 8381 -19438
rect 9233 -19622 11725 -18667
rect 12577 -19622 15069 -18667
rect 15922 -19622 18413 -18667
rect 19266 -19622 21757 -18667
rect 22610 -19622 25101 -18667
rect 25954 -19622 28445 -18667
rect 29299 -19622 31789 -18667
rect 32643 -19622 35133 -18667
rect 35987 -19622 38274 -18543
rect 6479 -19687 8381 -19622
rect 9824 -19687 11725 -19622
rect 13168 -19687 15069 -19622
rect 16513 -19687 18413 -19622
rect 19857 -19687 21757 -19622
rect 23201 -19687 25101 -19622
rect 26545 -19687 28445 -19622
rect 29890 -19687 31789 -19622
rect 33234 -19687 35133 -19622
rect 36578 -19687 38274 -19622
rect 7070 -19747 8381 -19687
rect 10415 -19747 11725 -19687
rect 13759 -19747 15069 -19687
rect 17104 -19747 18413 -19687
rect 20448 -19747 21757 -19687
rect 23792 -19747 25101 -19687
rect 27136 -19747 28445 -19687
rect 30481 -19747 31789 -19687
rect 33825 -19747 35133 -19687
rect 37169 -19747 38274 -19687
rect 7099 -19752 8381 -19747
rect 10444 -19752 11725 -19747
rect 13788 -19752 15069 -19747
rect 17133 -19752 18413 -19747
rect 20477 -19752 21757 -19747
rect 23821 -19752 25101 -19747
rect 27165 -19752 28445 -19747
rect 30510 -19752 31789 -19747
rect 33854 -19752 35133 -19747
rect 37198 -19752 38274 -19747
rect 2477 -19781 5013 -19763
rect 7234 -19770 8381 -19752
rect 10578 -19770 11725 -19752
rect 13922 -19770 15069 -19752
rect 17266 -19770 18413 -19752
rect 20610 -19770 21757 -19752
rect 23954 -19770 25101 -19752
rect 27298 -19770 28445 -19752
rect 30642 -19770 31789 -19752
rect 33986 -19770 35133 -19752
rect 37330 -19770 38274 -19752
rect 7661 -19781 8381 -19770
rect 11006 -19781 11725 -19770
rect 14350 -19781 15069 -19770
rect 17695 -19781 18413 -19770
rect 21039 -19781 21757 -19770
rect 24383 -19781 25101 -19770
rect 27727 -19781 28445 -19770
rect 31072 -19781 31789 -19770
rect 34416 -19781 35133 -19770
rect 2477 -19813 5022 -19781
rect 2477 -19817 4984 -19813
rect 7661 -19817 8346 -19781
rect 11006 -19817 11690 -19781
rect 14350 -19817 15034 -19781
rect 17695 -19817 18378 -19781
rect 21039 -19817 21722 -19781
rect 24383 -19817 25066 -19781
rect 27727 -19817 28410 -19781
rect 31072 -19817 31754 -19781
rect 34416 -19817 35098 -19781
rect 37760 -19817 38274 -19770
rect 2477 -19825 4906 -19817
rect 4913 -19825 4947 -19817
rect 4980 -19825 4981 -19817
rect 2477 -19859 4947 -19825
rect 7855 -19835 8346 -19817
rect 11199 -19835 11690 -19817
rect 14543 -19835 15034 -19817
rect 17887 -19835 18378 -19817
rect 21231 -19835 21722 -19817
rect 24575 -19835 25066 -19817
rect 27919 -19835 28410 -19817
rect 31263 -19835 31754 -19817
rect 34607 -19835 35098 -19817
rect 37951 -19835 38274 -19817
rect 7894 -19859 8273 -19835
rect 11239 -19859 11617 -19835
rect 14583 -19859 14961 -19835
rect 17928 -19859 18305 -19835
rect 21272 -19859 21649 -19835
rect 24616 -19859 24993 -19835
rect 27960 -19859 28337 -19835
rect 31305 -19859 31681 -19835
rect 34649 -19859 35025 -19835
rect 37993 -19859 38274 -19835
rect 2477 -19871 4906 -19859
rect 4913 -19871 4947 -19859
rect 2477 -19880 4959 -19871
rect 3068 -19945 4959 -19880
rect 3659 -20005 4959 -19945
rect 3688 -20010 4959 -20005
rect 3812 -20028 4959 -20010
rect 4250 -20039 4959 -20028
rect 4250 -20075 4924 -20039
rect 4433 -20093 4924 -20075
<< error_ps >>
rect 38274 -19817 38424 -18543
rect 39331 -19622 39534 -18506
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
use idac8bit_binary_cs  x1
timestamp 1717439242
transform 1 0 0 0 1 -8000
box -79 -12195 429791 200
use idac4bit_unary_cs  x2
timestamp 1717439242
transform 1 0 1 0 1 -8000
box -90 -18645 37013 663926
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 dvdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 avss
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 iref
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 din0
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 din1
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 din2
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 din3
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 din4
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 din5
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 din6
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 din7
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 din8
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 din9
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 din10
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 din11
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 {}
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 clk
port 20 nsew
<< end >>
