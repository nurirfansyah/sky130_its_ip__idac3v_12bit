magic
tech sky130A
magscale 1 2
timestamp 1717480505
<< metal1 >>
rect 556 364992 638 672192
rect -980 -166 -780 34
rect -1004 -502 -804 -302
rect -970 -772 -770 -572
rect -984 -1098 -784 -898
rect -1038 -1432 -838 -1232
rect -1016 -1750 -816 -1550
rect -1066 -2130 -866 -1930
rect -160 -2388 -72 364992
rect 222 12 310 364992
rect 220 -2388 310 12
rect 556 -2388 644 364992
rect 936 211690 1024 672192
rect 942 -2388 1024 211690
rect 1272 -2388 1354 262592
rect 1634 -2388 1902 262592
rect 2182 -2388 2264 262592
use sky130_fd_pr__pfet_g5v0d10v5_BK8KVU  XM1
timestamp 1717439242
transform 1 0 75 0 1 181302
box -358 -183987 358 183987
use sky130_fd_pr__pfet_g5v0d10v5_AJ8KYZ  XM2
timestamp 1717439242
transform 1 0 790 0 1 334902
box -358 -337587 358 337587
use sky130_fd_pr__pfet_g5v0d10v5_GK83LR  XM3
timestamp 1717439242
transform 1 0 1505 0 1 130102
box -358 -132787 358 132787
use sky130_fd_pr__pfet_g5v0d10v5_GK83LR  XM4
timestamp 1717439242
transform 1 0 2031 0 1 130102
box -358 -132787 358 132787
<< labels >>
flabel metal1 -1066 -2130 -866 -1930 0 FreeSans 256 0 0 0 iout
port 6 nsew
flabel metal1 -1016 -1750 -816 -1550 0 FreeSans 256 0 0 0 iout_n
port 5 nsew
flabel metal1 -1038 -1432 -838 -1232 0 FreeSans 256 0 0 0 sw_bn
port 4 nsew
flabel metal1 -984 -1098 -784 -898 0 FreeSans 256 0 0 0 sw_b
port 3 nsew
flabel metal1 -970 -772 -770 -572 0 FreeSans 256 0 0 0 pcbias
port 2 nsew
flabel metal1 -1004 -502 -804 -302 0 FreeSans 256 0 0 0 pbias
port 1 nsew
flabel metal1 -980 -166 -780 34 0 FreeSans 256 0 0 0 avdd
port 0 nsew
<< end >>
