magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< error_p >>
rect 19685 -17967 19723 -17952
rect 22151 -18010 22189 -17985
rect 24617 -18053 24655 -18028
rect 27083 -18096 27121 -18071
rect 29549 -18139 29587 -18114
rect 32015 -18182 32053 -18157
rect 34481 -18225 34519 -18200
<< error_s >>
rect 3985 663814 4367 663848
rect 3889 356809 3937 663752
rect 4085 663676 4267 663710
rect 4069 663617 4071 663628
rect 4270 663617 4283 663628
rect 4023 661241 4071 663617
rect 4281 661241 4329 663617
rect 4085 661148 4267 661182
rect 4085 661040 4267 661074
rect 4069 660981 4071 660992
rect 4270 660981 4283 660992
rect 4023 658605 4071 660981
rect 4281 658605 4329 660981
rect 4085 658512 4267 658546
rect 4085 658404 4267 658438
rect 4069 658345 4071 658356
rect 4270 658345 4283 658356
rect 4023 655969 4071 658345
rect 4281 655969 4329 658345
rect 4085 655876 4267 655910
rect 4085 655768 4267 655802
rect 4069 655709 4071 655720
rect 4270 655709 4283 655720
rect 4023 653333 4071 655709
rect 4281 653333 4329 655709
rect 4085 653240 4267 653274
rect 4085 653132 4267 653166
rect 4069 653073 4071 653084
rect 4270 653073 4283 653084
rect 4023 650697 4071 653073
rect 4281 650697 4329 653073
rect 4085 650604 4267 650638
rect 4085 650496 4267 650530
rect 4069 650437 4071 650448
rect 4270 650437 4283 650448
rect 4023 648061 4071 650437
rect 4281 648061 4329 650437
rect 4085 647968 4267 648002
rect 4085 647860 4267 647894
rect 4069 647801 4071 647812
rect 4270 647801 4283 647812
rect 4023 645425 4071 647801
rect 4281 645425 4329 647801
rect 4085 645332 4267 645366
rect 4085 645224 4267 645258
rect 4069 645165 4071 645176
rect 4270 645165 4283 645176
rect 4023 642789 4071 645165
rect 4281 642789 4329 645165
rect 4085 642696 4267 642730
rect 4085 642588 4267 642622
rect 4069 642529 4071 642540
rect 4270 642529 4283 642540
rect 4023 640153 4071 642529
rect 4281 640153 4329 642529
rect 4085 640060 4267 640094
rect 4085 639952 4267 639986
rect 4069 639893 4071 639904
rect 4270 639893 4283 639904
rect 4023 637517 4071 639893
rect 4281 637517 4329 639893
rect 4085 637424 4267 637458
rect 4085 637316 4267 637350
rect 4069 637257 4071 637268
rect 4270 637257 4283 637268
rect 4023 634881 4071 637257
rect 4281 634881 4329 637257
rect 4085 634788 4267 634822
rect 4085 634680 4267 634714
rect 4069 634621 4071 634632
rect 4270 634621 4283 634632
rect 4023 632245 4071 634621
rect 4281 632245 4329 634621
rect 4085 632152 4267 632186
rect 4085 632044 4267 632078
rect 4069 631985 4071 631996
rect 4270 631985 4283 631996
rect 4023 629609 4071 631985
rect 4281 629609 4329 631985
rect 4085 629516 4267 629550
rect 4085 629408 4267 629442
rect 4069 629349 4071 629360
rect 4270 629349 4283 629360
rect 4023 626973 4071 629349
rect 4281 626973 4329 629349
rect 4085 626880 4267 626914
rect 4085 626772 4267 626806
rect 4069 626713 4071 626724
rect 4270 626713 4283 626724
rect 4023 624337 4071 626713
rect 4281 624337 4329 626713
rect 4085 624244 4267 624278
rect 4085 624136 4267 624170
rect 4069 624077 4071 624088
rect 4270 624077 4283 624088
rect 4023 621701 4071 624077
rect 4281 621701 4329 624077
rect 4085 621608 4267 621642
rect 4085 621500 4267 621534
rect 4069 621441 4071 621452
rect 4270 621441 4283 621452
rect 4023 619065 4071 621441
rect 4281 619065 4329 621441
rect 4085 618972 4267 619006
rect 4085 618864 4267 618898
rect 4069 618805 4071 618816
rect 4270 618805 4283 618816
rect 4023 616429 4071 618805
rect 4281 616429 4329 618805
rect 4085 616336 4267 616370
rect 4085 616228 4267 616262
rect 4069 616169 4071 616180
rect 4270 616169 4283 616180
rect 4023 613793 4071 616169
rect 4281 613793 4329 616169
rect 4085 613700 4267 613734
rect 4085 613592 4267 613626
rect 4069 613533 4071 613544
rect 4270 613533 4283 613544
rect 4023 611157 4071 613533
rect 4281 611157 4329 613533
rect 4085 611064 4267 611098
rect 4085 610956 4267 610990
rect 4069 610897 4071 610908
rect 4270 610897 4283 610908
rect 4023 608521 4071 610897
rect 4281 608521 4329 610897
rect 4085 608428 4267 608462
rect 4085 608320 4267 608354
rect 4069 608261 4071 608272
rect 4270 608261 4283 608272
rect 4023 605885 4071 608261
rect 4281 605885 4329 608261
rect 4085 605792 4267 605826
rect 4085 605684 4267 605718
rect 4069 605625 4071 605636
rect 4270 605625 4283 605636
rect 4023 603249 4071 605625
rect 4281 603249 4329 605625
rect 4085 603156 4267 603190
rect 4085 603048 4267 603082
rect 4069 602989 4071 603000
rect 4270 602989 4283 603000
rect 4023 600613 4071 602989
rect 4281 600613 4329 602989
rect 4085 600520 4267 600554
rect 4085 600412 4267 600446
rect 4069 600353 4071 600364
rect 4270 600353 4283 600364
rect 4023 597977 4071 600353
rect 4281 597977 4329 600353
rect 4085 597884 4267 597918
rect 4085 597776 4267 597810
rect 4069 597717 4071 597728
rect 4270 597717 4283 597728
rect 4023 595341 4071 597717
rect 4281 595341 4329 597717
rect 4085 595248 4267 595282
rect 4085 595140 4267 595174
rect 4069 595081 4071 595092
rect 4270 595081 4283 595092
rect 4023 592705 4071 595081
rect 4281 592705 4329 595081
rect 4085 592612 4267 592646
rect 4085 592504 4267 592538
rect 4069 592445 4071 592456
rect 4270 592445 4283 592456
rect 4023 590069 4071 592445
rect 4281 590069 4329 592445
rect 4085 589976 4267 590010
rect 4085 589868 4267 589902
rect 4069 589809 4071 589820
rect 4270 589809 4283 589820
rect 4023 587433 4071 589809
rect 4281 587433 4329 589809
rect 4085 587340 4267 587374
rect 4085 587232 4267 587266
rect 4069 587173 4071 587184
rect 4270 587173 4283 587184
rect 4023 584797 4071 587173
rect 4281 584797 4329 587173
rect 4085 584704 4267 584738
rect 4085 584596 4267 584630
rect 4069 584537 4071 584548
rect 4270 584537 4283 584548
rect 4023 582161 4071 584537
rect 4281 582161 4329 584537
rect 4085 582068 4267 582102
rect 4085 581960 4267 581994
rect 4069 581901 4071 581912
rect 4270 581901 4283 581912
rect 4023 579525 4071 581901
rect 4281 579525 4329 581901
rect 4085 579432 4267 579466
rect 4085 579324 4267 579358
rect 4069 579265 4071 579276
rect 4270 579265 4283 579276
rect 4023 576889 4071 579265
rect 4281 576889 4329 579265
rect 4085 576796 4267 576830
rect 4085 576688 4267 576722
rect 4069 576629 4071 576640
rect 4270 576629 4283 576640
rect 4023 574253 4071 576629
rect 4281 574253 4329 576629
rect 4085 574160 4267 574194
rect 4085 574052 4267 574086
rect 4069 573993 4071 574004
rect 4270 573993 4283 574004
rect 4023 571617 4071 573993
rect 4281 571617 4329 573993
rect 4085 571524 4267 571558
rect 4085 571416 4267 571450
rect 4069 571357 4071 571368
rect 4270 571357 4283 571368
rect 4023 568981 4071 571357
rect 4281 568981 4329 571357
rect 4085 568888 4267 568922
rect 4085 568780 4267 568814
rect 4069 568721 4071 568732
rect 4270 568721 4283 568732
rect 4023 566345 4071 568721
rect 4281 566345 4329 568721
rect 4085 566252 4267 566286
rect 4085 566144 4267 566178
rect 4069 566085 4071 566096
rect 4270 566085 4283 566096
rect 4023 563709 4071 566085
rect 4281 563709 4329 566085
rect 4085 563616 4267 563650
rect 4085 563508 4267 563542
rect 4069 563449 4071 563460
rect 4270 563449 4283 563460
rect 4023 561073 4071 563449
rect 4281 561073 4329 563449
rect 4085 560980 4267 561014
rect 4085 560872 4267 560906
rect 4069 560813 4071 560824
rect 4270 560813 4283 560824
rect 4023 558437 4071 560813
rect 4281 558437 4329 560813
rect 4085 558344 4267 558378
rect 4085 558236 4267 558270
rect 4069 558177 4071 558188
rect 4270 558177 4283 558188
rect 4023 555801 4071 558177
rect 4281 555801 4329 558177
rect 4085 555708 4267 555742
rect 4085 555600 4267 555634
rect 4069 555541 4071 555552
rect 4270 555541 4283 555552
rect 4023 553165 4071 555541
rect 4281 553165 4329 555541
rect 4085 553072 4267 553106
rect 4085 552964 4267 552998
rect 4069 552905 4071 552916
rect 4270 552905 4283 552916
rect 4023 550529 4071 552905
rect 4281 550529 4329 552905
rect 4085 550436 4267 550470
rect 4085 550328 4267 550362
rect 4069 550269 4071 550280
rect 4270 550269 4283 550280
rect 4023 547893 4071 550269
rect 4281 547893 4329 550269
rect 4085 547800 4267 547834
rect 4085 547692 4267 547726
rect 4069 547633 4071 547644
rect 4270 547633 4283 547644
rect 4023 545257 4071 547633
rect 4281 545257 4329 547633
rect 4085 545164 4267 545198
rect 4085 545056 4267 545090
rect 4069 544997 4071 545008
rect 4270 544997 4283 545008
rect 4023 542621 4071 544997
rect 4281 542621 4329 544997
rect 4085 542528 4267 542562
rect 4085 542420 4267 542454
rect 4069 542361 4071 542372
rect 4270 542361 4283 542372
rect 4023 539985 4071 542361
rect 4281 539985 4329 542361
rect 4085 539892 4267 539926
rect 4085 539784 4267 539818
rect 4069 539725 4071 539736
rect 4270 539725 4283 539736
rect 4023 537349 4071 539725
rect 4281 537349 4329 539725
rect 4085 537256 4267 537290
rect 4085 537148 4267 537182
rect 4069 537089 4071 537100
rect 4270 537089 4283 537100
rect 4023 534713 4071 537089
rect 4281 534713 4329 537089
rect 4085 534620 4267 534654
rect 4085 534512 4267 534546
rect 4069 534453 4071 534464
rect 4270 534453 4283 534464
rect 4023 532077 4071 534453
rect 4281 532077 4329 534453
rect 4085 531984 4267 532018
rect 4085 531876 4267 531910
rect 4069 531817 4071 531828
rect 4270 531817 4283 531828
rect 4023 529441 4071 531817
rect 4281 529441 4329 531817
rect 4085 529348 4267 529382
rect 4085 529240 4267 529274
rect 4069 529181 4071 529192
rect 4270 529181 4283 529192
rect 4023 526805 4071 529181
rect 4281 526805 4329 529181
rect 4085 526712 4267 526746
rect 4085 526604 4267 526638
rect 4069 526545 4071 526556
rect 4270 526545 4283 526556
rect 4023 524169 4071 526545
rect 4281 524169 4329 526545
rect 4085 524076 4267 524110
rect 4085 523968 4267 524002
rect 4069 523909 4071 523920
rect 4270 523909 4283 523920
rect 4023 521533 4071 523909
rect 4281 521533 4329 523909
rect 4085 521440 4267 521474
rect 4085 521332 4267 521366
rect 4069 521273 4071 521284
rect 4270 521273 4283 521284
rect 4023 518897 4071 521273
rect 4281 518897 4329 521273
rect 4085 518804 4267 518838
rect 4085 518696 4267 518730
rect 4069 518637 4071 518648
rect 4270 518637 4283 518648
rect 4023 516261 4071 518637
rect 4281 516261 4329 518637
rect 4085 516168 4267 516202
rect 4085 516060 4267 516094
rect 4069 516001 4071 516012
rect 4270 516001 4283 516012
rect 4023 513625 4071 516001
rect 4281 513625 4329 516001
rect 4085 513532 4267 513566
rect 4085 513424 4267 513458
rect 4069 513365 4071 513376
rect 4270 513365 4283 513376
rect 4023 510989 4071 513365
rect 4281 510989 4329 513365
rect 4085 510896 4267 510930
rect 4085 510788 4267 510822
rect 4069 510729 4071 510740
rect 4270 510729 4283 510740
rect 4023 508353 4071 510729
rect 4281 508353 4329 510729
rect 4085 508260 4267 508294
rect 4085 508152 4267 508186
rect 4069 508093 4071 508104
rect 4270 508093 4283 508104
rect 4023 505717 4071 508093
rect 4281 505717 4329 508093
rect 4085 505624 4267 505658
rect 4085 505516 4267 505550
rect 4069 505457 4071 505468
rect 4270 505457 4283 505468
rect 4023 503081 4071 505457
rect 4281 503081 4329 505457
rect 4085 502988 4267 503022
rect 4085 502880 4267 502914
rect 4069 502821 4071 502832
rect 4270 502821 4283 502832
rect 4023 500445 4071 502821
rect 4281 500445 4329 502821
rect 4085 500352 4267 500386
rect 4085 500244 4267 500278
rect 4069 500185 4071 500196
rect 4270 500185 4283 500196
rect 4023 497809 4071 500185
rect 4281 497809 4329 500185
rect 4085 497716 4267 497750
rect 4085 497608 4267 497642
rect 4069 497549 4071 497560
rect 4270 497549 4283 497560
rect 4023 495173 4071 497549
rect 4281 495173 4329 497549
rect 4085 495080 4267 495114
rect 4085 494972 4267 495006
rect 4069 494913 4071 494924
rect 4270 494913 4283 494924
rect 4023 492537 4071 494913
rect 4281 492537 4329 494913
rect 4085 492444 4267 492478
rect 4085 492336 4267 492370
rect 4069 492277 4071 492288
rect 4270 492277 4283 492288
rect 4023 489901 4071 492277
rect 4281 489901 4329 492277
rect 4085 489808 4267 489842
rect 4085 489700 4267 489734
rect 4069 489641 4071 489652
rect 4270 489641 4283 489652
rect 4023 487265 4071 489641
rect 4281 487265 4329 489641
rect 4085 487172 4267 487206
rect 4085 487064 4267 487098
rect 4069 487005 4071 487016
rect 4270 487005 4283 487016
rect 4023 484629 4071 487005
rect 4281 484629 4329 487005
rect 4085 484536 4267 484570
rect 4085 484428 4267 484462
rect 4069 484369 4071 484380
rect 4270 484369 4283 484380
rect 4023 481993 4071 484369
rect 4281 481993 4329 484369
rect 4085 481900 4267 481934
rect 4085 481792 4267 481826
rect 4069 481733 4071 481744
rect 4270 481733 4283 481744
rect 4023 479357 4071 481733
rect 4281 479357 4329 481733
rect 4085 479264 4267 479298
rect 4085 479156 4267 479190
rect 4069 479097 4071 479108
rect 4270 479097 4283 479108
rect 4023 476721 4071 479097
rect 4281 476721 4329 479097
rect 4085 476628 4267 476662
rect 4085 476520 4267 476554
rect 4069 476461 4071 476472
rect 4270 476461 4283 476472
rect 4023 474085 4071 476461
rect 4281 474085 4329 476461
rect 4085 473992 4267 474026
rect 4085 473884 4267 473918
rect 4069 473825 4071 473836
rect 4270 473825 4283 473836
rect 4023 471449 4071 473825
rect 4281 471449 4329 473825
rect 4085 471356 4267 471390
rect 4085 471248 4267 471282
rect 4069 471189 4071 471200
rect 4270 471189 4283 471200
rect 4023 468813 4071 471189
rect 4281 468813 4329 471189
rect 4085 468720 4267 468754
rect 4085 468612 4267 468646
rect 4069 468553 4071 468564
rect 4270 468553 4283 468564
rect 4023 466177 4071 468553
rect 4281 466177 4329 468553
rect 4085 466084 4267 466118
rect 4085 465976 4267 466010
rect 4069 465917 4071 465928
rect 4270 465917 4283 465928
rect 4023 463541 4071 465917
rect 4281 463541 4329 465917
rect 4085 463448 4267 463482
rect 4085 463340 4267 463374
rect 4069 463281 4071 463292
rect 4270 463281 4283 463292
rect 4023 460905 4071 463281
rect 4281 460905 4329 463281
rect 4085 460812 4267 460846
rect 4085 460704 4267 460738
rect 4069 460645 4071 460656
rect 4270 460645 4283 460656
rect 4023 458269 4071 460645
rect 4281 458269 4329 460645
rect 4085 458176 4267 458210
rect 4085 458068 4267 458102
rect 4069 458009 4071 458020
rect 4270 458009 4283 458020
rect 4023 455633 4071 458009
rect 4281 455633 4329 458009
rect 4085 455540 4267 455574
rect 4085 455432 4267 455466
rect 4069 455373 4071 455384
rect 4270 455373 4283 455384
rect 4023 452997 4071 455373
rect 4281 452997 4329 455373
rect 4085 452904 4267 452938
rect 4085 452796 4267 452830
rect 4069 452737 4071 452748
rect 4270 452737 4283 452748
rect 4023 450361 4071 452737
rect 4281 450361 4329 452737
rect 4085 450268 4267 450302
rect 4085 450160 4267 450194
rect 4069 450101 4071 450112
rect 4270 450101 4283 450112
rect 4023 447725 4071 450101
rect 4281 447725 4329 450101
rect 4085 447632 4267 447666
rect 4085 447524 4267 447558
rect 4069 447465 4071 447476
rect 4270 447465 4283 447476
rect 4023 445089 4071 447465
rect 4281 445089 4329 447465
rect 4085 444996 4267 445030
rect 4085 444888 4267 444922
rect 4069 444829 4071 444840
rect 4270 444829 4283 444840
rect 4023 442453 4071 444829
rect 4281 442453 4329 444829
rect 4085 442360 4267 442394
rect 4085 442252 4267 442286
rect 4069 442193 4071 442204
rect 4270 442193 4283 442204
rect 4023 439817 4071 442193
rect 4281 439817 4329 442193
rect 4085 439724 4267 439758
rect 4085 439616 4267 439650
rect 4069 439557 4071 439568
rect 4270 439557 4283 439568
rect 4023 437181 4071 439557
rect 4281 437181 4329 439557
rect 4085 437088 4267 437122
rect 4085 436980 4267 437014
rect 4069 436921 4071 436932
rect 4270 436921 4283 436932
rect 4023 434545 4071 436921
rect 4281 434545 4329 436921
rect 4085 434452 4267 434486
rect 4085 434344 4267 434378
rect 4069 434285 4071 434296
rect 4270 434285 4283 434296
rect 4023 431909 4071 434285
rect 4281 431909 4329 434285
rect 4085 431816 4267 431850
rect 4085 431708 4267 431742
rect 4069 431649 4071 431660
rect 4270 431649 4283 431660
rect 4023 429273 4071 431649
rect 4281 429273 4329 431649
rect 4085 429180 4267 429214
rect 4085 429072 4267 429106
rect 4069 429013 4071 429024
rect 4270 429013 4283 429024
rect 4023 426637 4071 429013
rect 4281 426637 4329 429013
rect 4085 426544 4267 426578
rect 4085 426436 4267 426470
rect 4069 426377 4071 426388
rect 4270 426377 4283 426388
rect 4023 424001 4071 426377
rect 4281 424001 4329 426377
rect 4085 423908 4267 423942
rect 4085 423800 4267 423834
rect 4069 423741 4071 423752
rect 4270 423741 4283 423752
rect 4023 421365 4071 423741
rect 4281 421365 4329 423741
rect 4085 421272 4267 421306
rect 4085 421164 4267 421198
rect 4069 421105 4071 421116
rect 4270 421105 4283 421116
rect 4023 418729 4071 421105
rect 4281 418729 4329 421105
rect 4085 418636 4267 418670
rect 4085 418528 4267 418562
rect 4069 418469 4071 418480
rect 4270 418469 4283 418480
rect 4023 416093 4071 418469
rect 4281 416093 4329 418469
rect 4085 416000 4267 416034
rect 4085 415892 4267 415926
rect 4069 415833 4071 415844
rect 4270 415833 4283 415844
rect 4023 413457 4071 415833
rect 4281 413457 4329 415833
rect 4085 413364 4267 413398
rect 4085 413256 4267 413290
rect 4069 413197 4071 413208
rect 4270 413197 4283 413208
rect 4023 410821 4071 413197
rect 4281 410821 4329 413197
rect 4085 410728 4267 410762
rect 4085 410620 4267 410654
rect 4069 410561 4071 410572
rect 4270 410561 4283 410572
rect 4023 408185 4071 410561
rect 4281 408185 4329 410561
rect 4085 408092 4267 408126
rect 4085 407984 4267 408018
rect 4069 407925 4071 407936
rect 4270 407925 4283 407936
rect 4023 405549 4071 407925
rect 4281 405549 4329 407925
rect 4085 405456 4267 405490
rect 4085 405348 4267 405382
rect 4069 405289 4071 405300
rect 4270 405289 4283 405300
rect 4023 402913 4071 405289
rect 4281 402913 4329 405289
rect 4085 402820 4267 402854
rect 4085 402712 4267 402746
rect 4069 402653 4071 402664
rect 4270 402653 4283 402664
rect 4023 400277 4071 402653
rect 4281 400277 4329 402653
rect 4085 400184 4267 400218
rect 4085 400076 4267 400110
rect 4069 400017 4071 400028
rect 4270 400017 4283 400028
rect 4023 397641 4071 400017
rect 4281 397641 4329 400017
rect 4085 397548 4267 397582
rect 4085 397440 4267 397474
rect 4069 397381 4071 397392
rect 4270 397381 4283 397392
rect 4023 395005 4071 397381
rect 4281 395005 4329 397381
rect 4085 394912 4267 394946
rect 4085 394804 4267 394838
rect 4069 394745 4071 394756
rect 4270 394745 4283 394756
rect 4023 392369 4071 394745
rect 4281 392369 4329 394745
rect 4085 392276 4267 392310
rect 4085 392168 4267 392202
rect 4069 392109 4071 392120
rect 4270 392109 4283 392120
rect 4023 389733 4071 392109
rect 4281 389733 4329 392109
rect 4085 389640 4267 389674
rect 4085 389532 4267 389566
rect 4069 389473 4071 389484
rect 4270 389473 4283 389484
rect 4023 387097 4071 389473
rect 4281 387097 4329 389473
rect 4085 387004 4267 387038
rect 4085 386896 4267 386930
rect 4069 386837 4071 386848
rect 4270 386837 4283 386848
rect 4023 384461 4071 386837
rect 4281 384461 4329 386837
rect 4085 384368 4267 384402
rect 4085 384260 4267 384294
rect 4069 384201 4071 384212
rect 4270 384201 4283 384212
rect 4023 381825 4071 384201
rect 4281 381825 4329 384201
rect 4085 381732 4267 381766
rect 4085 381624 4267 381658
rect 4069 381565 4071 381576
rect 4270 381565 4283 381576
rect 4023 379189 4071 381565
rect 4281 379189 4329 381565
rect 4085 379096 4267 379130
rect 4085 378988 4267 379022
rect 4069 378929 4071 378940
rect 4270 378929 4283 378940
rect 4023 376553 4071 378929
rect 4281 376553 4329 378929
rect 4085 376460 4267 376494
rect 4085 376352 4267 376386
rect 4069 376293 4071 376304
rect 4270 376293 4283 376304
rect 4023 373917 4071 376293
rect 4281 373917 4329 376293
rect 4085 373824 4267 373858
rect 4085 373716 4267 373750
rect 4069 373657 4071 373668
rect 4270 373657 4283 373668
rect 4023 371281 4071 373657
rect 4281 371281 4329 373657
rect 4085 371188 4267 371222
rect 4085 371080 4267 371114
rect 4069 371021 4071 371032
rect 4270 371021 4283 371032
rect 4023 368645 4071 371021
rect 4281 368645 4329 371021
rect 4085 368552 4267 368586
rect 4085 368444 4267 368478
rect 4069 368385 4071 368396
rect 4270 368385 4283 368396
rect 4023 366009 4071 368385
rect 4281 366009 4329 368385
rect 4085 365916 4267 365950
rect 4085 365808 4267 365842
rect 4069 365749 4071 365760
rect 4270 365749 4283 365760
rect 4023 363373 4071 365749
rect 4281 363373 4329 365749
rect 4085 363280 4267 363314
rect 4085 363172 4267 363206
rect 4069 363113 4071 363124
rect 4270 363113 4283 363124
rect 4023 360737 4071 363113
rect 4281 360737 4329 363113
rect 4085 360644 4267 360678
rect 4085 360536 4267 360570
rect 4069 360477 4071 360488
rect 4270 360477 4283 360488
rect 4023 358101 4071 360477
rect 4281 358101 4329 360477
rect 4085 358008 4267 358042
rect 4085 357900 4267 357934
rect 4069 357841 4071 357852
rect 4270 357841 4283 357852
rect 3364 356709 3746 356743
rect 3823 356647 3854 356755
rect 3268 198583 3316 356647
rect 3464 356571 3646 356605
rect 3448 356512 3450 356523
rect 3649 356512 3662 356523
rect 3402 355336 3450 356512
rect 3660 355336 3708 356512
rect 3464 355243 3646 355277
rect 3464 355135 3646 355169
rect 3448 355076 3450 355087
rect 3649 355076 3662 355087
rect 3402 353900 3450 355076
rect 3660 353900 3708 355076
rect 3464 353807 3646 353841
rect 3464 353699 3646 353733
rect 3448 353640 3450 353651
rect 3649 353640 3662 353651
rect 3402 352464 3450 353640
rect 3660 352464 3708 353640
rect 3464 352371 3646 352405
rect 3464 352263 3646 352297
rect 3448 352204 3450 352215
rect 3649 352204 3662 352215
rect 3402 351028 3450 352204
rect 3660 351028 3708 352204
rect 3794 352118 3854 356647
rect 3877 352118 3937 356809
rect 4023 355465 4071 357841
rect 4281 355465 4329 357841
rect 4085 355372 4267 355406
rect 4085 355264 4267 355298
rect 4069 355205 4071 355216
rect 4270 355205 4283 355216
rect 4023 352829 4071 355205
rect 4281 352829 4329 355205
rect 4085 352736 4267 352770
rect 4085 352628 4267 352662
rect 4069 352569 4071 352580
rect 4270 352569 4283 352580
rect 4023 352118 4071 352569
rect 4281 352118 4329 352569
rect 4415 352118 4463 663752
rect 3794 352053 4480 352118
rect 3464 350935 3646 350969
rect 3464 350827 3646 350861
rect 3448 350768 3450 350779
rect 3649 350768 3662 350779
rect 3402 349592 3450 350768
rect 3660 349592 3708 350768
rect 3464 349499 3646 349533
rect 3464 349391 3646 349425
rect 3448 349332 3450 349343
rect 3649 349332 3662 349343
rect 3402 348156 3450 349332
rect 3660 348156 3708 349332
rect 3464 348063 3646 348097
rect 3464 347955 3646 347989
rect 3448 347896 3450 347907
rect 3649 347896 3662 347907
rect 3402 346720 3450 347896
rect 3660 346720 3708 347896
rect 3464 346627 3646 346661
rect 3464 346519 3646 346553
rect 3448 346460 3450 346471
rect 3649 346460 3662 346471
rect 3402 345284 3450 346460
rect 3660 345284 3708 346460
rect 3464 345191 3646 345225
rect 3464 345083 3646 345117
rect 3448 345024 3450 345035
rect 3649 345024 3662 345035
rect 3402 343848 3450 345024
rect 3660 343848 3708 345024
rect 3464 343755 3646 343789
rect 3464 343647 3646 343681
rect 3448 343588 3450 343599
rect 3649 343588 3662 343599
rect 3402 342412 3450 343588
rect 3660 342412 3708 343588
rect 3464 342319 3646 342353
rect 3464 342211 3646 342245
rect 3448 342152 3450 342163
rect 3649 342152 3662 342163
rect 3402 340976 3450 342152
rect 3660 340976 3708 342152
rect 3464 340883 3646 340917
rect 3464 340775 3646 340809
rect 3448 340716 3450 340727
rect 3649 340716 3662 340727
rect 3402 339540 3450 340716
rect 3660 339540 3708 340716
rect 3464 339447 3646 339481
rect 3464 339339 3646 339373
rect 3448 339280 3450 339291
rect 3649 339280 3662 339291
rect 3402 338104 3450 339280
rect 3660 338104 3708 339280
rect 3464 338011 3646 338045
rect 3464 337903 3646 337937
rect 3448 337844 3450 337855
rect 3649 337844 3662 337855
rect 3402 336668 3450 337844
rect 3660 336668 3708 337844
rect 3464 336575 3646 336609
rect 3464 336467 3646 336501
rect 3448 336408 3450 336419
rect 3649 336408 3662 336419
rect 3402 335232 3450 336408
rect 3660 335232 3708 336408
rect 3464 335139 3646 335173
rect 3464 335031 3646 335065
rect 3448 334972 3450 334983
rect 3649 334972 3662 334983
rect 3402 333796 3450 334972
rect 3660 333796 3708 334972
rect 3464 333703 3646 333737
rect 3464 333595 3646 333629
rect 3448 333536 3450 333547
rect 3649 333536 3662 333547
rect 3402 332360 3450 333536
rect 3660 332360 3708 333536
rect 3464 332267 3646 332301
rect 3464 332159 3646 332193
rect 3448 332100 3450 332111
rect 3649 332100 3662 332111
rect 3402 330924 3450 332100
rect 3660 330924 3708 332100
rect 3464 330831 3646 330865
rect 3464 330723 3646 330757
rect 3448 330664 3450 330675
rect 3649 330664 3662 330675
rect 3402 329488 3450 330664
rect 3660 329488 3708 330664
rect 3464 329395 3646 329429
rect 3464 329287 3646 329321
rect 3448 329228 3450 329239
rect 3649 329228 3662 329239
rect 3402 328052 3450 329228
rect 3660 328052 3708 329228
rect 3464 327959 3646 327993
rect 3464 327851 3646 327885
rect 3448 327792 3450 327803
rect 3649 327792 3662 327803
rect 3402 326616 3450 327792
rect 3660 326616 3708 327792
rect 3464 326523 3646 326557
rect 3464 326415 3646 326449
rect 3448 326356 3450 326367
rect 3649 326356 3662 326367
rect 3402 325180 3450 326356
rect 3660 325180 3708 326356
rect 3464 325087 3646 325121
rect 3464 324979 3646 325013
rect 3448 324920 3450 324931
rect 3649 324920 3662 324931
rect 3402 323744 3450 324920
rect 3660 323744 3708 324920
rect 3464 323651 3646 323685
rect 3464 323543 3646 323577
rect 3448 323484 3450 323495
rect 3649 323484 3662 323495
rect 3402 322308 3450 323484
rect 3660 322308 3708 323484
rect 3464 322215 3646 322249
rect 3464 322107 3646 322141
rect 3448 322048 3450 322059
rect 3649 322048 3662 322059
rect 3402 320872 3450 322048
rect 3660 320872 3708 322048
rect 3464 320779 3646 320813
rect 3464 320671 3646 320705
rect 3448 320612 3450 320623
rect 3649 320612 3662 320623
rect 3402 319436 3450 320612
rect 3660 319436 3708 320612
rect 3464 319343 3646 319377
rect 3464 319235 3646 319269
rect 3448 319176 3450 319187
rect 3649 319176 3662 319187
rect 3402 318000 3450 319176
rect 3660 318000 3708 319176
rect 3464 317907 3646 317941
rect 3464 317799 3646 317833
rect 3448 317740 3450 317751
rect 3649 317740 3662 317751
rect 3402 316564 3450 317740
rect 3660 316564 3708 317740
rect 3464 316471 3646 316505
rect 3464 316363 3646 316397
rect 3448 316304 3450 316315
rect 3649 316304 3662 316315
rect 3402 315128 3450 316304
rect 3660 315128 3708 316304
rect 3464 315035 3646 315069
rect 3464 314927 3646 314961
rect 3448 314868 3450 314879
rect 3649 314868 3662 314879
rect 3402 313692 3450 314868
rect 3660 313692 3708 314868
rect 3464 313599 3646 313633
rect 3464 313491 3646 313525
rect 3448 313432 3450 313443
rect 3649 313432 3662 313443
rect 3402 312256 3450 313432
rect 3660 312256 3708 313432
rect 3464 312163 3646 312197
rect 3464 312055 3646 312089
rect 3448 311996 3450 312007
rect 3649 311996 3662 312007
rect 3402 310820 3450 311996
rect 3660 310820 3708 311996
rect 3464 310727 3646 310761
rect 3464 310619 3646 310653
rect 3448 310560 3450 310571
rect 3649 310560 3662 310571
rect 3402 309384 3450 310560
rect 3660 309384 3708 310560
rect 3464 309291 3646 309325
rect 3464 309183 3646 309217
rect 3448 309124 3450 309135
rect 3649 309124 3662 309135
rect 3402 307948 3450 309124
rect 3660 307948 3708 309124
rect 3464 307855 3646 307889
rect 3464 307747 3646 307781
rect 3448 307688 3450 307699
rect 3649 307688 3662 307699
rect 3402 306512 3450 307688
rect 3660 306512 3708 307688
rect 3464 306419 3646 306453
rect 3464 306311 3646 306345
rect 3448 306252 3450 306263
rect 3649 306252 3662 306263
rect 3402 305076 3450 306252
rect 3660 305076 3708 306252
rect 3464 304983 3646 305017
rect 3464 304875 3646 304909
rect 3448 304816 3450 304827
rect 3649 304816 3662 304827
rect 3402 303640 3450 304816
rect 3660 303640 3708 304816
rect 3464 303547 3646 303581
rect 3464 303439 3646 303473
rect 3448 303380 3450 303391
rect 3649 303380 3662 303391
rect 3402 302204 3450 303380
rect 3660 302204 3708 303380
rect 3464 302111 3646 302145
rect 3464 302003 3646 302037
rect 3448 301944 3450 301955
rect 3649 301944 3662 301955
rect 3402 300768 3450 301944
rect 3660 300768 3708 301944
rect 3464 300675 3646 300709
rect 3464 300567 3646 300601
rect 3448 300508 3450 300519
rect 3649 300508 3662 300519
rect 3402 299332 3450 300508
rect 3660 299332 3708 300508
rect 3464 299239 3646 299273
rect 3464 299131 3646 299165
rect 3448 299072 3450 299083
rect 3649 299072 3662 299083
rect 3402 297896 3450 299072
rect 3660 297896 3708 299072
rect 3464 297803 3646 297837
rect 3464 297695 3646 297729
rect 3448 297636 3450 297647
rect 3649 297636 3662 297647
rect 3402 296460 3450 297636
rect 3660 296460 3708 297636
rect 3464 296367 3646 296401
rect 3464 296259 3646 296293
rect 3448 296200 3450 296211
rect 3649 296200 3662 296211
rect 3402 295024 3450 296200
rect 3660 295024 3708 296200
rect 3464 294931 3646 294965
rect 3464 294823 3646 294857
rect 3448 294764 3450 294775
rect 3649 294764 3662 294775
rect 3402 293588 3450 294764
rect 3660 293588 3708 294764
rect 3464 293495 3646 293529
rect 3464 293387 3646 293421
rect 3448 293328 3450 293339
rect 3649 293328 3662 293339
rect 3402 292152 3450 293328
rect 3660 292152 3708 293328
rect 3464 292059 3646 292093
rect 3464 291951 3646 291985
rect 3448 291892 3450 291903
rect 3649 291892 3662 291903
rect 3402 290716 3450 291892
rect 3660 290716 3708 291892
rect 3464 290623 3646 290657
rect 3464 290515 3646 290549
rect 3448 290456 3450 290467
rect 3649 290456 3662 290467
rect 3402 289280 3450 290456
rect 3660 289280 3708 290456
rect 3464 289187 3646 289221
rect 3464 289079 3646 289113
rect 3448 289020 3450 289031
rect 3649 289020 3662 289031
rect 3402 287844 3450 289020
rect 3660 287844 3708 289020
rect 3464 287751 3646 287785
rect 3464 287643 3646 287677
rect 3448 287584 3450 287595
rect 3649 287584 3662 287595
rect 3402 286408 3450 287584
rect 3660 286408 3708 287584
rect 3464 286315 3646 286349
rect 3464 286207 3646 286241
rect 3448 286148 3450 286159
rect 3649 286148 3662 286159
rect 3402 284972 3450 286148
rect 3660 284972 3708 286148
rect 3464 284879 3646 284913
rect 3464 284771 3646 284805
rect 3448 284712 3450 284723
rect 3649 284712 3662 284723
rect 3402 283536 3450 284712
rect 3660 283536 3708 284712
rect 3464 283443 3646 283477
rect 3464 283335 3646 283369
rect 3448 283276 3450 283287
rect 3649 283276 3662 283287
rect 3402 282100 3450 283276
rect 3660 282100 3708 283276
rect 3464 282007 3646 282041
rect 3464 281899 3646 281933
rect 3448 281840 3450 281851
rect 3649 281840 3662 281851
rect 3402 280664 3450 281840
rect 3660 280664 3708 281840
rect 3464 280571 3646 280605
rect 3464 280463 3646 280497
rect 3448 280404 3450 280415
rect 3649 280404 3662 280415
rect 3402 279228 3450 280404
rect 3660 279228 3708 280404
rect 3464 279135 3646 279169
rect 3464 279027 3646 279061
rect 3448 278968 3450 278979
rect 3649 278968 3662 278979
rect 3402 277792 3450 278968
rect 3660 277792 3708 278968
rect 3464 277699 3646 277733
rect 3464 277591 3646 277625
rect 3448 277532 3450 277543
rect 3649 277532 3662 277543
rect 3402 276356 3450 277532
rect 3660 276356 3708 277532
rect 3464 276263 3646 276297
rect 3464 276155 3646 276189
rect 3448 276096 3450 276107
rect 3649 276096 3662 276107
rect 3402 274920 3450 276096
rect 3660 274920 3708 276096
rect 3464 274827 3646 274861
rect 3464 274719 3646 274753
rect 3448 274660 3450 274671
rect 3649 274660 3662 274671
rect 3402 273484 3450 274660
rect 3660 273484 3708 274660
rect 3464 273391 3646 273425
rect 3464 273283 3646 273317
rect 3448 273224 3450 273235
rect 3649 273224 3662 273235
rect 3402 272048 3450 273224
rect 3660 272048 3708 273224
rect 3464 271955 3646 271989
rect 3464 271847 3646 271881
rect 3448 271788 3450 271799
rect 3649 271788 3662 271799
rect 3402 270612 3450 271788
rect 3660 270612 3708 271788
rect 3464 270519 3646 270553
rect 3464 270411 3646 270445
rect 3448 270352 3450 270363
rect 3649 270352 3662 270363
rect 3402 269176 3450 270352
rect 3660 269176 3708 270352
rect 3464 269083 3646 269117
rect 3464 268975 3646 269009
rect 3448 268916 3450 268927
rect 3649 268916 3662 268927
rect 3402 267740 3450 268916
rect 3660 267740 3708 268916
rect 3464 267647 3646 267681
rect 3464 267539 3646 267573
rect 3448 267480 3450 267491
rect 3649 267480 3662 267491
rect 3402 266304 3450 267480
rect 3660 266304 3708 267480
rect 3464 266211 3646 266245
rect 3464 266103 3646 266137
rect 3448 266044 3450 266055
rect 3649 266044 3662 266055
rect 3402 264868 3450 266044
rect 3660 264868 3708 266044
rect 3464 264775 3646 264809
rect 3464 264667 3646 264701
rect 3448 264608 3450 264619
rect 3649 264608 3662 264619
rect 3402 263432 3450 264608
rect 3660 263432 3708 264608
rect 3464 263339 3646 263373
rect 3464 263231 3646 263265
rect 3448 263172 3450 263183
rect 3649 263172 3662 263183
rect 3402 261996 3450 263172
rect 3660 261996 3708 263172
rect 3464 261903 3646 261937
rect 3464 261795 3646 261829
rect 3448 261736 3450 261747
rect 3649 261736 3662 261747
rect 3402 260560 3450 261736
rect 3660 260560 3708 261736
rect 3464 260467 3646 260501
rect 3464 260359 3646 260393
rect 3448 260300 3450 260311
rect 3649 260300 3662 260311
rect 3402 259124 3450 260300
rect 3660 259124 3708 260300
rect 3464 259031 3646 259065
rect 3464 258923 3646 258957
rect 3448 258864 3450 258875
rect 3649 258864 3662 258875
rect 3402 257688 3450 258864
rect 3660 257688 3708 258864
rect 3464 257595 3646 257629
rect 3464 257487 3646 257521
rect 3448 257428 3450 257439
rect 3649 257428 3662 257439
rect 3402 256252 3450 257428
rect 3660 256252 3708 257428
rect 3464 256159 3646 256193
rect 3464 256051 3646 256085
rect 3448 255992 3450 256003
rect 3649 255992 3662 256003
rect 3402 254816 3450 255992
rect 3660 254816 3708 255992
rect 3464 254723 3646 254757
rect 3464 254615 3646 254649
rect 3448 254556 3450 254567
rect 3649 254556 3662 254567
rect 3402 253380 3450 254556
rect 3660 253380 3708 254556
rect 3794 254231 4541 352053
rect 4545 351971 4927 352005
rect 5006 351909 5023 351971
rect 4975 351869 5023 351909
rect 4645 351833 4827 351867
rect 4571 351783 4583 351795
rect 4629 351783 4631 351794
rect 4830 351783 4843 351794
rect 4889 351783 4901 351795
rect 4571 350607 4631 351783
rect 4841 350607 4901 351783
rect 4571 350595 4583 350607
rect 4889 350595 4901 350607
rect 4645 350523 4827 350557
rect 4963 350521 5023 351869
rect 4975 350451 5023 350521
rect 4645 350415 4827 350449
rect 4571 350365 4583 350377
rect 4629 350365 4631 350376
rect 4830 350365 4843 350376
rect 4889 350365 4901 350377
rect 4571 349189 4631 350365
rect 4841 349189 4901 350365
rect 4571 349177 4583 349189
rect 4889 349177 4901 349189
rect 4645 349105 4827 349139
rect 4963 349103 5023 350451
rect 4975 349033 5023 349103
rect 4645 348997 4827 349031
rect 4571 348947 4583 348959
rect 4629 348947 4631 348958
rect 4830 348947 4843 348958
rect 4889 348947 4901 348959
rect 4571 347771 4631 348947
rect 4841 347771 4901 348947
rect 4571 347759 4583 347771
rect 4889 347759 4901 347771
rect 4645 347687 4827 347721
rect 4963 347685 5023 349033
rect 4975 347615 5023 347685
rect 4645 347579 4827 347613
rect 4571 347529 4583 347541
rect 4629 347529 4631 347540
rect 4830 347529 4843 347540
rect 4889 347529 4901 347541
rect 4571 346353 4631 347529
rect 4841 346353 4901 347529
rect 4571 346341 4583 346353
rect 4889 346341 4901 346353
rect 4645 346269 4827 346303
rect 4963 346267 5023 347615
rect 4975 346197 5023 346267
rect 4645 346161 4827 346195
rect 4571 346111 4583 346123
rect 4629 346111 4631 346122
rect 4830 346111 4843 346122
rect 4889 346111 4901 346123
rect 4571 344935 4631 346111
rect 4841 344935 4901 346111
rect 4571 344923 4583 344935
rect 4889 344923 4901 344935
rect 4645 344851 4827 344885
rect 4963 344849 5023 346197
rect 4975 344779 5023 344849
rect 4645 344743 4827 344777
rect 4571 344693 4583 344705
rect 4629 344693 4631 344704
rect 4830 344693 4843 344704
rect 4889 344693 4901 344705
rect 4571 343517 4631 344693
rect 4841 343517 4901 344693
rect 4571 343505 4583 343517
rect 4889 343505 4901 343517
rect 4645 343433 4827 343467
rect 4963 343431 5023 344779
rect 4975 343361 5023 343431
rect 4645 343325 4827 343359
rect 4571 343275 4583 343287
rect 4629 343275 4631 343286
rect 4830 343275 4843 343286
rect 4889 343275 4901 343287
rect 4571 342099 4631 343275
rect 4841 342099 4901 343275
rect 4571 342087 4583 342099
rect 4889 342087 4901 342099
rect 4645 342015 4827 342049
rect 4963 342013 5023 343361
rect 4975 341943 5023 342013
rect 4645 341907 4827 341941
rect 4571 341857 4583 341869
rect 4629 341857 4631 341868
rect 4830 341857 4843 341868
rect 4889 341857 4901 341869
rect 4571 340681 4631 341857
rect 4841 340681 4901 341857
rect 4571 340669 4583 340681
rect 4889 340669 4901 340681
rect 4645 340597 4827 340631
rect 4963 340595 5023 341943
rect 4975 340525 5023 340595
rect 4645 340489 4827 340523
rect 4571 340439 4583 340451
rect 4629 340439 4631 340450
rect 4830 340439 4843 340450
rect 4889 340439 4901 340451
rect 4571 339263 4631 340439
rect 4841 339263 4901 340439
rect 4571 339251 4583 339263
rect 4889 339251 4901 339263
rect 4645 339179 4827 339213
rect 4963 339177 5023 340525
rect 4975 339107 5023 339177
rect 4645 339071 4827 339105
rect 4571 339021 4583 339033
rect 4629 339021 4631 339032
rect 4830 339021 4843 339032
rect 4889 339021 4901 339033
rect 4571 337845 4631 339021
rect 4841 337845 4901 339021
rect 4571 337833 4583 337845
rect 4889 337833 4901 337845
rect 4645 337761 4827 337795
rect 4963 337759 5023 339107
rect 4975 337689 5023 337759
rect 4645 337653 4827 337687
rect 4571 337603 4583 337615
rect 4629 337603 4631 337614
rect 4830 337603 4843 337614
rect 4889 337603 4901 337615
rect 4571 336427 4631 337603
rect 4841 336427 4901 337603
rect 4571 336415 4583 336427
rect 4889 336415 4901 336427
rect 4645 336343 4827 336377
rect 4963 336341 5023 337689
rect 4975 336271 5023 336341
rect 4645 336235 4827 336269
rect 4571 336185 4583 336197
rect 4629 336185 4631 336196
rect 4830 336185 4843 336196
rect 4889 336185 4901 336197
rect 4571 335009 4631 336185
rect 4841 335009 4901 336185
rect 4571 334997 4583 335009
rect 4889 334997 4901 335009
rect 4645 334925 4827 334959
rect 4963 334923 5023 336271
rect 4975 334853 5023 334923
rect 4645 334817 4827 334851
rect 4571 334767 4583 334779
rect 4629 334767 4631 334778
rect 4830 334767 4843 334778
rect 4889 334767 4901 334779
rect 4571 333591 4631 334767
rect 4841 333591 4901 334767
rect 4571 333579 4583 333591
rect 4889 333579 4901 333591
rect 4645 333507 4827 333541
rect 4963 333505 5023 334853
rect 4975 333435 5023 333505
rect 4645 333399 4827 333433
rect 4571 333349 4583 333361
rect 4629 333349 4631 333360
rect 4830 333349 4843 333360
rect 4889 333349 4901 333361
rect 4571 332173 4631 333349
rect 4841 332173 4901 333349
rect 4571 332161 4583 332173
rect 4889 332161 4901 332173
rect 4645 332089 4827 332123
rect 4963 332087 5023 333435
rect 4975 332017 5023 332087
rect 4645 331981 4827 332015
rect 4571 331931 4583 331943
rect 4629 331931 4631 331942
rect 4830 331931 4843 331942
rect 4889 331931 4901 331943
rect 4571 330755 4631 331931
rect 4841 330755 4901 331931
rect 4571 330743 4583 330755
rect 4889 330743 4901 330755
rect 4645 330671 4827 330705
rect 4963 330669 5023 332017
rect 4975 330599 5023 330669
rect 4645 330563 4827 330597
rect 4571 330513 4583 330525
rect 4629 330513 4631 330524
rect 4830 330513 4843 330524
rect 4889 330513 4901 330525
rect 4571 329337 4631 330513
rect 4841 329337 4901 330513
rect 4571 329325 4583 329337
rect 4889 329325 4901 329337
rect 4645 329253 4827 329287
rect 4963 329251 5023 330599
rect 4975 329181 5023 329251
rect 4645 329145 4827 329179
rect 4571 329095 4583 329107
rect 4629 329095 4631 329106
rect 4830 329095 4843 329106
rect 4889 329095 4901 329107
rect 4571 327919 4631 329095
rect 4841 327919 4901 329095
rect 4571 327907 4583 327919
rect 4889 327907 4901 327919
rect 4645 327835 4827 327869
rect 4963 327833 5023 329181
rect 4975 327763 5023 327833
rect 4645 327727 4827 327761
rect 4571 327677 4583 327689
rect 4629 327677 4631 327688
rect 4830 327677 4843 327688
rect 4889 327677 4901 327689
rect 4571 326501 4631 327677
rect 4841 326501 4901 327677
rect 4571 326489 4583 326501
rect 4889 326489 4901 326501
rect 4645 326417 4827 326451
rect 4963 326415 5023 327763
rect 4975 326345 5023 326415
rect 4645 326309 4827 326343
rect 4571 326259 4583 326271
rect 4629 326259 4631 326270
rect 4830 326259 4843 326270
rect 4889 326259 4901 326271
rect 4571 325083 4631 326259
rect 4841 325083 4901 326259
rect 4571 325071 4583 325083
rect 4889 325071 4901 325083
rect 4645 324999 4827 325033
rect 4963 324997 5023 326345
rect 4975 324927 5023 324997
rect 4645 324891 4827 324925
rect 4571 324841 4583 324853
rect 4629 324841 4631 324852
rect 4830 324841 4843 324852
rect 4889 324841 4901 324853
rect 4571 323665 4631 324841
rect 4841 323665 4901 324841
rect 4571 323653 4583 323665
rect 4889 323653 4901 323665
rect 4645 323581 4827 323615
rect 4963 323579 5023 324927
rect 4975 323509 5023 323579
rect 4645 323473 4827 323507
rect 4571 323423 4583 323435
rect 4629 323423 4631 323434
rect 4830 323423 4843 323434
rect 4889 323423 4901 323435
rect 4571 322247 4631 323423
rect 4841 322247 4901 323423
rect 4571 322235 4583 322247
rect 4889 322235 4901 322247
rect 4645 322163 4827 322197
rect 4963 322161 5023 323509
rect 4975 322091 5023 322161
rect 4645 322055 4827 322089
rect 4571 322005 4583 322017
rect 4629 322005 4631 322016
rect 4830 322005 4843 322016
rect 4889 322005 4901 322017
rect 4571 320829 4631 322005
rect 4841 320829 4901 322005
rect 4571 320817 4583 320829
rect 4889 320817 4901 320829
rect 4645 320745 4827 320779
rect 4963 320743 5023 322091
rect 4975 320673 5023 320743
rect 4645 320637 4827 320671
rect 4571 320587 4583 320599
rect 4629 320587 4631 320598
rect 4830 320587 4843 320598
rect 4889 320587 4901 320599
rect 4571 319411 4631 320587
rect 4841 319411 4901 320587
rect 4571 319399 4583 319411
rect 4889 319399 4901 319411
rect 4645 319327 4827 319361
rect 4963 319325 5023 320673
rect 4975 319255 5023 319325
rect 4645 319219 4827 319253
rect 4571 319169 4583 319181
rect 4629 319169 4631 319180
rect 4830 319169 4843 319180
rect 4889 319169 4901 319181
rect 4571 317993 4631 319169
rect 4841 317993 4901 319169
rect 4571 317981 4583 317993
rect 4889 317981 4901 317993
rect 4645 317909 4827 317943
rect 4963 317907 5023 319255
rect 4975 317837 5023 317907
rect 4645 317801 4827 317835
rect 4571 317751 4583 317763
rect 4629 317751 4631 317762
rect 4830 317751 4843 317762
rect 4889 317751 4901 317763
rect 4571 316575 4631 317751
rect 4841 316575 4901 317751
rect 4571 316563 4583 316575
rect 4889 316563 4901 316575
rect 4645 316491 4827 316525
rect 4963 316489 5023 317837
rect 4975 316419 5023 316489
rect 4645 316383 4827 316417
rect 4571 316333 4583 316345
rect 4629 316333 4631 316344
rect 4830 316333 4843 316344
rect 4889 316333 4901 316345
rect 4571 315157 4631 316333
rect 4841 315157 4901 316333
rect 4571 315145 4583 315157
rect 4889 315145 4901 315157
rect 4645 315073 4827 315107
rect 4963 315071 5023 316419
rect 4975 315001 5023 315071
rect 4645 314965 4827 314999
rect 4571 314915 4583 314927
rect 4629 314915 4631 314926
rect 4830 314915 4843 314926
rect 4889 314915 4901 314927
rect 4571 313739 4631 314915
rect 4841 313739 4901 314915
rect 4571 313727 4583 313739
rect 4889 313727 4901 313739
rect 4645 313655 4827 313689
rect 4963 313653 5023 315001
rect 4975 313583 5023 313653
rect 4645 313547 4827 313581
rect 4571 313497 4583 313509
rect 4629 313497 4631 313508
rect 4830 313497 4843 313508
rect 4889 313497 4901 313509
rect 4571 312321 4631 313497
rect 4841 312321 4901 313497
rect 4571 312309 4583 312321
rect 4889 312309 4901 312321
rect 4645 312237 4827 312271
rect 4963 312235 5023 313583
rect 4975 312165 5023 312235
rect 4645 312129 4827 312163
rect 4571 312079 4583 312091
rect 4629 312079 4631 312090
rect 4830 312079 4843 312090
rect 4889 312079 4901 312091
rect 4571 310903 4631 312079
rect 4841 310903 4901 312079
rect 4571 310891 4583 310903
rect 4889 310891 4901 310903
rect 4645 310819 4827 310853
rect 4963 310817 5023 312165
rect 4975 310747 5023 310817
rect 4645 310711 4827 310745
rect 4571 310661 4583 310673
rect 4629 310661 4631 310672
rect 4830 310661 4843 310672
rect 4889 310661 4901 310673
rect 4571 309485 4631 310661
rect 4841 309485 4901 310661
rect 4571 309473 4583 309485
rect 4889 309473 4901 309485
rect 4645 309401 4827 309435
rect 4963 309399 5023 310747
rect 4975 309329 5023 309399
rect 4645 309293 4827 309327
rect 4571 309243 4583 309255
rect 4629 309243 4631 309254
rect 4830 309243 4843 309254
rect 4889 309243 4901 309255
rect 4571 308067 4631 309243
rect 4841 308067 4901 309243
rect 4571 308055 4583 308067
rect 4889 308055 4901 308067
rect 4645 307983 4827 308017
rect 4963 307981 5023 309329
rect 4975 307911 5023 307981
rect 4645 307875 4827 307909
rect 4571 307825 4583 307837
rect 4629 307825 4631 307836
rect 4830 307825 4843 307836
rect 4889 307825 4901 307837
rect 4571 306649 4631 307825
rect 4841 306649 4901 307825
rect 4571 306637 4583 306649
rect 4889 306637 4901 306649
rect 4645 306565 4827 306599
rect 4963 306563 5023 307911
rect 4975 306493 5023 306563
rect 4645 306457 4827 306491
rect 4571 306407 4583 306419
rect 4629 306407 4631 306418
rect 4830 306407 4843 306418
rect 4889 306407 4901 306419
rect 4571 305231 4631 306407
rect 4841 305231 4901 306407
rect 4571 305219 4583 305231
rect 4889 305219 4901 305231
rect 4645 305147 4827 305181
rect 4963 305145 5023 306493
rect 4975 305075 5023 305145
rect 4645 305039 4827 305073
rect 4571 304989 4583 305001
rect 4629 304989 4631 305000
rect 4830 304989 4843 305000
rect 4889 304989 4901 305001
rect 4571 303813 4631 304989
rect 4841 303813 4901 304989
rect 4571 303801 4583 303813
rect 4889 303801 4901 303813
rect 4645 303729 4827 303763
rect 4963 303727 5023 305075
rect 4975 303657 5023 303727
rect 4645 303621 4827 303655
rect 4571 303571 4583 303583
rect 4629 303571 4631 303582
rect 4830 303571 4843 303582
rect 4889 303571 4901 303583
rect 4571 302395 4631 303571
rect 4841 302395 4901 303571
rect 4571 302383 4583 302395
rect 4889 302383 4901 302395
rect 4645 302311 4827 302345
rect 4963 302309 5023 303657
rect 4975 302239 5023 302309
rect 4645 302203 4827 302237
rect 4571 302153 4583 302165
rect 4629 302153 4631 302164
rect 4830 302153 4843 302164
rect 4889 302153 4901 302165
rect 4571 300977 4631 302153
rect 4841 300977 4901 302153
rect 4571 300965 4583 300977
rect 4889 300965 4901 300977
rect 4645 300893 4827 300927
rect 4963 300891 5023 302239
rect 4975 300821 5023 300891
rect 4645 300785 4827 300819
rect 4571 300735 4583 300747
rect 4629 300735 4631 300746
rect 4830 300735 4843 300746
rect 4889 300735 4901 300747
rect 4571 299559 4631 300735
rect 4841 299559 4901 300735
rect 4571 299547 4583 299559
rect 4889 299547 4901 299559
rect 4645 299475 4827 299509
rect 4963 299473 5023 300821
rect 4975 299403 5023 299473
rect 4645 299367 4827 299401
rect 4571 299317 4583 299329
rect 4629 299317 4631 299328
rect 4830 299317 4843 299328
rect 4889 299317 4901 299329
rect 4571 298141 4631 299317
rect 4841 298141 4901 299317
rect 4571 298129 4583 298141
rect 4889 298129 4901 298141
rect 4645 298057 4827 298091
rect 4963 298055 5023 299403
rect 4975 297985 5023 298055
rect 4645 297949 4827 297983
rect 4571 297899 4583 297911
rect 4629 297899 4631 297910
rect 4830 297899 4843 297910
rect 4889 297899 4901 297911
rect 4571 296723 4631 297899
rect 4841 296723 4901 297899
rect 4571 296711 4583 296723
rect 4889 296711 4901 296723
rect 4645 296639 4827 296673
rect 4963 296637 5023 297985
rect 4975 296567 5023 296637
rect 4645 296531 4827 296565
rect 4571 296481 4583 296493
rect 4629 296481 4631 296492
rect 4830 296481 4843 296492
rect 4889 296481 4901 296493
rect 4571 295305 4631 296481
rect 4841 295305 4901 296481
rect 4571 295293 4583 295305
rect 4889 295293 4901 295305
rect 4645 295221 4827 295255
rect 4963 295219 5023 296567
rect 4975 295149 5023 295219
rect 4645 295113 4827 295147
rect 4571 295063 4583 295075
rect 4629 295063 4631 295074
rect 4830 295063 4843 295074
rect 4889 295063 4901 295075
rect 4571 293887 4631 295063
rect 4841 293887 4901 295063
rect 4571 293875 4583 293887
rect 4889 293875 4901 293887
rect 4645 293803 4827 293837
rect 4963 293801 5023 295149
rect 4975 293731 5023 293801
rect 4645 293695 4827 293729
rect 4571 293645 4583 293657
rect 4629 293645 4631 293656
rect 4830 293645 4843 293656
rect 4889 293645 4901 293657
rect 4571 292469 4631 293645
rect 4841 292469 4901 293645
rect 4571 292457 4583 292469
rect 4889 292457 4901 292469
rect 4645 292385 4827 292419
rect 4963 292383 5023 293731
rect 4975 292313 5023 292383
rect 4645 292277 4827 292311
rect 4571 292227 4583 292239
rect 4629 292227 4631 292238
rect 4830 292227 4843 292238
rect 4889 292227 4901 292239
rect 4571 291051 4631 292227
rect 4841 291051 4901 292227
rect 4571 291039 4583 291051
rect 4889 291039 4901 291051
rect 4645 290967 4827 291001
rect 4963 290965 5023 292313
rect 4975 290895 5023 290965
rect 4645 290859 4827 290893
rect 4571 290809 4583 290821
rect 4629 290809 4631 290820
rect 4830 290809 4843 290820
rect 4889 290809 4901 290821
rect 4571 289633 4631 290809
rect 4841 289633 4901 290809
rect 4571 289621 4583 289633
rect 4889 289621 4901 289633
rect 4645 289549 4827 289583
rect 4963 289547 5023 290895
rect 4975 289477 5023 289547
rect 4645 289441 4827 289475
rect 4571 289391 4583 289403
rect 4629 289391 4631 289402
rect 4830 289391 4843 289402
rect 4889 289391 4901 289403
rect 4571 288215 4631 289391
rect 4841 288215 4901 289391
rect 4571 288203 4583 288215
rect 4889 288203 4901 288215
rect 4645 288131 4827 288165
rect 4963 288129 5023 289477
rect 4975 288059 5023 288129
rect 4645 288023 4827 288057
rect 4571 287973 4583 287985
rect 4629 287973 4631 287984
rect 4830 287973 4843 287984
rect 4889 287973 4901 287985
rect 4571 286797 4631 287973
rect 4841 286797 4901 287973
rect 4571 286785 4583 286797
rect 4889 286785 4901 286797
rect 4645 286713 4827 286747
rect 4963 286711 5023 288059
rect 4975 286641 5023 286711
rect 4645 286605 4827 286639
rect 4571 286555 4583 286567
rect 4629 286555 4631 286566
rect 4830 286555 4843 286566
rect 4889 286555 4901 286567
rect 4571 285379 4631 286555
rect 4841 285379 4901 286555
rect 4571 285367 4583 285379
rect 4889 285367 4901 285379
rect 4645 285295 4827 285329
rect 4963 285293 5023 286641
rect 4975 285223 5023 285293
rect 4645 285187 4827 285221
rect 4571 285137 4583 285149
rect 4629 285137 4631 285148
rect 4830 285137 4843 285148
rect 4889 285137 4901 285149
rect 4571 283961 4631 285137
rect 4841 283961 4901 285137
rect 4571 283949 4583 283961
rect 4889 283949 4901 283961
rect 4645 283877 4827 283911
rect 4963 283875 5023 285223
rect 4975 283805 5023 283875
rect 4645 283769 4827 283803
rect 4571 283719 4583 283731
rect 4629 283719 4631 283730
rect 4830 283719 4843 283730
rect 4889 283719 4901 283731
rect 4571 282543 4631 283719
rect 4841 282543 4901 283719
rect 4571 282531 4583 282543
rect 4889 282531 4901 282543
rect 4645 282459 4827 282493
rect 4963 282457 5023 283805
rect 4975 282387 5023 282457
rect 4645 282351 4827 282385
rect 4571 282301 4583 282313
rect 4629 282301 4631 282312
rect 4830 282301 4843 282312
rect 4889 282301 4901 282313
rect 4571 281125 4631 282301
rect 4841 281125 4901 282301
rect 4571 281113 4583 281125
rect 4889 281113 4901 281125
rect 4645 281041 4827 281075
rect 4963 281039 5023 282387
rect 4975 280969 5023 281039
rect 4645 280933 4827 280967
rect 4571 280883 4583 280895
rect 4629 280883 4631 280894
rect 4830 280883 4843 280894
rect 4889 280883 4901 280895
rect 4571 279707 4631 280883
rect 4841 279707 4901 280883
rect 4571 279695 4583 279707
rect 4889 279695 4901 279707
rect 4645 279623 4827 279657
rect 4963 279621 5023 280969
rect 4975 279551 5023 279621
rect 4645 279515 4827 279549
rect 4571 279465 4583 279477
rect 4629 279465 4631 279476
rect 4830 279465 4843 279476
rect 4889 279465 4901 279477
rect 4571 278289 4631 279465
rect 4841 278289 4901 279465
rect 4571 278277 4583 278289
rect 4889 278277 4901 278289
rect 4645 278205 4827 278239
rect 4963 278203 5023 279551
rect 4975 278133 5023 278203
rect 4645 278097 4827 278131
rect 4571 278047 4583 278059
rect 4629 278047 4631 278058
rect 4830 278047 4843 278058
rect 4889 278047 4901 278059
rect 4571 276871 4631 278047
rect 4841 276871 4901 278047
rect 4571 276859 4583 276871
rect 4889 276859 4901 276871
rect 4645 276787 4827 276821
rect 4963 276785 5023 278133
rect 4975 276715 5023 276785
rect 4645 276679 4827 276713
rect 4571 276629 4583 276641
rect 4629 276629 4631 276640
rect 4830 276629 4843 276640
rect 4889 276629 4901 276641
rect 4571 275453 4631 276629
rect 4841 275453 4901 276629
rect 4571 275441 4583 275453
rect 4889 275441 4901 275453
rect 4645 275369 4827 275403
rect 4963 275367 5023 276715
rect 4975 275297 5023 275367
rect 4645 275261 4827 275295
rect 4571 275211 4583 275223
rect 4629 275211 4631 275222
rect 4830 275211 4843 275222
rect 4889 275211 4901 275223
rect 4571 274035 4631 275211
rect 4841 274035 4901 275211
rect 4571 274023 4583 274035
rect 4889 274023 4901 274035
rect 4645 273951 4827 273985
rect 4963 273949 5023 275297
rect 4975 273879 5023 273949
rect 4645 273843 4827 273877
rect 4571 273793 4583 273805
rect 4629 273793 4631 273804
rect 4830 273793 4843 273804
rect 4889 273793 4901 273805
rect 4571 272617 4631 273793
rect 4841 272617 4901 273793
rect 4571 272605 4583 272617
rect 4889 272605 4901 272617
rect 4645 272533 4827 272567
rect 4963 272531 5023 273879
rect 4975 272461 5023 272531
rect 4645 272425 4827 272459
rect 4571 272375 4583 272387
rect 4629 272375 4631 272386
rect 4830 272375 4843 272386
rect 4889 272375 4901 272387
rect 4571 271199 4631 272375
rect 4841 271199 4901 272375
rect 4571 271187 4583 271199
rect 4889 271187 4901 271199
rect 4645 271115 4827 271149
rect 4963 271113 5023 272461
rect 4975 271043 5023 271113
rect 4645 271007 4827 271041
rect 4571 270957 4583 270969
rect 4629 270957 4631 270968
rect 4830 270957 4843 270968
rect 4889 270957 4901 270969
rect 4571 269781 4631 270957
rect 4841 269781 4901 270957
rect 4571 269769 4583 269781
rect 4889 269769 4901 269781
rect 4645 269697 4827 269731
rect 4963 269695 5023 271043
rect 4975 269625 5023 269695
rect 4645 269589 4827 269623
rect 4571 269539 4583 269551
rect 4629 269539 4631 269550
rect 4830 269539 4843 269550
rect 4889 269539 4901 269551
rect 4571 268363 4631 269539
rect 4841 268363 4901 269539
rect 4571 268351 4583 268363
rect 4889 268351 4901 268363
rect 4645 268279 4827 268313
rect 4963 268277 5023 269625
rect 4975 268207 5023 268277
rect 4645 268171 4827 268205
rect 4571 268121 4583 268133
rect 4629 268121 4631 268132
rect 4830 268121 4843 268132
rect 4889 268121 4901 268133
rect 4571 266945 4631 268121
rect 4841 266945 4901 268121
rect 4571 266933 4583 266945
rect 4889 266933 4901 266945
rect 4645 266861 4827 266895
rect 4963 266859 5023 268207
rect 4975 266789 5023 266859
rect 4645 266753 4827 266787
rect 4571 266703 4583 266715
rect 4629 266703 4631 266714
rect 4830 266703 4843 266714
rect 4889 266703 4901 266715
rect 4571 265527 4631 266703
rect 4841 265527 4901 266703
rect 4571 265515 4583 265527
rect 4889 265515 4901 265527
rect 4645 265443 4827 265477
rect 4963 265441 5023 266789
rect 4975 265371 5023 265441
rect 4645 265335 4827 265369
rect 4571 265285 4583 265297
rect 4629 265285 4631 265296
rect 4830 265285 4843 265296
rect 4889 265285 4901 265297
rect 4571 264109 4631 265285
rect 4841 264109 4901 265285
rect 4571 264097 4583 264109
rect 4889 264097 4901 264109
rect 4645 264025 4827 264059
rect 4963 264023 5023 265371
rect 4975 263953 5023 264023
rect 4645 263917 4827 263951
rect 4571 263867 4583 263879
rect 4629 263867 4631 263878
rect 4830 263867 4843 263878
rect 4889 263867 4901 263879
rect 4571 262691 4631 263867
rect 4841 262691 4901 263867
rect 4571 262679 4583 262691
rect 4889 262679 4901 262691
rect 4645 262607 4827 262641
rect 4963 262605 5023 263953
rect 4975 262535 5023 262605
rect 4645 262499 4827 262533
rect 4571 262449 4583 262461
rect 4629 262449 4631 262460
rect 4830 262449 4843 262460
rect 4889 262449 4901 262461
rect 4571 261273 4631 262449
rect 4841 261273 4901 262449
rect 4571 261261 4583 261273
rect 4889 261261 4901 261273
rect 4645 261189 4827 261223
rect 4963 261187 5023 262535
rect 4975 261117 5023 261187
rect 4645 261081 4827 261115
rect 4571 261031 4583 261043
rect 4629 261031 4631 261042
rect 4830 261031 4843 261042
rect 4889 261031 4901 261043
rect 4571 259855 4631 261031
rect 4841 259855 4901 261031
rect 4571 259843 4583 259855
rect 4889 259843 4901 259855
rect 4645 259771 4827 259805
rect 4963 259769 5023 261117
rect 4975 259699 5023 259769
rect 4645 259663 4827 259697
rect 4571 259613 4583 259625
rect 4629 259613 4631 259624
rect 4830 259613 4843 259624
rect 4889 259613 4901 259625
rect 4571 258437 4631 259613
rect 4841 258437 4901 259613
rect 4571 258425 4583 258437
rect 4889 258425 4901 258437
rect 4645 258353 4827 258387
rect 4963 258351 5023 259699
rect 4975 258281 5023 258351
rect 4645 258245 4827 258279
rect 4571 258195 4583 258207
rect 4629 258195 4631 258206
rect 4830 258195 4843 258206
rect 4889 258195 4901 258207
rect 4571 257019 4631 258195
rect 4841 257019 4901 258195
rect 4571 257007 4583 257019
rect 4889 257007 4901 257019
rect 4645 256935 4827 256969
rect 4963 256933 5023 258281
rect 4975 256863 5023 256933
rect 4645 256827 4827 256861
rect 4571 256777 4583 256789
rect 4629 256777 4631 256788
rect 4830 256777 4843 256788
rect 4889 256777 4901 256789
rect 4571 255601 4631 256777
rect 4841 255601 4901 256777
rect 4571 255589 4583 255601
rect 4889 255589 4901 255601
rect 4645 255517 4827 255551
rect 4963 255515 5023 256863
rect 4975 255445 5023 255515
rect 4645 255409 4827 255443
rect 4571 255359 4583 255371
rect 4629 255359 4631 255370
rect 4830 255359 4843 255370
rect 4889 255359 4901 255371
rect 4571 254231 4631 255359
rect 4841 254231 4901 255359
rect 4963 254231 5023 255445
rect 5040 351844 5057 351940
rect 5136 351906 5518 351940
rect 5040 351804 5088 351844
rect 5566 351804 5614 351844
rect 5040 350456 5100 351804
rect 5236 351768 5418 351802
rect 5162 351718 5174 351730
rect 5220 351718 5222 351729
rect 5421 351718 5434 351729
rect 5480 351718 5492 351730
rect 5162 350542 5222 351718
rect 5432 350542 5492 351718
rect 5162 350530 5174 350542
rect 5480 350530 5492 350542
rect 5236 350458 5418 350492
rect 5554 350456 5614 351804
rect 5040 350386 5088 350456
rect 5566 350386 5614 350456
rect 5040 349038 5100 350386
rect 5236 350350 5418 350384
rect 5162 350300 5174 350312
rect 5220 350300 5222 350311
rect 5421 350300 5434 350311
rect 5480 350300 5492 350312
rect 5162 349124 5222 350300
rect 5432 349124 5492 350300
rect 5162 349112 5174 349124
rect 5480 349112 5492 349124
rect 5236 349040 5418 349074
rect 5554 349038 5614 350386
rect 5040 348968 5088 349038
rect 5566 348968 5614 349038
rect 5040 347620 5100 348968
rect 5236 348932 5418 348966
rect 5162 348882 5174 348894
rect 5220 348882 5222 348893
rect 5421 348882 5434 348893
rect 5480 348882 5492 348894
rect 5162 347706 5222 348882
rect 5432 347706 5492 348882
rect 5162 347694 5174 347706
rect 5480 347694 5492 347706
rect 5236 347622 5418 347656
rect 5554 347620 5614 348968
rect 5040 347550 5088 347620
rect 5566 347550 5614 347620
rect 5040 346202 5100 347550
rect 5236 347514 5418 347548
rect 5162 347464 5174 347476
rect 5220 347464 5222 347475
rect 5421 347464 5434 347475
rect 5480 347464 5492 347476
rect 5162 346288 5222 347464
rect 5432 346288 5492 347464
rect 5162 346276 5174 346288
rect 5480 346276 5492 346288
rect 5236 346204 5418 346238
rect 5554 346202 5614 347550
rect 5040 346132 5088 346202
rect 5566 346132 5614 346202
rect 5040 344784 5100 346132
rect 5236 346096 5418 346130
rect 5162 346046 5174 346058
rect 5220 346046 5222 346057
rect 5421 346046 5434 346057
rect 5480 346046 5492 346058
rect 5162 344870 5222 346046
rect 5432 344870 5492 346046
rect 5162 344858 5174 344870
rect 5480 344858 5492 344870
rect 5236 344786 5418 344820
rect 5554 344784 5614 346132
rect 5040 344714 5088 344784
rect 5566 344714 5614 344784
rect 5040 343366 5100 344714
rect 5236 344678 5418 344712
rect 5162 344628 5174 344640
rect 5220 344628 5222 344639
rect 5421 344628 5434 344639
rect 5480 344628 5492 344640
rect 5162 343452 5222 344628
rect 5432 343452 5492 344628
rect 5162 343440 5174 343452
rect 5480 343440 5492 343452
rect 5236 343368 5418 343402
rect 5554 343366 5614 344714
rect 5040 343296 5088 343366
rect 5566 343296 5614 343366
rect 5040 341948 5100 343296
rect 5236 343260 5418 343294
rect 5162 343210 5174 343222
rect 5220 343210 5222 343221
rect 5421 343210 5434 343221
rect 5480 343210 5492 343222
rect 5162 342034 5222 343210
rect 5432 342034 5492 343210
rect 5162 342022 5174 342034
rect 5480 342022 5492 342034
rect 5236 341950 5418 341984
rect 5554 341948 5614 343296
rect 5040 341878 5088 341948
rect 5566 341878 5614 341948
rect 5040 340530 5100 341878
rect 5236 341842 5418 341876
rect 5162 341792 5174 341804
rect 5220 341792 5222 341803
rect 5421 341792 5434 341803
rect 5480 341792 5492 341804
rect 5162 340616 5222 341792
rect 5432 340616 5492 341792
rect 5162 340604 5174 340616
rect 5480 340604 5492 340616
rect 5236 340532 5418 340566
rect 5554 340530 5614 341878
rect 5040 340460 5088 340530
rect 5566 340460 5614 340530
rect 5040 339112 5100 340460
rect 5236 340424 5418 340458
rect 5162 340374 5174 340386
rect 5220 340374 5222 340385
rect 5421 340374 5434 340385
rect 5480 340374 5492 340386
rect 5162 339198 5222 340374
rect 5432 339198 5492 340374
rect 5162 339186 5174 339198
rect 5480 339186 5492 339198
rect 5236 339114 5418 339148
rect 5554 339112 5614 340460
rect 5040 339042 5088 339112
rect 5566 339042 5614 339112
rect 5040 337694 5100 339042
rect 5236 339006 5418 339040
rect 5162 338956 5174 338968
rect 5220 338956 5222 338967
rect 5421 338956 5434 338967
rect 5480 338956 5492 338968
rect 5162 337780 5222 338956
rect 5432 337780 5492 338956
rect 5162 337768 5174 337780
rect 5480 337768 5492 337780
rect 5236 337696 5418 337730
rect 5554 337694 5614 339042
rect 5040 337624 5088 337694
rect 5566 337624 5614 337694
rect 5040 336276 5100 337624
rect 5236 337588 5418 337622
rect 5162 337538 5174 337550
rect 5220 337538 5222 337549
rect 5421 337538 5434 337549
rect 5480 337538 5492 337550
rect 5162 336362 5222 337538
rect 5432 336362 5492 337538
rect 5162 336350 5174 336362
rect 5480 336350 5492 336362
rect 5236 336278 5418 336312
rect 5554 336276 5614 337624
rect 5040 336206 5088 336276
rect 5566 336206 5614 336276
rect 5040 334858 5100 336206
rect 5236 336170 5418 336204
rect 5162 336120 5174 336132
rect 5220 336120 5222 336131
rect 5421 336120 5434 336131
rect 5480 336120 5492 336132
rect 5162 334944 5222 336120
rect 5432 334944 5492 336120
rect 5162 334932 5174 334944
rect 5480 334932 5492 334944
rect 5236 334860 5418 334894
rect 5554 334858 5614 336206
rect 5040 334788 5088 334858
rect 5566 334788 5614 334858
rect 5040 333440 5100 334788
rect 5236 334752 5418 334786
rect 5162 334702 5174 334714
rect 5220 334702 5222 334713
rect 5421 334702 5434 334713
rect 5480 334702 5492 334714
rect 5162 333526 5222 334702
rect 5432 333526 5492 334702
rect 5162 333514 5174 333526
rect 5480 333514 5492 333526
rect 5236 333442 5418 333476
rect 5554 333440 5614 334788
rect 5040 333370 5088 333440
rect 5566 333370 5614 333440
rect 5040 332022 5100 333370
rect 5236 333334 5418 333368
rect 5162 333284 5174 333296
rect 5220 333284 5222 333295
rect 5421 333284 5434 333295
rect 5480 333284 5492 333296
rect 5162 332108 5222 333284
rect 5432 332108 5492 333284
rect 5162 332096 5174 332108
rect 5480 332096 5492 332108
rect 5236 332024 5418 332058
rect 5554 332022 5614 333370
rect 5040 331952 5088 332022
rect 5566 331952 5614 332022
rect 5040 330604 5100 331952
rect 5236 331916 5418 331950
rect 5162 331866 5174 331878
rect 5220 331866 5222 331877
rect 5421 331866 5434 331877
rect 5480 331866 5492 331878
rect 5162 330690 5222 331866
rect 5432 330690 5492 331866
rect 5162 330678 5174 330690
rect 5480 330678 5492 330690
rect 5236 330606 5418 330640
rect 5554 330604 5614 331952
rect 5040 330534 5088 330604
rect 5566 330534 5614 330604
rect 5040 329186 5100 330534
rect 5236 330498 5418 330532
rect 5162 330448 5174 330460
rect 5220 330448 5222 330459
rect 5421 330448 5434 330459
rect 5480 330448 5492 330460
rect 5162 329272 5222 330448
rect 5432 329272 5492 330448
rect 5162 329260 5174 329272
rect 5480 329260 5492 329272
rect 5236 329188 5418 329222
rect 5554 329186 5614 330534
rect 5040 329116 5088 329186
rect 5566 329116 5614 329186
rect 5040 327768 5100 329116
rect 5236 329080 5418 329114
rect 5162 329030 5174 329042
rect 5220 329030 5222 329041
rect 5421 329030 5434 329041
rect 5480 329030 5492 329042
rect 5162 327854 5222 329030
rect 5432 327854 5492 329030
rect 5162 327842 5174 327854
rect 5480 327842 5492 327854
rect 5236 327770 5418 327804
rect 5554 327768 5614 329116
rect 5040 327698 5088 327768
rect 5566 327698 5614 327768
rect 5040 326350 5100 327698
rect 5236 327662 5418 327696
rect 5162 327612 5174 327624
rect 5220 327612 5222 327623
rect 5421 327612 5434 327623
rect 5480 327612 5492 327624
rect 5162 326436 5222 327612
rect 5432 326436 5492 327612
rect 5162 326424 5174 326436
rect 5480 326424 5492 326436
rect 5236 326352 5418 326386
rect 5554 326350 5614 327698
rect 5040 326280 5088 326350
rect 5566 326280 5614 326350
rect 5040 324932 5100 326280
rect 5236 326244 5418 326278
rect 5162 326194 5174 326206
rect 5220 326194 5222 326205
rect 5421 326194 5434 326205
rect 5480 326194 5492 326206
rect 5162 325018 5222 326194
rect 5432 325018 5492 326194
rect 5162 325006 5174 325018
rect 5480 325006 5492 325018
rect 5236 324934 5418 324968
rect 5554 324932 5614 326280
rect 5040 324862 5088 324932
rect 5566 324862 5614 324932
rect 5040 323514 5100 324862
rect 5236 324826 5418 324860
rect 5162 324776 5174 324788
rect 5220 324776 5222 324787
rect 5421 324776 5434 324787
rect 5480 324776 5492 324788
rect 5162 323600 5222 324776
rect 5432 323600 5492 324776
rect 5162 323588 5174 323600
rect 5480 323588 5492 323600
rect 5236 323516 5418 323550
rect 5554 323514 5614 324862
rect 5040 323444 5088 323514
rect 5566 323444 5614 323514
rect 5040 322096 5100 323444
rect 5236 323408 5418 323442
rect 5162 323358 5174 323370
rect 5220 323358 5222 323369
rect 5421 323358 5434 323369
rect 5480 323358 5492 323370
rect 5162 322182 5222 323358
rect 5432 322182 5492 323358
rect 5162 322170 5174 322182
rect 5480 322170 5492 322182
rect 5236 322098 5418 322132
rect 5554 322096 5614 323444
rect 5040 322026 5088 322096
rect 5566 322026 5614 322096
rect 5040 320678 5100 322026
rect 5236 321990 5418 322024
rect 5162 321940 5174 321952
rect 5220 321940 5222 321951
rect 5421 321940 5434 321951
rect 5480 321940 5492 321952
rect 5162 320764 5222 321940
rect 5432 320764 5492 321940
rect 5162 320752 5174 320764
rect 5480 320752 5492 320764
rect 5236 320680 5418 320714
rect 5554 320678 5614 322026
rect 5040 320608 5088 320678
rect 5566 320608 5614 320678
rect 5040 319260 5100 320608
rect 5236 320572 5418 320606
rect 5162 320522 5174 320534
rect 5220 320522 5222 320533
rect 5421 320522 5434 320533
rect 5480 320522 5492 320534
rect 5162 319346 5222 320522
rect 5432 319346 5492 320522
rect 5162 319334 5174 319346
rect 5480 319334 5492 319346
rect 5236 319262 5418 319296
rect 5554 319260 5614 320608
rect 5040 319190 5088 319260
rect 5566 319190 5614 319260
rect 5040 317842 5100 319190
rect 5236 319154 5418 319188
rect 5162 319104 5174 319116
rect 5220 319104 5222 319115
rect 5421 319104 5434 319115
rect 5480 319104 5492 319116
rect 5162 317928 5222 319104
rect 5432 317928 5492 319104
rect 5162 317916 5174 317928
rect 5480 317916 5492 317928
rect 5236 317844 5418 317878
rect 5554 317842 5614 319190
rect 5040 317772 5088 317842
rect 5566 317772 5614 317842
rect 5040 316424 5100 317772
rect 5236 317736 5418 317770
rect 5162 317686 5174 317698
rect 5220 317686 5222 317697
rect 5421 317686 5434 317697
rect 5480 317686 5492 317698
rect 5162 316510 5222 317686
rect 5432 316510 5492 317686
rect 5162 316498 5174 316510
rect 5480 316498 5492 316510
rect 5236 316426 5418 316460
rect 5554 316424 5614 317772
rect 5040 316354 5088 316424
rect 5566 316354 5614 316424
rect 5040 315006 5100 316354
rect 5236 316318 5418 316352
rect 5162 316268 5174 316280
rect 5220 316268 5222 316279
rect 5421 316268 5434 316279
rect 5480 316268 5492 316280
rect 5162 315092 5222 316268
rect 5432 315092 5492 316268
rect 5162 315080 5174 315092
rect 5480 315080 5492 315092
rect 5236 315008 5418 315042
rect 5554 315006 5614 316354
rect 5040 314936 5088 315006
rect 5566 314936 5614 315006
rect 5040 313588 5100 314936
rect 5236 314900 5418 314934
rect 5162 314850 5174 314862
rect 5220 314850 5222 314861
rect 5421 314850 5434 314861
rect 5480 314850 5492 314862
rect 5162 313674 5222 314850
rect 5432 313674 5492 314850
rect 5162 313662 5174 313674
rect 5480 313662 5492 313674
rect 5236 313590 5418 313624
rect 5554 313588 5614 314936
rect 5040 313518 5088 313588
rect 5566 313518 5614 313588
rect 5040 312170 5100 313518
rect 5236 313482 5418 313516
rect 5162 313432 5174 313444
rect 5220 313432 5222 313443
rect 5421 313432 5434 313443
rect 5480 313432 5492 313444
rect 5162 312256 5222 313432
rect 5432 312256 5492 313432
rect 5162 312244 5174 312256
rect 5480 312244 5492 312256
rect 5236 312172 5418 312206
rect 5554 312170 5614 313518
rect 5040 312100 5088 312170
rect 5566 312100 5614 312170
rect 5040 310752 5100 312100
rect 5236 312064 5418 312098
rect 5162 312014 5174 312026
rect 5220 312014 5222 312025
rect 5421 312014 5434 312025
rect 5480 312014 5492 312026
rect 5162 310838 5222 312014
rect 5432 310838 5492 312014
rect 5162 310826 5174 310838
rect 5480 310826 5492 310838
rect 5236 310754 5418 310788
rect 5554 310752 5614 312100
rect 5040 310682 5088 310752
rect 5566 310682 5614 310752
rect 5040 309334 5100 310682
rect 5236 310646 5418 310680
rect 5162 310596 5174 310608
rect 5220 310596 5222 310607
rect 5421 310596 5434 310607
rect 5480 310596 5492 310608
rect 5162 309420 5222 310596
rect 5432 309420 5492 310596
rect 5162 309408 5174 309420
rect 5480 309408 5492 309420
rect 5236 309336 5418 309370
rect 5554 309334 5614 310682
rect 5040 309264 5088 309334
rect 5566 309264 5614 309334
rect 5040 307916 5100 309264
rect 5236 309228 5418 309262
rect 5162 309178 5174 309190
rect 5220 309178 5222 309189
rect 5421 309178 5434 309189
rect 5480 309178 5492 309190
rect 5162 308002 5222 309178
rect 5432 308002 5492 309178
rect 5162 307990 5174 308002
rect 5480 307990 5492 308002
rect 5236 307918 5418 307952
rect 5554 307916 5614 309264
rect 5040 307846 5088 307916
rect 5566 307846 5614 307916
rect 5040 306498 5100 307846
rect 5236 307810 5418 307844
rect 5162 307760 5174 307772
rect 5220 307760 5222 307771
rect 5421 307760 5434 307771
rect 5480 307760 5492 307772
rect 5162 306584 5222 307760
rect 5432 306584 5492 307760
rect 5162 306572 5174 306584
rect 5480 306572 5492 306584
rect 5236 306500 5418 306534
rect 5554 306498 5614 307846
rect 5040 306428 5088 306498
rect 5566 306428 5614 306498
rect 5040 305080 5100 306428
rect 5236 306392 5418 306426
rect 5162 306342 5174 306354
rect 5220 306342 5222 306353
rect 5421 306342 5434 306353
rect 5480 306342 5492 306354
rect 5162 305166 5222 306342
rect 5432 305166 5492 306342
rect 5162 305154 5174 305166
rect 5480 305154 5492 305166
rect 5236 305082 5418 305116
rect 5554 305080 5614 306428
rect 5040 305010 5088 305080
rect 5566 305010 5614 305080
rect 5040 303662 5100 305010
rect 5236 304974 5418 305008
rect 5162 304924 5174 304936
rect 5220 304924 5222 304935
rect 5421 304924 5434 304935
rect 5480 304924 5492 304936
rect 5162 303748 5222 304924
rect 5432 303748 5492 304924
rect 5162 303736 5174 303748
rect 5480 303736 5492 303748
rect 5236 303664 5418 303698
rect 5554 303662 5614 305010
rect 5040 303592 5088 303662
rect 5566 303592 5614 303662
rect 5040 302244 5100 303592
rect 5236 303556 5418 303590
rect 5162 303506 5174 303518
rect 5220 303506 5222 303517
rect 5421 303506 5434 303517
rect 5480 303506 5492 303518
rect 5162 302330 5222 303506
rect 5432 302330 5492 303506
rect 5162 302318 5174 302330
rect 5480 302318 5492 302330
rect 5236 302246 5418 302280
rect 5554 302244 5614 303592
rect 5040 302174 5088 302244
rect 5566 302174 5614 302244
rect 5040 300826 5100 302174
rect 5236 302138 5418 302172
rect 5162 302088 5174 302100
rect 5220 302088 5222 302099
rect 5421 302088 5434 302099
rect 5480 302088 5492 302100
rect 5162 300912 5222 302088
rect 5432 300912 5492 302088
rect 5162 300900 5174 300912
rect 5480 300900 5492 300912
rect 5236 300828 5418 300862
rect 5554 300826 5614 302174
rect 5040 300756 5088 300826
rect 5566 300756 5614 300826
rect 5040 299408 5100 300756
rect 5236 300720 5418 300754
rect 5162 300670 5174 300682
rect 5220 300670 5222 300681
rect 5421 300670 5434 300681
rect 5480 300670 5492 300682
rect 5162 299494 5222 300670
rect 5432 299494 5492 300670
rect 5162 299482 5174 299494
rect 5480 299482 5492 299494
rect 5236 299410 5418 299444
rect 5554 299408 5614 300756
rect 5040 299338 5088 299408
rect 5566 299338 5614 299408
rect 5040 297990 5100 299338
rect 5236 299302 5418 299336
rect 5162 299252 5174 299264
rect 5220 299252 5222 299263
rect 5421 299252 5434 299263
rect 5480 299252 5492 299264
rect 5162 298076 5222 299252
rect 5432 298076 5492 299252
rect 5162 298064 5174 298076
rect 5480 298064 5492 298076
rect 5236 297992 5418 298026
rect 5554 297990 5614 299338
rect 5040 297920 5088 297990
rect 5566 297920 5614 297990
rect 5040 296572 5100 297920
rect 5236 297884 5418 297918
rect 5162 297834 5174 297846
rect 5220 297834 5222 297845
rect 5421 297834 5434 297845
rect 5480 297834 5492 297846
rect 5162 296658 5222 297834
rect 5432 296658 5492 297834
rect 5162 296646 5174 296658
rect 5480 296646 5492 296658
rect 5236 296574 5418 296608
rect 5554 296572 5614 297920
rect 5040 296502 5088 296572
rect 5566 296502 5614 296572
rect 5040 295154 5100 296502
rect 5236 296466 5418 296500
rect 5162 296416 5174 296428
rect 5220 296416 5222 296427
rect 5421 296416 5434 296427
rect 5480 296416 5492 296428
rect 5162 295240 5222 296416
rect 5432 295240 5492 296416
rect 5162 295228 5174 295240
rect 5480 295228 5492 295240
rect 5236 295156 5418 295190
rect 5554 295154 5614 296502
rect 5040 295084 5088 295154
rect 5566 295084 5614 295154
rect 5040 293736 5100 295084
rect 5236 295048 5418 295082
rect 5162 294998 5174 295010
rect 5220 294998 5222 295009
rect 5421 294998 5434 295009
rect 5480 294998 5492 295010
rect 5162 293822 5222 294998
rect 5432 293822 5492 294998
rect 5162 293810 5174 293822
rect 5480 293810 5492 293822
rect 5236 293738 5418 293772
rect 5554 293736 5614 295084
rect 5040 293666 5088 293736
rect 5566 293666 5614 293736
rect 5040 292318 5100 293666
rect 5236 293630 5418 293664
rect 5162 293580 5174 293592
rect 5220 293580 5222 293591
rect 5421 293580 5434 293591
rect 5480 293580 5492 293592
rect 5162 292404 5222 293580
rect 5432 292404 5492 293580
rect 5162 292392 5174 292404
rect 5480 292392 5492 292404
rect 5236 292320 5418 292354
rect 5554 292318 5614 293666
rect 5040 292248 5088 292318
rect 5566 292248 5614 292318
rect 5040 290900 5100 292248
rect 5236 292212 5418 292246
rect 5162 292162 5174 292174
rect 5220 292162 5222 292173
rect 5421 292162 5434 292173
rect 5480 292162 5492 292174
rect 5162 290986 5222 292162
rect 5432 290986 5492 292162
rect 5162 290974 5174 290986
rect 5480 290974 5492 290986
rect 5236 290902 5418 290936
rect 5554 290900 5614 292248
rect 5040 290830 5088 290900
rect 5566 290830 5614 290900
rect 5040 289482 5100 290830
rect 5236 290794 5418 290828
rect 5162 290744 5174 290756
rect 5220 290744 5222 290755
rect 5421 290744 5434 290755
rect 5480 290744 5492 290756
rect 5162 289568 5222 290744
rect 5432 289568 5492 290744
rect 5162 289556 5174 289568
rect 5480 289556 5492 289568
rect 5236 289484 5418 289518
rect 5554 289482 5614 290830
rect 5040 289412 5088 289482
rect 5566 289412 5614 289482
rect 5040 288064 5100 289412
rect 5236 289376 5418 289410
rect 5162 289326 5174 289338
rect 5220 289326 5222 289337
rect 5421 289326 5434 289337
rect 5480 289326 5492 289338
rect 5162 288150 5222 289326
rect 5432 288150 5492 289326
rect 5162 288138 5174 288150
rect 5480 288138 5492 288150
rect 5236 288066 5418 288100
rect 5554 288064 5614 289412
rect 5040 287994 5088 288064
rect 5566 287994 5614 288064
rect 5040 286646 5100 287994
rect 5236 287958 5418 287992
rect 5162 287908 5174 287920
rect 5220 287908 5222 287919
rect 5421 287908 5434 287919
rect 5480 287908 5492 287920
rect 5162 286732 5222 287908
rect 5432 286732 5492 287908
rect 5162 286720 5174 286732
rect 5480 286720 5492 286732
rect 5236 286648 5418 286682
rect 5554 286646 5614 287994
rect 5040 286576 5088 286646
rect 5566 286576 5614 286646
rect 5040 285228 5100 286576
rect 5236 286540 5418 286574
rect 5162 286490 5174 286502
rect 5220 286490 5222 286501
rect 5421 286490 5434 286501
rect 5480 286490 5492 286502
rect 5162 285314 5222 286490
rect 5432 285314 5492 286490
rect 5162 285302 5174 285314
rect 5480 285302 5492 285314
rect 5236 285230 5418 285264
rect 5554 285228 5614 286576
rect 5040 285158 5088 285228
rect 5566 285158 5614 285228
rect 5040 283810 5100 285158
rect 5236 285122 5418 285156
rect 5162 285072 5174 285084
rect 5220 285072 5222 285083
rect 5421 285072 5434 285083
rect 5480 285072 5492 285084
rect 5162 283896 5222 285072
rect 5432 283896 5492 285072
rect 5162 283884 5174 283896
rect 5480 283884 5492 283896
rect 5236 283812 5418 283846
rect 5554 283810 5614 285158
rect 5040 283740 5088 283810
rect 5566 283740 5614 283810
rect 5040 282392 5100 283740
rect 5236 283704 5418 283738
rect 5162 283654 5174 283666
rect 5220 283654 5222 283665
rect 5421 283654 5434 283665
rect 5480 283654 5492 283666
rect 5162 282478 5222 283654
rect 5432 282478 5492 283654
rect 5162 282466 5174 282478
rect 5480 282466 5492 282478
rect 5236 282394 5418 282428
rect 5554 282392 5614 283740
rect 5040 282322 5088 282392
rect 5566 282322 5614 282392
rect 5040 280974 5100 282322
rect 5236 282286 5418 282320
rect 5162 282236 5174 282248
rect 5220 282236 5222 282247
rect 5421 282236 5434 282247
rect 5480 282236 5492 282248
rect 5162 281060 5222 282236
rect 5432 281060 5492 282236
rect 5162 281048 5174 281060
rect 5480 281048 5492 281060
rect 5236 280976 5418 281010
rect 5554 280974 5614 282322
rect 5040 280904 5088 280974
rect 5566 280904 5614 280974
rect 5040 279556 5100 280904
rect 5236 280868 5418 280902
rect 5162 280818 5174 280830
rect 5220 280818 5222 280829
rect 5421 280818 5434 280829
rect 5480 280818 5492 280830
rect 5162 279642 5222 280818
rect 5432 279642 5492 280818
rect 5162 279630 5174 279642
rect 5480 279630 5492 279642
rect 5236 279558 5418 279592
rect 5554 279556 5614 280904
rect 5040 279486 5088 279556
rect 5566 279486 5614 279556
rect 5040 278138 5100 279486
rect 5236 279450 5418 279484
rect 5162 279400 5174 279412
rect 5220 279400 5222 279411
rect 5421 279400 5434 279411
rect 5480 279400 5492 279412
rect 5162 278224 5222 279400
rect 5432 278224 5492 279400
rect 5162 278212 5174 278224
rect 5480 278212 5492 278224
rect 5236 278140 5418 278174
rect 5554 278138 5614 279486
rect 5040 278068 5088 278138
rect 5566 278068 5614 278138
rect 5040 276720 5100 278068
rect 5236 278032 5418 278066
rect 5162 277982 5174 277994
rect 5220 277982 5222 277993
rect 5421 277982 5434 277993
rect 5480 277982 5492 277994
rect 5162 276806 5222 277982
rect 5432 276806 5492 277982
rect 5162 276794 5174 276806
rect 5480 276794 5492 276806
rect 5236 276722 5418 276756
rect 5554 276720 5614 278068
rect 5040 276650 5088 276720
rect 5566 276650 5614 276720
rect 5040 275302 5100 276650
rect 5236 276614 5418 276648
rect 5162 276564 5174 276576
rect 5220 276564 5222 276575
rect 5421 276564 5434 276575
rect 5480 276564 5492 276576
rect 5162 275388 5222 276564
rect 5432 275388 5492 276564
rect 5162 275376 5174 275388
rect 5480 275376 5492 275388
rect 5236 275304 5418 275338
rect 5554 275302 5614 276650
rect 5040 275232 5088 275302
rect 5566 275232 5614 275302
rect 5040 273884 5100 275232
rect 5236 275196 5418 275230
rect 5162 275146 5174 275158
rect 5220 275146 5222 275157
rect 5421 275146 5434 275157
rect 5480 275146 5492 275158
rect 5162 273970 5222 275146
rect 5432 273970 5492 275146
rect 5162 273958 5174 273970
rect 5480 273958 5492 273970
rect 5236 273886 5418 273920
rect 5554 273884 5614 275232
rect 5040 273814 5088 273884
rect 5566 273814 5614 273884
rect 5040 272466 5100 273814
rect 5236 273778 5418 273812
rect 5162 273728 5174 273740
rect 5220 273728 5222 273739
rect 5421 273728 5434 273739
rect 5480 273728 5492 273740
rect 5162 272552 5222 273728
rect 5432 272552 5492 273728
rect 5162 272540 5174 272552
rect 5480 272540 5492 272552
rect 5236 272468 5418 272502
rect 5554 272466 5614 273814
rect 5040 272396 5088 272466
rect 5566 272396 5614 272466
rect 5040 271048 5100 272396
rect 5236 272360 5418 272394
rect 5162 272310 5174 272322
rect 5220 272310 5222 272321
rect 5421 272310 5434 272321
rect 5480 272310 5492 272322
rect 5162 271134 5222 272310
rect 5432 271134 5492 272310
rect 5162 271122 5174 271134
rect 5480 271122 5492 271134
rect 5236 271050 5418 271084
rect 5554 271048 5614 272396
rect 5040 270978 5088 271048
rect 5566 270978 5614 271048
rect 5040 269630 5100 270978
rect 5236 270942 5418 270976
rect 5162 270892 5174 270904
rect 5220 270892 5222 270903
rect 5421 270892 5434 270903
rect 5480 270892 5492 270904
rect 5162 269716 5222 270892
rect 5432 269716 5492 270892
rect 5162 269704 5174 269716
rect 5480 269704 5492 269716
rect 5236 269632 5418 269666
rect 5554 269630 5614 270978
rect 5040 269560 5088 269630
rect 5566 269560 5614 269630
rect 5040 268212 5100 269560
rect 5236 269524 5418 269558
rect 5162 269474 5174 269486
rect 5220 269474 5222 269485
rect 5421 269474 5434 269485
rect 5480 269474 5492 269486
rect 5162 268298 5222 269474
rect 5432 268298 5492 269474
rect 5162 268286 5174 268298
rect 5480 268286 5492 268298
rect 5236 268214 5418 268248
rect 5554 268212 5614 269560
rect 5040 268142 5088 268212
rect 5566 268142 5614 268212
rect 5040 266794 5100 268142
rect 5236 268106 5418 268140
rect 5162 268056 5174 268068
rect 5220 268056 5222 268067
rect 5421 268056 5434 268067
rect 5480 268056 5492 268068
rect 5162 266880 5222 268056
rect 5432 266880 5492 268056
rect 5162 266868 5174 266880
rect 5480 266868 5492 266880
rect 5236 266796 5418 266830
rect 5554 266794 5614 268142
rect 5040 266724 5088 266794
rect 5566 266724 5614 266794
rect 5040 265376 5100 266724
rect 5236 266688 5418 266722
rect 5162 266638 5174 266650
rect 5220 266638 5222 266649
rect 5421 266638 5434 266649
rect 5480 266638 5492 266650
rect 5162 265462 5222 266638
rect 5432 265462 5492 266638
rect 5162 265450 5174 265462
rect 5480 265450 5492 265462
rect 5236 265378 5418 265412
rect 5554 265376 5614 266724
rect 5040 265306 5088 265376
rect 5566 265306 5614 265376
rect 5040 263958 5100 265306
rect 5236 265270 5418 265304
rect 5162 265220 5174 265232
rect 5220 265220 5222 265231
rect 5421 265220 5434 265231
rect 5480 265220 5492 265232
rect 5162 264044 5222 265220
rect 5432 264044 5492 265220
rect 5162 264032 5174 264044
rect 5480 264032 5492 264044
rect 5236 263960 5418 263994
rect 5554 263958 5614 265306
rect 5040 263888 5088 263958
rect 5566 263888 5614 263958
rect 5040 262540 5100 263888
rect 5236 263852 5418 263886
rect 5162 263802 5174 263814
rect 5220 263802 5222 263813
rect 5421 263802 5434 263813
rect 5480 263802 5492 263814
rect 5162 262626 5222 263802
rect 5432 262626 5492 263802
rect 5162 262614 5174 262626
rect 5480 262614 5492 262626
rect 5236 262542 5418 262576
rect 5554 262540 5614 263888
rect 5040 262470 5088 262540
rect 5566 262470 5614 262540
rect 5040 261122 5100 262470
rect 5236 262434 5418 262468
rect 5162 262384 5174 262396
rect 5220 262384 5222 262395
rect 5421 262384 5434 262395
rect 5480 262384 5492 262396
rect 5162 261208 5222 262384
rect 5432 261208 5492 262384
rect 5162 261196 5174 261208
rect 5480 261196 5492 261208
rect 5236 261124 5418 261158
rect 5554 261122 5614 262470
rect 5040 261052 5088 261122
rect 5566 261052 5614 261122
rect 5040 259704 5100 261052
rect 5236 261016 5418 261050
rect 5162 260966 5174 260978
rect 5220 260966 5222 260977
rect 5421 260966 5434 260977
rect 5480 260966 5492 260978
rect 5162 259790 5222 260966
rect 5432 259790 5492 260966
rect 5162 259778 5174 259790
rect 5480 259778 5492 259790
rect 5236 259706 5418 259740
rect 5554 259704 5614 261052
rect 5040 259634 5088 259704
rect 5566 259634 5614 259704
rect 5040 258286 5100 259634
rect 5236 259598 5418 259632
rect 5162 259548 5174 259560
rect 5220 259548 5222 259559
rect 5421 259548 5434 259559
rect 5480 259548 5492 259560
rect 5162 258372 5222 259548
rect 5432 258372 5492 259548
rect 5162 258360 5174 258372
rect 5480 258360 5492 258372
rect 5236 258288 5418 258322
rect 5554 258286 5614 259634
rect 5040 258216 5088 258286
rect 5566 258216 5614 258286
rect 5040 256868 5100 258216
rect 5236 258180 5418 258214
rect 5162 258130 5174 258142
rect 5220 258130 5222 258141
rect 5421 258130 5434 258141
rect 5480 258130 5492 258142
rect 5162 256954 5222 258130
rect 5432 256954 5492 258130
rect 5162 256942 5174 256954
rect 5480 256942 5492 256954
rect 5236 256870 5418 256904
rect 5554 256868 5614 258216
rect 5040 256798 5088 256868
rect 5566 256798 5614 256868
rect 5040 255450 5100 256798
rect 5236 256762 5418 256796
rect 5162 256712 5174 256724
rect 5220 256712 5222 256723
rect 5421 256712 5434 256723
rect 5480 256712 5492 256724
rect 5162 255536 5222 256712
rect 5432 255536 5492 256712
rect 5162 255524 5174 255536
rect 5480 255524 5492 255536
rect 5236 255452 5418 255486
rect 5554 255450 5614 256798
rect 5040 255380 5088 255450
rect 5566 255380 5614 255450
rect 5040 254231 5100 255380
rect 5236 255344 5418 255378
rect 5162 255294 5174 255306
rect 5220 255294 5222 255305
rect 5421 255294 5434 255305
rect 5480 255294 5492 255306
rect 5162 254231 5222 255294
rect 3794 254136 5222 254231
rect 5432 254136 5492 255294
rect 5554 254136 5614 255380
rect 3794 254012 5662 254136
rect 3464 253287 3646 253321
rect 3464 253179 3646 253213
rect 3448 253120 3450 253131
rect 3649 253120 3662 253131
rect 3402 251944 3450 253120
rect 3660 251944 3708 253120
rect 3464 251851 3646 251885
rect 3464 251743 3646 251777
rect 3448 251684 3450 251695
rect 3649 251684 3662 251695
rect 3402 250508 3450 251684
rect 3660 250508 3708 251684
rect 3464 250415 3646 250449
rect 3464 250307 3646 250341
rect 3448 250248 3450 250259
rect 3649 250248 3662 250259
rect 3402 249072 3450 250248
rect 3660 249072 3708 250248
rect 3464 248979 3646 249013
rect 3464 248871 3646 248905
rect 3448 248812 3450 248823
rect 3649 248812 3662 248823
rect 3402 247636 3450 248812
rect 3660 247636 3708 248812
rect 3464 247543 3646 247577
rect 3464 247435 3646 247469
rect 3448 247376 3450 247387
rect 3649 247376 3662 247387
rect 3402 246200 3450 247376
rect 3660 246200 3708 247376
rect 3464 246107 3646 246141
rect 3464 245999 3646 246033
rect 3448 245940 3450 245951
rect 3649 245940 3662 245951
rect 3402 244764 3450 245940
rect 3660 244764 3708 245940
rect 3464 244671 3646 244705
rect 3464 244563 3646 244597
rect 3448 244504 3450 244515
rect 3649 244504 3662 244515
rect 3402 243328 3450 244504
rect 3660 243328 3708 244504
rect 3464 243235 3646 243269
rect 3464 243127 3646 243161
rect 3448 243068 3450 243079
rect 3649 243068 3662 243079
rect 3402 241892 3450 243068
rect 3660 241892 3708 243068
rect 3464 241799 3646 241833
rect 3464 241691 3646 241725
rect 3448 241632 3450 241643
rect 3649 241632 3662 241643
rect 3402 240456 3450 241632
rect 3660 240456 3708 241632
rect 3464 240363 3646 240397
rect 3464 240255 3646 240289
rect 3448 240196 3450 240207
rect 3649 240196 3662 240207
rect 3402 239020 3450 240196
rect 3660 239020 3708 240196
rect 3464 238927 3646 238961
rect 3464 238819 3646 238853
rect 3448 238760 3450 238771
rect 3649 238760 3662 238771
rect 3402 237584 3450 238760
rect 3660 237584 3708 238760
rect 3464 237491 3646 237525
rect 3464 237383 3646 237417
rect 3448 237324 3450 237335
rect 3649 237324 3662 237335
rect 3402 236148 3450 237324
rect 3660 236148 3708 237324
rect 3464 236055 3646 236089
rect 3464 235947 3646 235981
rect 3448 235888 3450 235899
rect 3649 235888 3662 235899
rect 3402 234712 3450 235888
rect 3660 234712 3708 235888
rect 3464 234619 3646 234653
rect 3464 234511 3646 234545
rect 3448 234452 3450 234463
rect 3649 234452 3662 234463
rect 3402 233276 3450 234452
rect 3660 233276 3708 234452
rect 3464 233183 3646 233217
rect 3464 233075 3646 233109
rect 3448 233016 3450 233027
rect 3649 233016 3662 233027
rect 3402 231840 3450 233016
rect 3660 231840 3708 233016
rect 3464 231747 3646 231781
rect 3464 231639 3646 231673
rect 3448 231580 3450 231591
rect 3649 231580 3662 231591
rect 3402 230404 3450 231580
rect 3660 230404 3708 231580
rect 3464 230311 3646 230345
rect 3464 230203 3646 230237
rect 3448 230144 3450 230155
rect 3649 230144 3662 230155
rect 3402 228968 3450 230144
rect 3660 228968 3708 230144
rect 3464 228875 3646 228909
rect 3464 228767 3646 228801
rect 3448 228708 3450 228719
rect 3649 228708 3662 228719
rect 3402 227532 3450 228708
rect 3660 227532 3708 228708
rect 3464 227439 3646 227473
rect 3464 227331 3646 227365
rect 3448 227272 3450 227283
rect 3649 227272 3662 227283
rect 3402 226096 3450 227272
rect 3660 226096 3708 227272
rect 3464 226003 3646 226037
rect 3464 225895 3646 225929
rect 3448 225836 3450 225847
rect 3649 225836 3662 225847
rect 3402 224660 3450 225836
rect 3660 224660 3708 225836
rect 3464 224567 3646 224601
rect 3464 224459 3646 224493
rect 3448 224400 3450 224411
rect 3649 224400 3662 224411
rect 3402 223224 3450 224400
rect 3660 223224 3708 224400
rect 3464 223131 3646 223165
rect 3464 223023 3646 223057
rect 3448 222964 3450 222975
rect 3649 222964 3662 222975
rect 3402 221788 3450 222964
rect 3660 221788 3708 222964
rect 3464 221695 3646 221729
rect 3464 221587 3646 221621
rect 3448 221528 3450 221539
rect 3649 221528 3662 221539
rect 3402 220352 3450 221528
rect 3660 220352 3708 221528
rect 3464 220259 3646 220293
rect 3464 220151 3646 220185
rect 3448 220092 3450 220103
rect 3649 220092 3662 220103
rect 3402 218916 3450 220092
rect 3660 218916 3708 220092
rect 3464 218823 3646 218857
rect 3464 218715 3646 218749
rect 3448 218656 3450 218667
rect 3649 218656 3662 218667
rect 3402 217480 3450 218656
rect 3660 217480 3708 218656
rect 3464 217387 3646 217421
rect 3464 217279 3646 217313
rect 3448 217220 3450 217231
rect 3649 217220 3662 217231
rect 3402 216044 3450 217220
rect 3660 216044 3708 217220
rect 3464 215951 3646 215985
rect 3464 215843 3646 215877
rect 3448 215784 3450 215795
rect 3649 215784 3662 215795
rect 3402 214608 3450 215784
rect 3660 214608 3708 215784
rect 3464 214515 3646 214549
rect 3464 214407 3646 214441
rect 3448 214348 3450 214359
rect 3649 214348 3662 214359
rect 3402 213172 3450 214348
rect 3660 213172 3708 214348
rect 3464 213079 3646 213113
rect 3464 212971 3646 213005
rect 3448 212912 3450 212923
rect 3649 212912 3662 212923
rect 3402 211736 3450 212912
rect 3660 211736 3708 212912
rect 3464 211643 3646 211677
rect 3464 211535 3646 211569
rect 3448 211476 3450 211487
rect 3649 211476 3662 211487
rect 3402 210300 3450 211476
rect 3660 210300 3708 211476
rect 3464 210207 3646 210241
rect 3464 210099 3646 210133
rect 3448 210040 3450 210051
rect 3649 210040 3662 210051
rect 3402 208864 3450 210040
rect 3660 208864 3708 210040
rect 3464 208771 3646 208805
rect 3464 208663 3646 208697
rect 3448 208604 3450 208615
rect 3649 208604 3662 208615
rect 3402 207428 3450 208604
rect 3660 207428 3708 208604
rect 3464 207335 3646 207369
rect 3464 207227 3646 207261
rect 3448 207168 3450 207179
rect 3649 207168 3662 207179
rect 3402 205992 3450 207168
rect 3660 205992 3708 207168
rect 3464 205899 3646 205933
rect 3464 205791 3646 205825
rect 3448 205732 3450 205743
rect 3649 205732 3662 205743
rect 3402 204556 3450 205732
rect 3660 204556 3708 205732
rect 3464 204463 3646 204497
rect 3464 204355 3646 204389
rect 3448 204296 3450 204307
rect 3649 204296 3662 204307
rect 3402 203120 3450 204296
rect 3660 203120 3708 204296
rect 3464 203027 3646 203061
rect 3464 202919 3646 202953
rect 3448 202860 3450 202871
rect 3649 202860 3662 202871
rect 3402 201684 3450 202860
rect 3660 201684 3708 202860
rect 3464 201591 3646 201625
rect 3464 201483 3646 201517
rect 3448 201424 3450 201435
rect 3649 201424 3662 201435
rect 3402 200248 3450 201424
rect 3660 200248 3708 201424
rect 3464 200155 3646 200189
rect 3464 200047 3646 200081
rect 3448 199988 3450 199999
rect 3649 199988 3662 199999
rect 3402 198812 3450 199988
rect 3660 198812 3708 199988
rect 3464 198719 3646 198753
rect 3464 198611 3646 198645
rect 3794 198583 5717 254012
rect -10 -4475 24 -2475
rect 112 -4379 428 -4367
rect 516 -4379 550 -2475
rect 3219 -4079 5717 198583
rect 3190 -4127 5717 -4079
rect 1267 -4161 5717 -4127
rect 112 -4413 670 -4379
rect 112 -4425 428 -4413
rect -12 -5121 24 -4475
rect 124 -4483 158 -4425
rect 124 -4585 164 -4483
rect 382 -4501 428 -4470
rect 516 -4479 550 -4413
rect 516 -4490 554 -4479
rect 168 -4517 170 -4501
rect 172 -4517 192 -4511
rect 370 -4517 428 -4501
rect 168 -4551 428 -4517
rect 124 -4610 158 -4585
rect 122 -4986 158 -4610
rect 168 -4598 170 -4551
rect 172 -4557 192 -4551
rect 370 -4598 428 -4551
rect 504 -4501 515 -4490
rect 516 -4501 562 -4490
rect 122 -5121 156 -4986
rect 162 -4998 164 -4972
rect 168 -4986 169 -4598
rect 382 -4986 416 -4598
rect 504 -4814 562 -4501
rect 1123 -4796 2826 -4301
rect 3190 -4394 5717 -4161
rect 3190 -4488 5783 -4394
rect 3190 -4796 5835 -4488
rect 1123 -4814 5835 -4796
rect 162 -5026 192 -5000
rect 354 -5045 401 -4998
rect 170 -5079 401 -5045
rect -12 -5129 22 -5121
rect 93 -5129 156 -5121
rect 504 -5129 5835 -4814
rect 6433 -4954 6578 -4943
rect 6433 -4988 6541 -4954
rect 6433 -5000 6578 -4988
rect 6433 -5059 6491 -5000
rect -26 -5215 5835 -5129
rect -12 -5223 22 -5215
rect 88 -5217 5835 -5215
rect 110 -5223 5835 -5217
rect -12 -5228 5835 -5223
rect -12 -5349 22 -5228
rect 110 -5229 5835 -5228
rect 317 -5251 5835 -5229
rect 325 -5257 5835 -5251
rect 323 -5291 5835 -5257
rect 325 -5349 5835 -5291
rect -59 -6032 5835 -5349
rect 5842 -6032 5889 -5095
rect -59 -6465 6027 -6032
rect 515 -6478 6027 -6465
rect 532 -6495 6027 -6478
rect 595 -6528 598 -6495
rect 611 -6535 648 -6501
rect 653 -6535 658 -6495
rect 687 -6516 744 -6495
rect 773 -6501 896 -6495
rect 653 -6593 656 -6535
rect 611 -6637 648 -6603
rect 653 -6637 658 -6593
rect 653 -6653 656 -6637
rect 687 -6681 690 -6516
rect 697 -6535 734 -6516
rect 697 -6641 734 -6607
rect 741 -6681 744 -6516
rect 775 -6516 896 -6501
rect 775 -6593 778 -6516
rect 783 -6535 820 -6516
rect 1052 -6519 1089 -6495
rect 1097 -6519 1100 -6495
rect 1159 -6501 1245 -6495
rect 1253 -6501 1256 -6495
rect 1364 -6501 1401 -6495
rect 1409 -6501 1412 -6495
rect 1520 -6501 1557 -6495
rect 1565 -6501 1568 -6495
rect 1676 -6501 1713 -6495
rect 1721 -6501 1724 -6495
rect 1832 -6501 1869 -6495
rect 2219 -6501 2256 -6495
rect 2287 -6501 2324 -6495
rect 2355 -6501 2392 -6495
rect 2423 -6501 2460 -6495
rect 2491 -6501 2528 -6495
rect 2559 -6501 2596 -6495
rect 2627 -6501 2664 -6495
rect 2695 -6501 6027 -6495
rect 1159 -6533 1877 -6501
rect 2199 -6513 6027 -6501
rect 1159 -6547 1903 -6533
rect 1159 -6559 1877 -6547
rect 2160 -6552 6027 -6513
rect 2160 -6559 5835 -6552
rect 773 -6603 778 -6593
rect 1052 -6601 1089 -6567
rect 1097 -6601 1100 -6559
rect 1197 -6567 1200 -6559
rect 1208 -6601 1245 -6567
rect 1253 -6601 1256 -6559
rect 1353 -6567 1356 -6559
rect 1364 -6601 1401 -6567
rect 1409 -6601 1412 -6559
rect 1509 -6567 1512 -6559
rect 1520 -6601 1557 -6567
rect 1565 -6601 1568 -6559
rect 1665 -6567 1668 -6559
rect 1676 -6601 1713 -6567
rect 1721 -6601 1724 -6559
rect 1821 -6567 1824 -6559
rect 2731 -6563 5835 -6559
rect 1832 -6601 1869 -6567
rect 2196 -6581 2317 -6578
rect 2386 -6581 5835 -6563
rect 775 -6653 778 -6603
rect 783 -6637 820 -6603
rect 2246 -6628 2283 -6594
rect 2291 -6628 2294 -6586
rect 2391 -6594 2394 -6586
rect 2402 -6628 2439 -6594
rect 2447 -6628 2450 -6586
rect 2703 -6594 2706 -6586
rect 2731 -6590 5835 -6581
rect 1052 -6681 1089 -6647
rect 1097 -6681 1100 -6636
rect 1197 -6647 1200 -6636
rect 1208 -6681 1245 -6647
rect 1253 -6681 1256 -6636
rect 1353 -6647 1356 -6636
rect 1364 -6681 1401 -6647
rect 1409 -6681 1412 -6636
rect 1509 -6647 1512 -6636
rect 1520 -6681 1557 -6647
rect 1565 -6681 1568 -6636
rect 1665 -6647 1668 -6636
rect 1676 -6681 1713 -6647
rect 1721 -6681 1724 -6636
rect 1821 -6647 1824 -6636
rect 1832 -6681 1869 -6647
rect 625 -6727 662 -6693
rect 697 -6715 734 -6681
rect 769 -6727 806 -6693
rect 1016 -6715 1053 -6681
rect 1088 -6715 1125 -6681
rect 1328 -6715 1365 -6681
rect 1400 -6715 1437 -6681
rect 1640 -6715 1677 -6681
rect 1712 -6715 1749 -6681
rect 2246 -6728 2283 -6694
rect 2291 -6728 2294 -6683
rect 2391 -6694 2394 -6683
rect 2438 -6694 2439 -6628
rect 2402 -6728 2439 -6694
rect 2447 -6728 2450 -6683
rect 2202 -6764 2239 -6730
rect 2274 -6764 2311 -6730
rect 2438 -6744 2439 -6728
rect 2472 -6764 2473 -6633
rect 2547 -6664 2550 -6653
rect 2558 -6698 2595 -6664
rect 2603 -6698 2606 -6653
rect 2478 -6764 2515 -6730
rect 2550 -6764 2587 -6730
rect 2622 -6764 2659 -6730
rect 2664 -6764 2665 -6633
rect 2698 -6744 2699 -6599
rect 2714 -6628 2751 -6594
rect 2759 -6628 2762 -6590
rect 2859 -6594 2919 -6590
rect 2862 -6633 2919 -6594
rect 3099 -6647 3136 -6613
rect 3144 -6647 3147 -6602
rect 2703 -6694 2706 -6683
rect 2714 -6728 2751 -6694
rect 2759 -6728 2762 -6683
rect 2859 -6694 2862 -6683
rect 2870 -6728 2907 -6694
rect 3099 -6715 3136 -6681
rect 3144 -6715 3147 -6670
rect 2860 -6764 2897 -6730
rect 3190 -6776 5835 -6590
rect 31 -6817 68 -6783
rect 127 -6817 164 -6783
rect 223 -6817 260 -6783
rect 319 -6817 356 -6783
rect 415 -6817 452 -6783
rect 511 -6817 548 -6783
rect 607 -6817 644 -6783
rect 703 -6817 740 -6783
rect 799 -6817 836 -6783
rect 895 -6817 932 -6783
rect 991 -6817 1028 -6783
rect 1087 -6817 1124 -6783
rect 1183 -6817 1220 -6783
rect 1279 -6817 1316 -6783
rect 1375 -6817 1412 -6783
rect 1471 -6817 1508 -6783
rect 1567 -6817 1604 -6783
rect 1663 -6817 1700 -6783
rect 1759 -6817 1796 -6783
rect 1855 -6817 1892 -6783
rect 1951 -6817 1988 -6783
rect 2047 -6817 2084 -6783
rect 3031 -6810 3068 -6776
rect 3103 -6810 3140 -6776
rect 3175 -6810 5835 -6776
rect 3190 -6816 5835 -6810
rect 3190 -6819 5783 -6816
rect 5788 -6819 5835 -6816
rect 5842 -6638 5888 -6552
rect 5842 -6724 5900 -6638
rect 5906 -6650 5922 -6552
rect 5976 -6717 5988 -6578
rect 5842 -6758 5920 -6724
rect 5842 -6788 5900 -6758
rect 5842 -6814 5873 -6788
rect 5842 -6819 5889 -6814
rect 2209 -6860 2246 -6826
rect 2305 -6860 2342 -6826
rect 2401 -6860 2438 -6826
rect 2497 -6860 2534 -6826
rect 2593 -6860 2630 -6826
rect 2689 -6860 2726 -6826
rect 2785 -6860 2822 -6826
rect 2881 -6860 2918 -6826
rect 3190 -6853 5889 -6819
rect 5905 -6853 5942 -6819
rect 3190 -6858 5783 -6853
rect 5788 -6858 5835 -6853
rect 3043 -6903 3080 -6869
rect 3139 -6903 3176 -6869
rect 3190 -6874 5835 -6858
rect 3190 -6912 5783 -6874
rect 5842 -6912 5889 -6853
rect 3190 -6928 5889 -6912
rect 3190 -6929 5783 -6928
rect 3219 -6972 5783 -6929
rect 5797 -6946 5834 -6928
rect 5893 -6946 5930 -6912
rect 5950 -6927 5964 -6893
rect 6367 -6939 6491 -5059
rect 6567 -6773 6578 -5173
rect 39 -7603 87 -7569
rect 135 -7603 183 -7569
rect 231 -7603 279 -7569
rect 327 -7603 375 -7569
rect 423 -7603 471 -7569
rect 500 -7603 502 -7569
rect 554 -7646 556 -7612
rect 585 -7646 633 -7612
rect 681 -7646 729 -7612
rect 777 -7646 825 -7612
rect 873 -7646 921 -7612
rect 969 -7646 1017 -7612
rect 1065 -7646 1113 -7612
rect 1161 -7646 1209 -7612
rect 1238 -7646 1240 -7612
rect 141 -7665 155 -7657
rect 218 -7665 230 -7649
rect 252 -7657 264 -7649
rect 306 -7657 316 -7649
rect 241 -7665 264 -7657
rect 297 -7665 316 -7657
rect 32 -7699 80 -7665
rect 96 -7699 155 -7665
rect 176 -7699 230 -7665
rect 141 -7748 155 -7737
rect 96 -7782 155 -7748
rect 141 -7832 155 -7821
rect 96 -7866 155 -7832
rect 141 -7915 155 -7904
rect 96 -7949 155 -7915
rect 218 -7965 230 -7699
rect 252 -7699 316 -7665
rect 252 -7737 264 -7699
rect 306 -7737 316 -7699
rect 241 -7748 264 -7737
rect 297 -7748 316 -7737
rect 252 -7782 316 -7748
rect 252 -7821 264 -7782
rect 306 -7821 316 -7782
rect 241 -7832 264 -7821
rect 297 -7832 316 -7821
rect 252 -7866 316 -7832
rect 252 -7904 264 -7866
rect 306 -7904 316 -7866
rect 241 -7915 264 -7904
rect 297 -7915 316 -7904
rect 252 -7949 316 -7915
rect 241 -7983 264 -7949
rect 252 -7999 264 -7983
rect 161 -8063 209 -8029
rect 218 -8090 225 -8013
rect 252 -8095 259 -7999
rect 283 -8131 297 -7983
rect 306 -7999 316 -7949
rect 340 -7665 350 -7649
rect 397 -7665 411 -7657
rect 340 -7699 394 -7665
rect 408 -7699 466 -7665
rect 1292 -7689 1294 -7655
rect 1323 -7689 1371 -7655
rect 1419 -7689 1467 -7655
rect 1515 -7689 1563 -7655
rect 1592 -7689 1594 -7655
rect 340 -7965 350 -7699
rect 1116 -7708 1128 -7692
rect 1150 -7700 1162 -7692
rect 1139 -7708 1162 -7700
rect 397 -7748 411 -7737
rect 576 -7742 624 -7708
rect 648 -7742 696 -7708
rect 720 -7742 768 -7708
rect 864 -7742 912 -7708
rect 936 -7742 1056 -7708
rect 1080 -7742 1128 -7708
rect 408 -7782 456 -7748
rect 397 -7832 411 -7821
rect 973 -7825 1021 -7791
rect 408 -7866 456 -7832
rect 397 -7915 411 -7904
rect 408 -7949 456 -7915
rect 683 -7941 697 -7930
rect 638 -7975 697 -7941
rect 760 -7992 772 -7874
rect 794 -7930 806 -7908
rect 783 -7941 806 -7930
rect 830 -7941 842 -7908
rect 794 -7975 842 -7941
rect 794 -8026 806 -7975
rect 830 -8026 842 -7975
rect 864 -7992 876 -7875
rect 961 -7916 968 -7875
rect 973 -7909 1021 -7875
rect 973 -7992 1021 -7958
rect 1116 -7992 1128 -7742
rect 1150 -7742 1198 -7708
rect 1646 -7732 1648 -7698
rect 1677 -7732 1725 -7698
rect 1773 -7732 1821 -7698
rect 1869 -7732 1917 -7698
rect 1946 -7732 1948 -7698
rect 1150 -7780 1162 -7742
rect 1389 -7751 1403 -7743
rect 1489 -7751 1503 -7743
rect 1139 -7791 1162 -7780
rect 1316 -7785 1436 -7751
rect 1500 -7785 1548 -7751
rect 2000 -7775 2002 -7741
rect 2031 -7775 2079 -7741
rect 2127 -7775 2175 -7741
rect 2223 -7775 2271 -7741
rect 2319 -7775 2367 -7741
rect 2415 -7775 2463 -7741
rect 2492 -7775 2494 -7741
rect 3219 -7784 5717 -6972
rect 6367 -6975 6480 -6939
rect 6433 -6993 6480 -6975
rect 1150 -7825 1198 -7791
rect 1743 -7794 1757 -7786
rect 1843 -7794 1857 -7786
rect 1150 -7864 1162 -7825
rect 1389 -7834 1403 -7823
rect 1489 -7834 1503 -7823
rect 1670 -7828 1790 -7794
rect 1854 -7828 1902 -7794
rect 2546 -7818 2548 -7784
rect 2577 -7818 2625 -7784
rect 2673 -7818 2721 -7784
rect 2769 -7818 2817 -7784
rect 2865 -7818 2913 -7784
rect 2961 -7818 3009 -7784
rect 3057 -7818 3105 -7784
rect 3153 -7818 5717 -7784
rect 1139 -7875 1162 -7864
rect 1344 -7868 1403 -7834
rect 1500 -7868 1548 -7834
rect 2133 -7837 2147 -7829
rect 2210 -7837 2222 -7821
rect 2244 -7829 2256 -7821
rect 2298 -7829 2308 -7821
rect 2233 -7837 2256 -7829
rect 2289 -7837 2308 -7829
rect 1150 -7909 1198 -7875
rect 1743 -7877 1757 -7866
rect 1843 -7877 1857 -7866
rect 2024 -7871 2072 -7837
rect 2088 -7871 2147 -7837
rect 2168 -7871 2222 -7837
rect 1150 -7947 1162 -7909
rect 1389 -7918 1403 -7907
rect 1489 -7918 1503 -7907
rect 1698 -7911 1757 -7877
rect 1854 -7911 1902 -7877
rect 1139 -7958 1162 -7947
rect 1344 -7952 1403 -7918
rect 1500 -7952 1548 -7918
rect 2133 -7920 2147 -7909
rect 1150 -7992 1198 -7958
rect 1743 -7961 1757 -7950
rect 1843 -7961 1857 -7950
rect 2088 -7954 2147 -7920
rect 1150 -8026 1162 -7992
rect 1389 -8001 1403 -7990
rect 1489 -8001 1503 -7990
rect 1698 -7995 1757 -7961
rect 1854 -7995 1902 -7961
rect 403 -8045 415 -8029
rect 141 -8147 155 -8139
rect 96 -8181 155 -8147
rect 283 -8199 302 -8131
rect 324 -8165 336 -8097
rect 369 -8129 381 -8061
rect 403 -8079 461 -8045
rect 403 -8095 415 -8079
rect 614 -8124 662 -8090
rect 383 -8147 397 -8139
rect 394 -8181 442 -8147
rect 614 -8192 662 -8158
rect 141 -8247 155 -8236
rect 96 -8281 155 -8247
rect 283 -8287 297 -8199
rect 663 -8208 675 -8074
rect 383 -8247 397 -8236
rect 697 -8242 709 -8048
rect 737 -8064 751 -8053
rect 733 -8095 751 -8064
rect 1059 -8082 1107 -8048
rect 394 -8281 442 -8247
rect 637 -8277 651 -8266
rect 32 -8321 80 -8287
rect 104 -8321 152 -8287
rect 176 -8321 224 -8287
rect 248 -8315 297 -8287
rect 592 -8311 651 -8277
rect 733 -8278 745 -8095
rect 779 -8098 793 -8095
rect 1116 -8098 1123 -8028
rect 767 -8281 793 -8098
rect 795 -8146 843 -8112
rect 1150 -8132 1157 -8026
rect 1344 -8035 1403 -8001
rect 1500 -8035 1548 -8001
rect 2133 -8004 2147 -7993
rect 1743 -8044 1757 -8033
rect 1843 -8044 1857 -8033
rect 2088 -8038 2147 -8004
rect 795 -8214 843 -8180
rect 847 -8281 859 -8146
rect 1409 -8149 1457 -8115
rect 1461 -8176 1473 -8099
rect 881 -8266 893 -8178
rect 1043 -8194 1057 -8186
rect 998 -8228 1057 -8194
rect 1143 -8198 1157 -8187
rect 1154 -8232 1202 -8198
rect 1495 -8210 1507 -8065
rect 1698 -8078 1757 -8044
rect 1854 -8078 1902 -8044
rect 2133 -8087 2147 -8076
rect 1763 -8192 1811 -8158
rect 1815 -8219 1827 -8142
rect 1393 -8237 1407 -8229
rect 1493 -8237 1507 -8229
rect 879 -8277 893 -8266
rect 1348 -8271 1407 -8237
rect 1504 -8271 1552 -8237
rect 1849 -8253 1861 -8108
rect 2088 -8121 2147 -8087
rect 2210 -8137 2222 -7871
rect 2244 -7871 2308 -7837
rect 2244 -7909 2256 -7871
rect 2298 -7909 2308 -7871
rect 2233 -7920 2256 -7909
rect 2289 -7920 2308 -7909
rect 2244 -7954 2308 -7920
rect 2244 -7993 2256 -7954
rect 2298 -7993 2308 -7954
rect 2233 -8004 2256 -7993
rect 2289 -8004 2308 -7993
rect 2244 -8038 2308 -8004
rect 2244 -8076 2256 -8038
rect 2298 -8076 2308 -8038
rect 2233 -8087 2256 -8076
rect 2289 -8087 2308 -8076
rect 2244 -8121 2308 -8087
rect 2233 -8155 2256 -8121
rect 2244 -8171 2256 -8155
rect 2153 -8235 2201 -8201
rect 2210 -8262 2217 -8185
rect 2244 -8267 2251 -8171
rect 248 -8321 296 -8315
rect 779 -8362 793 -8281
rect 881 -8311 938 -8277
rect 1043 -8294 1057 -8283
rect 1143 -8290 1157 -8279
rect 1747 -8280 1761 -8272
rect 1847 -8280 1861 -8272
rect 998 -8328 1057 -8294
rect 1154 -8324 1202 -8290
rect 1702 -8314 1761 -8280
rect 1858 -8314 1906 -8280
rect 2275 -8303 2289 -8155
rect 2298 -8171 2308 -8121
rect 2332 -7837 2342 -7821
rect 2389 -7837 2403 -7829
rect 2332 -7871 2386 -7837
rect 2400 -7871 2458 -7837
rect 2332 -8137 2342 -7871
rect 3108 -7880 3120 -7864
rect 3142 -7872 3154 -7864
rect 3219 -7870 5717 -7818
rect 3131 -7880 3154 -7872
rect 2389 -7920 2403 -7909
rect 2568 -7914 2616 -7880
rect 2640 -7914 2688 -7880
rect 2712 -7914 2760 -7880
rect 2856 -7914 2904 -7880
rect 2928 -7914 3048 -7880
rect 3072 -7914 3120 -7880
rect 2400 -7954 2448 -7920
rect 2389 -8004 2403 -7993
rect 2965 -7997 3013 -7963
rect 2400 -8038 2448 -8004
rect 2389 -8087 2403 -8076
rect 2400 -8121 2448 -8087
rect 2675 -8113 2689 -8102
rect 2630 -8147 2689 -8113
rect 2752 -8164 2764 -8046
rect 2786 -8102 2798 -8080
rect 2775 -8113 2798 -8102
rect 2822 -8113 2834 -8080
rect 2786 -8147 2834 -8113
rect 2786 -8198 2798 -8147
rect 2822 -8198 2834 -8147
rect 2856 -8164 2868 -8047
rect 2953 -8088 2960 -8047
rect 2965 -8081 3013 -8047
rect 2965 -8164 3013 -8130
rect 3108 -8164 3120 -7914
rect 3142 -7914 3190 -7880
rect 3142 -7952 3154 -7914
rect 3131 -7963 3154 -7952
rect 3142 -7997 3190 -7963
rect 3142 -8036 3154 -7997
rect 3131 -8047 3154 -8036
rect 3142 -8081 3190 -8047
rect 3142 -8119 3154 -8081
rect 3131 -8130 3154 -8119
rect 3142 -8164 3190 -8130
rect 3142 -8198 3154 -8164
rect 3201 -8172 3202 -7872
rect 3219 -7904 5735 -7870
rect 5783 -7904 5831 -7870
rect 5879 -7904 5927 -7870
rect 5975 -7904 6023 -7870
rect 6071 -7904 6119 -7870
rect 6167 -7904 6215 -7870
rect 6263 -7904 6311 -7870
rect 6359 -7904 6407 -7870
rect 6455 -7904 6503 -7870
rect 6551 -7904 6599 -7870
rect 6647 -7904 6695 -7870
rect 6743 -7904 6791 -7870
rect 6820 -7904 6822 -7870
rect 3219 -7958 5717 -7904
rect 6874 -7947 6876 -7913
rect 6905 -7947 6953 -7913
rect 7001 -7947 7049 -7913
rect 7097 -7947 7145 -7913
rect 7193 -7947 7241 -7913
rect 7289 -7947 7337 -7913
rect 7385 -7947 7433 -7913
rect 7481 -7947 7529 -7913
rect 7577 -7947 7625 -7913
rect 7654 -7947 7656 -7913
rect 3219 -7966 5724 -7958
rect 5766 -7966 5780 -7958
rect 3219 -8023 5717 -7966
rect 5721 -7972 5780 -7966
rect 5826 -7972 5840 -7950
rect 5720 -8000 5780 -7972
rect 5720 -8006 5768 -8000
rect 5792 -8006 5840 -7972
rect 3219 -8034 5724 -8023
rect 5766 -8034 5780 -8023
rect 3219 -8137 5717 -8034
rect 5721 -8068 5780 -8034
rect 3219 -8148 5724 -8137
rect 5766 -8148 5780 -8137
rect 2395 -8217 2407 -8201
rect 2133 -8319 2147 -8311
rect 891 -8364 939 -8330
rect 963 -8364 1011 -8330
rect 1035 -8364 1083 -8330
rect 1393 -8337 1407 -8326
rect 1493 -8337 1507 -8326
rect 1348 -8371 1407 -8337
rect 1504 -8371 1552 -8337
rect 2088 -8353 2147 -8319
rect 39 -8417 87 -8383
rect 135 -8417 183 -8383
rect 231 -8417 279 -8383
rect 327 -8417 375 -8383
rect 423 -8417 471 -8383
rect 500 -8417 502 -8383
rect 1316 -8407 1364 -8373
rect 1388 -8407 1436 -8373
rect 1747 -8380 1761 -8369
rect 1847 -8380 1861 -8369
rect 2275 -8371 2294 -8303
rect 2316 -8337 2328 -8269
rect 2361 -8301 2373 -8233
rect 2395 -8251 2453 -8217
rect 2395 -8267 2407 -8251
rect 2606 -8296 2654 -8262
rect 2375 -8319 2389 -8311
rect 2386 -8353 2434 -8319
rect 2606 -8364 2654 -8330
rect 1702 -8414 1761 -8380
rect 1858 -8414 1906 -8380
rect 554 -8460 556 -8426
rect 585 -8460 633 -8426
rect 681 -8460 729 -8426
rect 777 -8460 825 -8426
rect 873 -8460 921 -8426
rect 969 -8460 1017 -8426
rect 1065 -8460 1113 -8426
rect 1161 -8460 1209 -8426
rect 1238 -8460 1240 -8426
rect 1670 -8450 1718 -8416
rect 1742 -8450 1790 -8416
rect 2133 -8419 2147 -8408
rect 2088 -8453 2147 -8419
rect 2275 -8459 2289 -8371
rect 2655 -8380 2667 -8246
rect 2375 -8419 2389 -8408
rect 2689 -8414 2701 -8220
rect 2729 -8236 2743 -8225
rect 2725 -8267 2743 -8236
rect 3051 -8254 3099 -8220
rect 2386 -8453 2434 -8419
rect 2629 -8449 2643 -8438
rect 1292 -8503 1294 -8469
rect 1323 -8503 1371 -8469
rect 1419 -8503 1467 -8469
rect 1515 -8503 1563 -8469
rect 1592 -8503 1594 -8469
rect 2024 -8493 2072 -8459
rect 2096 -8493 2144 -8459
rect 2168 -8493 2216 -8459
rect 2240 -8487 2289 -8459
rect 2584 -8483 2643 -8449
rect 2725 -8450 2737 -8267
rect 2771 -8270 2785 -8267
rect 3108 -8270 3115 -8200
rect 2759 -8453 2785 -8270
rect 2787 -8318 2835 -8284
rect 3142 -8304 3149 -8198
rect 3219 -8205 5717 -8148
rect 5721 -8182 5780 -8148
rect 3219 -8216 5724 -8205
rect 5766 -8216 5780 -8205
rect 3219 -8290 5717 -8216
rect 5721 -8250 5780 -8216
rect 5826 -8266 5840 -8006
rect 5860 -7958 5874 -7950
rect 5926 -7958 5940 -7950
rect 5860 -7966 5880 -7958
rect 5922 -7966 5940 -7958
rect 5860 -8023 5874 -7966
rect 5877 -8000 5940 -7966
rect 5926 -8023 5940 -8000
rect 5860 -8034 5880 -8023
rect 5922 -8034 5940 -8023
rect 5860 -8137 5874 -8034
rect 5877 -8068 5940 -8034
rect 5926 -8137 5940 -8068
rect 5860 -8148 5880 -8137
rect 5922 -8148 5940 -8137
rect 5860 -8205 5874 -8148
rect 5877 -8182 5940 -8148
rect 5877 -8205 5925 -8203
rect 5926 -8205 5940 -8182
rect 5860 -8216 5940 -8205
rect 2787 -8386 2835 -8352
rect 2839 -8453 2851 -8318
rect 3190 -8342 5717 -8290
rect 5777 -8342 5825 -8338
rect 2873 -8438 2885 -8350
rect 3190 -8358 5825 -8342
rect 3035 -8366 3049 -8358
rect 2990 -8400 3049 -8366
rect 3135 -8370 3149 -8359
rect 3181 -8370 5825 -8358
rect 3146 -8372 5825 -8370
rect 3146 -8385 5805 -8372
rect 3146 -8404 5783 -8385
rect 5826 -8388 5840 -8322
rect 2871 -8449 2885 -8438
rect 2240 -8493 2288 -8487
rect 1646 -8546 1648 -8512
rect 1677 -8546 1725 -8512
rect 1773 -8546 1821 -8512
rect 1869 -8546 1917 -8512
rect 1946 -8546 1948 -8512
rect 2771 -8534 2785 -8453
rect 2873 -8483 2930 -8449
rect 3035 -8466 3049 -8455
rect 3135 -8462 3149 -8451
rect 3181 -8462 5783 -8404
rect 5860 -8410 5874 -8216
rect 5877 -8250 5940 -8216
rect 5926 -8410 5940 -8250
rect 5960 -7972 5974 -7950
rect 6022 -7966 6036 -7958
rect 6078 -7966 6092 -7958
rect 6033 -7972 6092 -7966
rect 6138 -7972 6152 -7950
rect 5960 -8006 6008 -7972
rect 6032 -8000 6092 -7972
rect 6032 -8006 6080 -8000
rect 6104 -8006 6152 -7972
rect 5960 -8266 5974 -8006
rect 6022 -8034 6036 -8023
rect 6078 -8034 6092 -8023
rect 6033 -8068 6092 -8034
rect 6022 -8148 6036 -8137
rect 6078 -8148 6092 -8137
rect 6033 -8182 6092 -8148
rect 6022 -8216 6036 -8205
rect 6078 -8216 6092 -8205
rect 6033 -8250 6092 -8216
rect 6138 -8266 6152 -8006
rect 6172 -7958 6186 -7950
rect 6238 -7958 6252 -7950
rect 6172 -7966 6192 -7958
rect 6234 -7966 6252 -7958
rect 6172 -8023 6186 -7966
rect 6189 -8000 6252 -7966
rect 6238 -8023 6252 -8000
rect 6172 -8034 6192 -8023
rect 6234 -8034 6252 -8023
rect 6172 -8137 6186 -8034
rect 6189 -8068 6252 -8034
rect 6238 -8137 6252 -8068
rect 6172 -8148 6192 -8137
rect 6234 -8148 6252 -8137
rect 6172 -8205 6186 -8148
rect 6189 -8182 6252 -8148
rect 6189 -8205 6237 -8203
rect 6238 -8205 6252 -8182
rect 6172 -8216 6252 -8205
rect 5960 -8388 5974 -8322
rect 5976 -8351 6024 -8338
rect 6089 -8351 6137 -8338
rect 5976 -8372 6045 -8351
rect 5997 -8385 6045 -8372
rect 6069 -8372 6137 -8351
rect 6069 -8385 6117 -8372
rect 6138 -8388 6152 -8322
rect 5860 -8418 5879 -8410
rect 5921 -8418 5940 -8410
rect 6172 -8410 6186 -8216
rect 6189 -8250 6252 -8216
rect 6238 -8410 6252 -8250
rect 6272 -7972 6286 -7950
rect 6334 -7966 6348 -7958
rect 6390 -7966 6404 -7958
rect 6345 -7972 6404 -7966
rect 6450 -7972 6464 -7950
rect 6272 -8006 6320 -7972
rect 6344 -8000 6404 -7972
rect 6344 -8006 6392 -8000
rect 6416 -8006 6464 -7972
rect 6272 -8266 6286 -8006
rect 6334 -8034 6348 -8023
rect 6390 -8034 6404 -8023
rect 6345 -8068 6404 -8034
rect 6334 -8148 6348 -8137
rect 6390 -8148 6404 -8137
rect 6345 -8182 6404 -8148
rect 6334 -8216 6348 -8205
rect 6390 -8216 6404 -8205
rect 6345 -8250 6404 -8216
rect 6450 -8266 6464 -8006
rect 6484 -7958 6498 -7950
rect 6550 -7958 6564 -7950
rect 6484 -7966 6504 -7958
rect 6546 -7966 6564 -7958
rect 6484 -8023 6498 -7966
rect 6501 -8000 6564 -7966
rect 6550 -8023 6564 -8000
rect 6484 -8034 6504 -8023
rect 6546 -8034 6564 -8023
rect 6484 -8137 6498 -8034
rect 6501 -8068 6564 -8034
rect 6550 -8137 6564 -8068
rect 6484 -8148 6504 -8137
rect 6546 -8148 6564 -8137
rect 6484 -8205 6498 -8148
rect 6501 -8182 6564 -8148
rect 6501 -8205 6549 -8203
rect 6550 -8205 6564 -8182
rect 6484 -8216 6564 -8205
rect 6272 -8388 6286 -8322
rect 6288 -8351 6336 -8338
rect 6401 -8351 6449 -8338
rect 6288 -8372 6357 -8351
rect 6309 -8385 6357 -8372
rect 6381 -8372 6449 -8351
rect 6381 -8385 6429 -8372
rect 6450 -8388 6464 -8322
rect 2990 -8500 3049 -8466
rect 3146 -8496 5783 -8462
rect 2883 -8536 2931 -8502
rect 2955 -8536 3003 -8502
rect 3027 -8536 3075 -8502
rect 3181 -8508 5783 -8496
rect 2000 -8589 2002 -8555
rect 2031 -8589 2079 -8555
rect 2127 -8589 2175 -8555
rect 2223 -8589 2271 -8555
rect 2319 -8589 2367 -8555
rect 2415 -8589 2463 -8555
rect 2492 -8589 2494 -8555
rect 3190 -8598 5783 -8508
rect 5826 -8576 5840 -8422
rect 5860 -8481 5874 -8418
rect 5876 -8452 5940 -8418
rect 6080 -8422 6091 -8411
rect 6172 -8418 6191 -8410
rect 6233 -8418 6252 -8410
rect 6484 -8410 6498 -8216
rect 6501 -8250 6564 -8216
rect 6550 -8300 6564 -8250
rect 6584 -7972 6598 -7966
rect 6646 -7970 6660 -7959
rect 6657 -7972 6705 -7970
rect 6584 -8006 6641 -7972
rect 6657 -8004 6713 -7972
rect 7708 -7990 7710 -7956
rect 7739 -7990 7787 -7956
rect 7835 -7990 7883 -7956
rect 7931 -7990 7979 -7956
rect 8027 -7990 8075 -7956
rect 8123 -7990 8171 -7956
rect 8219 -7990 8267 -7956
rect 8315 -7990 8363 -7956
rect 8411 -7990 8459 -7956
rect 8507 -7990 8555 -7956
rect 8603 -7990 8651 -7956
rect 8699 -7990 8747 -7956
rect 8795 -7990 8843 -7956
rect 8891 -7990 8939 -7956
rect 8987 -7990 9035 -7956
rect 9083 -7990 9131 -7956
rect 9179 -7990 9227 -7956
rect 9275 -7990 9323 -7956
rect 9371 -7990 9419 -7956
rect 9467 -7990 9515 -7956
rect 9563 -7990 9611 -7956
rect 9659 -7990 9707 -7956
rect 9755 -7990 9803 -7956
rect 9851 -7990 9899 -7956
rect 9947 -7990 9995 -7956
rect 10043 -7990 10091 -7956
rect 10139 -7990 10187 -7956
rect 10235 -7990 10283 -7956
rect 10331 -7990 10379 -7956
rect 10408 -7990 10410 -7956
rect 7150 -8001 7162 -7993
rect 6665 -8006 6713 -8004
rect 6584 -8266 6598 -8006
rect 6987 -8009 7001 -8001
rect 7087 -8009 7101 -8001
rect 7143 -8009 7162 -8001
rect 6646 -8038 6660 -8027
rect 6657 -8072 6705 -8038
rect 6898 -8043 7018 -8009
rect 7098 -8043 7162 -8009
rect 7150 -8081 7162 -8043
rect 6987 -8092 7001 -8081
rect 7087 -8092 7101 -8081
rect 7143 -8092 7162 -8081
rect 6942 -8126 7001 -8092
rect 7098 -8126 7162 -8092
rect 6646 -8144 6660 -8133
rect 6657 -8178 6705 -8144
rect 7150 -8165 7162 -8126
rect 6987 -8176 7001 -8165
rect 7087 -8176 7101 -8165
rect 7143 -8176 7162 -8165
rect 6646 -8212 6660 -8201
rect 6942 -8210 7001 -8176
rect 7098 -8210 7162 -8176
rect 6657 -8246 6705 -8212
rect 7150 -8248 7162 -8210
rect 6987 -8259 7001 -8248
rect 7087 -8259 7101 -8248
rect 7143 -8259 7162 -8248
rect 6942 -8293 7001 -8259
rect 7098 -8293 7162 -8259
rect 7184 -8009 7196 -7993
rect 7243 -8009 7257 -8001
rect 7299 -8009 7313 -8001
rect 7376 -8009 7388 -7993
rect 7410 -8001 7422 -7993
rect 7464 -8001 7474 -7993
rect 7399 -8009 7422 -8001
rect 7455 -8009 7474 -8001
rect 7184 -8043 7238 -8009
rect 7254 -8043 7313 -8009
rect 7334 -8043 7388 -8009
rect 7184 -8288 7196 -8043
rect 7243 -8090 7257 -8079
rect 7299 -8090 7313 -8079
rect 7254 -8124 7313 -8090
rect 7243 -8173 7257 -8162
rect 7299 -8173 7313 -8162
rect 7254 -8207 7313 -8173
rect 7243 -8254 7257 -8243
rect 7299 -8254 7313 -8243
rect 7254 -8288 7313 -8254
rect 7376 -8288 7388 -8043
rect 7410 -8043 7474 -8009
rect 7410 -8081 7422 -8043
rect 7464 -8081 7474 -8043
rect 7399 -8092 7422 -8081
rect 7455 -8092 7474 -8081
rect 7410 -8126 7474 -8092
rect 7410 -8165 7422 -8126
rect 7464 -8165 7474 -8126
rect 7399 -8176 7422 -8165
rect 7455 -8176 7474 -8165
rect 7410 -8210 7474 -8176
rect 7410 -8248 7422 -8210
rect 7464 -8248 7474 -8210
rect 7399 -8259 7422 -8248
rect 7455 -8259 7474 -8248
rect 7150 -8322 7162 -8293
rect 7410 -8293 7474 -8259
rect 7498 -8009 7508 -7993
rect 7555 -8009 7569 -8001
rect 7498 -8043 7552 -8009
rect 7566 -8043 7624 -8009
rect 10462 -8033 10464 -7999
rect 10493 -8033 10541 -7999
rect 10589 -8033 10637 -7999
rect 10685 -8033 10733 -7999
rect 10781 -8033 10829 -7999
rect 10877 -8033 10925 -7999
rect 10973 -8033 11021 -7999
rect 11069 -8033 11117 -7999
rect 11165 -8033 11213 -7999
rect 11242 -8033 11244 -7999
rect 7498 -8288 7508 -8043
rect 7954 -8044 7968 -8036
rect 7794 -8056 7808 -8045
rect 7894 -8052 7908 -8044
rect 7950 -8052 7968 -8044
rect 7749 -8058 7808 -8056
rect 7555 -8090 7569 -8079
rect 7733 -8090 7853 -8058
rect 7905 -8086 7968 -8052
rect 7566 -8124 7614 -8090
rect 7733 -8092 7781 -8090
rect 7805 -8092 7853 -8090
rect 7954 -8109 7968 -8086
rect 7794 -8124 7808 -8113
rect 7894 -8120 7908 -8109
rect 7950 -8120 7968 -8109
rect 7749 -8158 7808 -8124
rect 7905 -8154 7968 -8120
rect 7555 -8173 7569 -8162
rect 7566 -8207 7614 -8173
rect 7794 -8230 7808 -8219
rect 7954 -8223 7968 -8154
rect 7555 -8254 7569 -8243
rect 7566 -8288 7614 -8254
rect 7749 -8264 7808 -8230
rect 7894 -8234 7908 -8223
rect 7950 -8234 7968 -8223
rect 7905 -8268 7968 -8234
rect 7410 -8322 7422 -8293
rect 7464 -8322 7474 -8293
rect 7794 -8298 7808 -8287
rect 7905 -8291 7953 -8289
rect 7954 -8291 7968 -8268
rect 7749 -8332 7808 -8298
rect 7894 -8302 7968 -8291
rect 7905 -8336 7968 -8302
rect 6550 -8410 6564 -8388
rect 5926 -8481 5940 -8452
rect 5860 -8492 5879 -8481
rect 5921 -8492 5940 -8481
rect 5860 -8542 5874 -8492
rect 5876 -8526 5940 -8492
rect 5926 -8542 5940 -8526
rect 5960 -8576 5974 -8422
rect 6032 -8456 6091 -8422
rect 6021 -8495 6035 -8484
rect 6077 -8495 6091 -8484
rect 6032 -8529 6091 -8495
rect 6138 -8576 6152 -8422
rect 6172 -8481 6186 -8418
rect 6188 -8452 6252 -8418
rect 6392 -8422 6403 -8411
rect 6484 -8418 6503 -8410
rect 6545 -8418 6564 -8410
rect 6238 -8481 6252 -8452
rect 6172 -8492 6191 -8481
rect 6233 -8492 6252 -8481
rect 6172 -8542 6186 -8492
rect 6188 -8526 6252 -8492
rect 6238 -8542 6252 -8526
rect 6272 -8576 6286 -8422
rect 6344 -8456 6403 -8422
rect 6333 -8495 6347 -8484
rect 6389 -8495 6403 -8484
rect 6344 -8529 6403 -8495
rect 6450 -8576 6464 -8422
rect 6484 -8481 6498 -8418
rect 6500 -8452 6564 -8418
rect 6550 -8481 6564 -8452
rect 6484 -8492 6503 -8481
rect 6545 -8492 6564 -8481
rect 6484 -8542 6498 -8492
rect 6500 -8526 6564 -8492
rect 6550 -8542 6564 -8526
rect 6584 -8576 6598 -8422
rect 6656 -8456 6704 -8422
rect 6915 -8428 6963 -8394
rect 6983 -8428 7031 -8394
rect 7051 -8428 7099 -8394
rect 7119 -8428 7167 -8394
rect 7187 -8428 7235 -8394
rect 7255 -8428 7303 -8394
rect 7323 -8428 7371 -8394
rect 7391 -8428 7439 -8394
rect 7443 -8428 7455 -8394
rect 7477 -8462 7489 -8360
rect 6645 -8495 6659 -8484
rect 6987 -8495 7001 -8487
rect 7087 -8495 7101 -8487
rect 7143 -8495 7157 -8487
rect 7399 -8495 7413 -8487
rect 7455 -8495 7469 -8487
rect 6656 -8529 6704 -8495
rect 6942 -8529 7001 -8495
rect 7098 -8498 7157 -8495
rect 7098 -8529 7146 -8498
rect 2546 -8632 2548 -8598
rect 2577 -8632 2625 -8598
rect 2673 -8632 2721 -8598
rect 2769 -8632 2817 -8598
rect 2865 -8632 2913 -8598
rect 2961 -8632 3009 -8598
rect 3057 -8632 3105 -8598
rect 3153 -8632 5783 -8598
rect 5792 -8616 5840 -8582
rect 5960 -8616 6008 -8582
rect 6032 -8616 6080 -8582
rect 6104 -8616 6152 -8582
rect 6272 -8616 6320 -8582
rect 6344 -8616 6392 -8582
rect 6416 -8616 6464 -8582
rect 6593 -8616 6641 -8582
rect 6665 -8616 6713 -8582
rect 6987 -8595 7001 -8584
rect 7087 -8595 7101 -8584
rect 7134 -8595 7146 -8529
rect 6942 -8629 7001 -8595
rect 7098 -8629 7146 -8595
rect 3190 -8658 5783 -8632
rect 3219 -8684 5783 -8658
rect 6898 -8665 6946 -8631
rect 6970 -8665 7018 -8631
rect 7134 -8645 7146 -8629
rect 7168 -8631 7180 -8534
rect 7243 -8565 7257 -8554
rect 7299 -8565 7313 -8554
rect 7254 -8599 7313 -8565
rect 7360 -8631 7372 -8534
rect 7168 -8665 7222 -8631
rect 7246 -8665 7294 -8631
rect 7318 -8665 7372 -8631
rect 7394 -8584 7406 -8500
rect 7410 -8529 7469 -8495
rect 7394 -8595 7413 -8584
rect 7455 -8595 7469 -8584
rect 7394 -8645 7406 -8595
rect 7410 -8629 7469 -8595
rect 7516 -8645 7525 -8445
rect 7550 -8487 7559 -8479
rect 7550 -8495 7569 -8487
rect 7550 -8584 7559 -8495
rect 7566 -8529 7614 -8495
rect 7954 -8496 7968 -8336
rect 7988 -8058 8002 -8036
rect 8050 -8052 8064 -8044
rect 8106 -8052 8120 -8044
rect 8061 -8058 8120 -8052
rect 8166 -8058 8180 -8036
rect 7988 -8092 8036 -8058
rect 8060 -8086 8120 -8058
rect 8060 -8092 8108 -8086
rect 8132 -8092 8180 -8058
rect 7988 -8352 8002 -8092
rect 8050 -8120 8064 -8109
rect 8106 -8120 8120 -8109
rect 8061 -8154 8120 -8120
rect 8050 -8234 8064 -8223
rect 8106 -8234 8120 -8223
rect 8061 -8268 8120 -8234
rect 8050 -8302 8064 -8291
rect 8106 -8302 8120 -8291
rect 8061 -8336 8120 -8302
rect 8166 -8352 8180 -8092
rect 8200 -8044 8214 -8036
rect 8266 -8044 8280 -8036
rect 8200 -8052 8220 -8044
rect 8262 -8052 8280 -8044
rect 8200 -8109 8214 -8052
rect 8217 -8086 8280 -8052
rect 8266 -8109 8280 -8086
rect 8200 -8120 8220 -8109
rect 8262 -8120 8280 -8109
rect 8200 -8223 8214 -8120
rect 8217 -8154 8280 -8120
rect 8266 -8223 8280 -8154
rect 8200 -8234 8220 -8223
rect 8262 -8234 8280 -8223
rect 8200 -8291 8214 -8234
rect 8217 -8268 8280 -8234
rect 8217 -8291 8265 -8289
rect 8266 -8291 8280 -8268
rect 8200 -8302 8280 -8291
rect 7988 -8474 8002 -8408
rect 8004 -8437 8052 -8424
rect 8117 -8437 8165 -8424
rect 8004 -8458 8075 -8437
rect 8027 -8471 8075 -8458
rect 8099 -8458 8165 -8437
rect 8099 -8471 8147 -8458
rect 8166 -8474 8180 -8408
rect 7793 -8508 7807 -8497
rect 7893 -8504 7907 -8496
rect 7949 -8504 7968 -8496
rect 8200 -8496 8214 -8302
rect 8217 -8336 8280 -8302
rect 8266 -8496 8280 -8336
rect 8300 -8058 8314 -8036
rect 8362 -8052 8376 -8044
rect 8418 -8052 8432 -8044
rect 8373 -8058 8432 -8052
rect 8478 -8058 8492 -8036
rect 8300 -8092 8348 -8058
rect 8372 -8086 8432 -8058
rect 8372 -8092 8420 -8086
rect 8444 -8092 8492 -8058
rect 8300 -8352 8314 -8092
rect 8362 -8120 8376 -8109
rect 8418 -8120 8432 -8109
rect 8373 -8154 8432 -8120
rect 8362 -8234 8376 -8223
rect 8418 -8234 8432 -8223
rect 8373 -8268 8432 -8234
rect 8362 -8302 8376 -8291
rect 8418 -8302 8432 -8291
rect 8373 -8336 8432 -8302
rect 8478 -8352 8492 -8092
rect 8512 -8044 8526 -8036
rect 8578 -8044 8592 -8036
rect 8512 -8052 8532 -8044
rect 8574 -8052 8592 -8044
rect 8512 -8109 8526 -8052
rect 8529 -8086 8592 -8052
rect 8578 -8109 8592 -8086
rect 8512 -8120 8532 -8109
rect 8574 -8120 8592 -8109
rect 8512 -8223 8526 -8120
rect 8529 -8154 8592 -8120
rect 8578 -8223 8592 -8154
rect 8512 -8234 8532 -8223
rect 8574 -8234 8592 -8223
rect 8512 -8291 8526 -8234
rect 8529 -8268 8592 -8234
rect 8529 -8291 8577 -8289
rect 8578 -8291 8592 -8268
rect 8512 -8302 8592 -8291
rect 8300 -8474 8314 -8408
rect 8316 -8437 8364 -8424
rect 8429 -8437 8477 -8424
rect 8316 -8458 8385 -8437
rect 8337 -8471 8385 -8458
rect 8409 -8458 8477 -8437
rect 8409 -8471 8457 -8458
rect 8478 -8474 8492 -8408
rect 7748 -8542 7807 -8508
rect 7904 -8538 7968 -8504
rect 8108 -8508 8119 -8497
rect 8200 -8504 8219 -8496
rect 8261 -8504 8280 -8496
rect 8512 -8496 8526 -8302
rect 8529 -8336 8592 -8302
rect 8578 -8496 8592 -8336
rect 8612 -8058 8626 -8036
rect 8674 -8052 8688 -8044
rect 8730 -8052 8744 -8044
rect 8685 -8058 8744 -8052
rect 8790 -8058 8804 -8036
rect 8612 -8092 8660 -8058
rect 8684 -8086 8744 -8058
rect 8684 -8092 8732 -8086
rect 8756 -8092 8804 -8058
rect 8612 -8352 8626 -8092
rect 8674 -8120 8688 -8109
rect 8730 -8120 8744 -8109
rect 8685 -8154 8744 -8120
rect 8674 -8234 8688 -8223
rect 8730 -8234 8744 -8223
rect 8685 -8268 8744 -8234
rect 8674 -8302 8688 -8291
rect 8730 -8302 8744 -8291
rect 8685 -8336 8744 -8302
rect 8790 -8352 8804 -8092
rect 8824 -8044 8838 -8036
rect 8890 -8044 8904 -8036
rect 8824 -8052 8844 -8044
rect 8886 -8052 8904 -8044
rect 8824 -8109 8838 -8052
rect 8841 -8086 8904 -8052
rect 8890 -8109 8904 -8086
rect 8824 -8120 8844 -8109
rect 8886 -8120 8904 -8109
rect 8824 -8223 8838 -8120
rect 8841 -8154 8904 -8120
rect 8890 -8223 8904 -8154
rect 8824 -8234 8844 -8223
rect 8886 -8234 8904 -8223
rect 8824 -8291 8838 -8234
rect 8841 -8268 8904 -8234
rect 8841 -8291 8889 -8289
rect 8890 -8291 8904 -8268
rect 8824 -8302 8904 -8291
rect 8612 -8474 8626 -8408
rect 8628 -8437 8676 -8424
rect 8741 -8437 8789 -8424
rect 8628 -8458 8697 -8437
rect 8649 -8471 8697 -8458
rect 8721 -8458 8789 -8437
rect 8721 -8471 8769 -8458
rect 8790 -8474 8804 -8408
rect 7954 -8567 7968 -8538
rect 7793 -8581 7807 -8570
rect 7893 -8578 7907 -8567
rect 7949 -8578 7968 -8567
rect 7550 -8595 7569 -8584
rect 7550 -8631 7559 -8595
rect 7566 -8629 7614 -8595
rect 7748 -8615 7807 -8581
rect 7904 -8612 7968 -8578
rect 7954 -8628 7968 -8612
rect 7168 -8671 7180 -8665
rect 7360 -8671 7372 -8665
rect 7550 -8665 7604 -8631
rect 7988 -8662 8002 -8508
rect 8060 -8542 8119 -8508
rect 8049 -8581 8063 -8570
rect 8105 -8581 8119 -8570
rect 8060 -8615 8119 -8581
rect 8166 -8662 8180 -8508
rect 8200 -8567 8214 -8504
rect 8216 -8538 8280 -8504
rect 8420 -8508 8431 -8497
rect 8512 -8504 8531 -8496
rect 8573 -8504 8592 -8496
rect 8824 -8496 8838 -8302
rect 8841 -8336 8904 -8302
rect 8890 -8496 8904 -8336
rect 8924 -8058 8938 -8036
rect 8986 -8052 9000 -8044
rect 9042 -8052 9056 -8044
rect 8997 -8058 9056 -8052
rect 9102 -8058 9116 -8036
rect 8924 -8092 8972 -8058
rect 8996 -8086 9056 -8058
rect 8996 -8092 9044 -8086
rect 9068 -8092 9116 -8058
rect 8924 -8352 8938 -8092
rect 8986 -8120 9000 -8109
rect 9042 -8120 9056 -8109
rect 8997 -8154 9056 -8120
rect 8986 -8234 9000 -8223
rect 9042 -8234 9056 -8223
rect 8997 -8268 9056 -8234
rect 8986 -8302 9000 -8291
rect 9042 -8302 9056 -8291
rect 8997 -8336 9056 -8302
rect 9102 -8352 9116 -8092
rect 9136 -8044 9150 -8036
rect 9202 -8044 9216 -8036
rect 9136 -8052 9156 -8044
rect 9198 -8052 9216 -8044
rect 9136 -8109 9150 -8052
rect 9153 -8086 9216 -8052
rect 9202 -8109 9216 -8086
rect 9136 -8120 9156 -8109
rect 9198 -8120 9216 -8109
rect 9136 -8223 9150 -8120
rect 9153 -8154 9216 -8120
rect 9202 -8223 9216 -8154
rect 9136 -8234 9156 -8223
rect 9198 -8234 9216 -8223
rect 9136 -8291 9150 -8234
rect 9153 -8268 9216 -8234
rect 9153 -8291 9201 -8289
rect 9202 -8291 9216 -8268
rect 9136 -8302 9216 -8291
rect 8924 -8474 8938 -8408
rect 8940 -8437 8988 -8424
rect 9053 -8437 9101 -8424
rect 8940 -8458 9009 -8437
rect 8961 -8471 9009 -8458
rect 9033 -8458 9101 -8437
rect 9033 -8471 9081 -8458
rect 9102 -8474 9116 -8408
rect 8266 -8567 8280 -8538
rect 8200 -8578 8219 -8567
rect 8261 -8578 8280 -8567
rect 8200 -8628 8214 -8578
rect 8216 -8612 8280 -8578
rect 8266 -8628 8280 -8612
rect 8300 -8662 8314 -8508
rect 8372 -8542 8431 -8508
rect 8361 -8581 8375 -8570
rect 8417 -8581 8431 -8570
rect 8372 -8615 8431 -8581
rect 8478 -8662 8492 -8508
rect 8512 -8567 8526 -8504
rect 8528 -8538 8592 -8504
rect 8732 -8508 8743 -8497
rect 8824 -8504 8843 -8496
rect 8885 -8504 8904 -8496
rect 9136 -8496 9150 -8302
rect 9153 -8336 9216 -8302
rect 9202 -8496 9216 -8336
rect 9236 -8058 9250 -8036
rect 9298 -8052 9312 -8044
rect 9354 -8052 9368 -8044
rect 9309 -8058 9368 -8052
rect 9414 -8058 9428 -8036
rect 9236 -8092 9284 -8058
rect 9308 -8086 9368 -8058
rect 9308 -8092 9356 -8086
rect 9380 -8092 9428 -8058
rect 9236 -8352 9250 -8092
rect 9298 -8120 9312 -8109
rect 9354 -8120 9368 -8109
rect 9309 -8154 9368 -8120
rect 9298 -8234 9312 -8223
rect 9354 -8234 9368 -8223
rect 9309 -8268 9368 -8234
rect 9298 -8302 9312 -8291
rect 9354 -8302 9368 -8291
rect 9309 -8336 9368 -8302
rect 9414 -8352 9428 -8092
rect 9448 -8044 9462 -8036
rect 9514 -8044 9528 -8036
rect 9448 -8052 9468 -8044
rect 9510 -8052 9528 -8044
rect 9448 -8109 9462 -8052
rect 9465 -8086 9528 -8052
rect 9514 -8109 9528 -8086
rect 9448 -8120 9468 -8109
rect 9510 -8120 9528 -8109
rect 9448 -8223 9462 -8120
rect 9465 -8154 9528 -8120
rect 9514 -8223 9528 -8154
rect 9448 -8234 9468 -8223
rect 9510 -8234 9528 -8223
rect 9448 -8291 9462 -8234
rect 9465 -8268 9528 -8234
rect 9465 -8291 9513 -8289
rect 9514 -8291 9528 -8268
rect 9448 -8302 9528 -8291
rect 9236 -8474 9250 -8408
rect 9252 -8437 9300 -8424
rect 9365 -8437 9413 -8424
rect 9252 -8458 9321 -8437
rect 9273 -8471 9321 -8458
rect 9345 -8458 9413 -8437
rect 9345 -8471 9393 -8458
rect 9414 -8474 9428 -8408
rect 8578 -8567 8592 -8538
rect 8512 -8578 8531 -8567
rect 8573 -8578 8592 -8567
rect 8512 -8628 8526 -8578
rect 8528 -8612 8592 -8578
rect 8578 -8628 8592 -8612
rect 8612 -8662 8626 -8508
rect 8684 -8542 8743 -8508
rect 8673 -8581 8687 -8570
rect 8729 -8581 8743 -8570
rect 8684 -8615 8743 -8581
rect 8790 -8662 8804 -8508
rect 8824 -8567 8838 -8504
rect 8840 -8538 8904 -8504
rect 9044 -8508 9055 -8497
rect 9136 -8504 9155 -8496
rect 9197 -8504 9216 -8496
rect 9448 -8496 9462 -8302
rect 9465 -8336 9528 -8302
rect 9514 -8496 9528 -8336
rect 9548 -8058 9562 -8036
rect 9610 -8052 9624 -8044
rect 9666 -8052 9680 -8044
rect 9621 -8058 9680 -8052
rect 9726 -8058 9740 -8036
rect 9548 -8092 9596 -8058
rect 9620 -8086 9680 -8058
rect 9620 -8092 9668 -8086
rect 9692 -8092 9740 -8058
rect 9548 -8352 9562 -8092
rect 9610 -8120 9624 -8109
rect 9666 -8120 9680 -8109
rect 9621 -8154 9680 -8120
rect 9610 -8234 9624 -8223
rect 9666 -8234 9680 -8223
rect 9621 -8268 9680 -8234
rect 9610 -8302 9624 -8291
rect 9666 -8302 9680 -8291
rect 9621 -8336 9680 -8302
rect 9726 -8352 9740 -8092
rect 9760 -8044 9774 -8036
rect 9826 -8044 9840 -8036
rect 9760 -8052 9780 -8044
rect 9822 -8052 9840 -8044
rect 9760 -8109 9774 -8052
rect 9777 -8086 9840 -8052
rect 9826 -8109 9840 -8086
rect 9760 -8120 9780 -8109
rect 9822 -8120 9840 -8109
rect 9760 -8223 9774 -8120
rect 9777 -8154 9840 -8120
rect 9826 -8223 9840 -8154
rect 9760 -8234 9780 -8223
rect 9822 -8234 9840 -8223
rect 9760 -8291 9774 -8234
rect 9777 -8268 9840 -8234
rect 9777 -8291 9825 -8289
rect 9826 -8291 9840 -8268
rect 9760 -8302 9840 -8291
rect 9548 -8474 9562 -8408
rect 9564 -8437 9612 -8424
rect 9677 -8437 9725 -8424
rect 9564 -8458 9633 -8437
rect 9585 -8471 9633 -8458
rect 9657 -8458 9725 -8437
rect 9657 -8471 9705 -8458
rect 9726 -8474 9740 -8408
rect 8890 -8567 8904 -8538
rect 8824 -8578 8843 -8567
rect 8885 -8578 8904 -8567
rect 8824 -8628 8838 -8578
rect 8840 -8612 8904 -8578
rect 8890 -8628 8904 -8612
rect 8924 -8662 8938 -8508
rect 8996 -8542 9055 -8508
rect 8985 -8581 8999 -8570
rect 9041 -8581 9055 -8570
rect 8996 -8615 9055 -8581
rect 9102 -8662 9116 -8508
rect 9136 -8567 9150 -8504
rect 9152 -8538 9216 -8504
rect 9356 -8508 9367 -8497
rect 9448 -8504 9467 -8496
rect 9509 -8504 9528 -8496
rect 9760 -8496 9774 -8302
rect 9777 -8336 9840 -8302
rect 9826 -8496 9840 -8336
rect 9860 -8058 9874 -8036
rect 9922 -8052 9936 -8044
rect 9978 -8052 9992 -8044
rect 9933 -8058 9992 -8052
rect 10038 -8058 10052 -8036
rect 9860 -8092 9908 -8058
rect 9932 -8086 9992 -8058
rect 9932 -8092 9980 -8086
rect 10004 -8092 10052 -8058
rect 9860 -8352 9874 -8092
rect 9922 -8120 9936 -8109
rect 9978 -8120 9992 -8109
rect 9933 -8154 9992 -8120
rect 9922 -8234 9936 -8223
rect 9978 -8234 9992 -8223
rect 9933 -8268 9992 -8234
rect 9922 -8302 9936 -8291
rect 9978 -8302 9992 -8291
rect 9933 -8336 9992 -8302
rect 10038 -8352 10052 -8092
rect 10072 -8044 10086 -8036
rect 10138 -8044 10152 -8036
rect 10072 -8052 10092 -8044
rect 10134 -8052 10152 -8044
rect 10072 -8109 10086 -8052
rect 10089 -8086 10152 -8052
rect 10138 -8109 10152 -8086
rect 10072 -8120 10092 -8109
rect 10134 -8120 10152 -8109
rect 10072 -8223 10086 -8120
rect 10089 -8154 10152 -8120
rect 10138 -8223 10152 -8154
rect 10072 -8234 10092 -8223
rect 10134 -8234 10152 -8223
rect 10072 -8291 10086 -8234
rect 10089 -8268 10152 -8234
rect 10089 -8291 10137 -8289
rect 10138 -8291 10152 -8268
rect 10072 -8302 10152 -8291
rect 9860 -8474 9874 -8408
rect 9876 -8437 9924 -8424
rect 9989 -8437 10037 -8424
rect 9876 -8458 9945 -8437
rect 9897 -8471 9945 -8458
rect 9969 -8458 10037 -8437
rect 9969 -8471 10017 -8458
rect 10038 -8474 10052 -8408
rect 9202 -8567 9216 -8538
rect 9136 -8578 9155 -8567
rect 9197 -8578 9216 -8567
rect 9136 -8628 9150 -8578
rect 9152 -8612 9216 -8578
rect 9202 -8628 9216 -8612
rect 9236 -8662 9250 -8508
rect 9308 -8542 9367 -8508
rect 9297 -8581 9311 -8570
rect 9353 -8581 9367 -8570
rect 9308 -8615 9367 -8581
rect 9414 -8662 9428 -8508
rect 9448 -8567 9462 -8504
rect 9464 -8538 9528 -8504
rect 9668 -8508 9679 -8497
rect 9760 -8504 9779 -8496
rect 9821 -8504 9840 -8496
rect 10072 -8496 10086 -8302
rect 10089 -8336 10152 -8302
rect 10138 -8386 10152 -8336
rect 10172 -8058 10186 -8052
rect 10234 -8056 10248 -8045
rect 10245 -8058 10293 -8056
rect 10172 -8092 10229 -8058
rect 10245 -8090 10301 -8058
rect 11296 -8076 11298 -8042
rect 11327 -8076 11375 -8042
rect 11423 -8076 11471 -8042
rect 11519 -8076 11567 -8042
rect 11615 -8076 11663 -8042
rect 11711 -8076 11759 -8042
rect 11807 -8076 11855 -8042
rect 11903 -8076 11951 -8042
rect 11999 -8076 12047 -8042
rect 12095 -8076 12143 -8042
rect 12191 -8076 12239 -8042
rect 12287 -8076 12335 -8042
rect 12383 -8076 12431 -8042
rect 12479 -8076 12527 -8042
rect 12575 -8076 12623 -8042
rect 12671 -8076 12719 -8042
rect 12767 -8076 12815 -8042
rect 12863 -8076 12911 -8042
rect 12959 -8076 13007 -8042
rect 13055 -8076 13103 -8042
rect 13151 -8076 13199 -8042
rect 13247 -8076 13295 -8042
rect 13343 -8076 13391 -8042
rect 13439 -8076 13487 -8042
rect 13535 -8076 13583 -8042
rect 13631 -8076 13679 -8042
rect 13727 -8076 13775 -8042
rect 13823 -8076 13871 -8042
rect 13919 -8076 13967 -8042
rect 13996 -8076 13998 -8042
rect 10738 -8087 10750 -8079
rect 10253 -8092 10301 -8090
rect 10172 -8352 10186 -8092
rect 10575 -8095 10589 -8087
rect 10675 -8095 10689 -8087
rect 10731 -8095 10750 -8087
rect 10234 -8124 10248 -8113
rect 10245 -8158 10293 -8124
rect 10486 -8129 10606 -8095
rect 10686 -8129 10750 -8095
rect 10738 -8167 10750 -8129
rect 10575 -8178 10589 -8167
rect 10675 -8178 10689 -8167
rect 10731 -8178 10750 -8167
rect 10530 -8212 10589 -8178
rect 10686 -8212 10750 -8178
rect 10234 -8230 10248 -8219
rect 10245 -8264 10293 -8230
rect 10738 -8251 10750 -8212
rect 10575 -8262 10589 -8251
rect 10675 -8262 10689 -8251
rect 10731 -8262 10750 -8251
rect 10234 -8298 10248 -8287
rect 10530 -8296 10589 -8262
rect 10686 -8296 10750 -8262
rect 10245 -8332 10293 -8298
rect 10738 -8334 10750 -8296
rect 10575 -8345 10589 -8334
rect 10675 -8345 10689 -8334
rect 10731 -8345 10750 -8334
rect 10530 -8379 10589 -8345
rect 10686 -8379 10750 -8345
rect 10772 -8095 10784 -8079
rect 10831 -8095 10845 -8087
rect 10887 -8095 10901 -8087
rect 10964 -8095 10976 -8079
rect 10998 -8087 11010 -8079
rect 11052 -8087 11062 -8079
rect 10987 -8095 11010 -8087
rect 11043 -8095 11062 -8087
rect 10772 -8129 10826 -8095
rect 10842 -8129 10901 -8095
rect 10922 -8129 10976 -8095
rect 10772 -8374 10784 -8129
rect 10831 -8176 10845 -8165
rect 10887 -8176 10901 -8165
rect 10842 -8210 10901 -8176
rect 10831 -8259 10845 -8248
rect 10887 -8259 10901 -8248
rect 10842 -8293 10901 -8259
rect 10831 -8340 10845 -8329
rect 10887 -8340 10901 -8329
rect 10842 -8374 10901 -8340
rect 10964 -8374 10976 -8129
rect 10998 -8129 11062 -8095
rect 10998 -8167 11010 -8129
rect 11052 -8167 11062 -8129
rect 10987 -8178 11010 -8167
rect 11043 -8178 11062 -8167
rect 10998 -8212 11062 -8178
rect 10998 -8251 11010 -8212
rect 11052 -8251 11062 -8212
rect 10987 -8262 11010 -8251
rect 11043 -8262 11062 -8251
rect 10998 -8296 11062 -8262
rect 10998 -8334 11010 -8296
rect 11052 -8334 11062 -8296
rect 10987 -8345 11010 -8334
rect 11043 -8345 11062 -8334
rect 10738 -8408 10750 -8379
rect 10998 -8379 11062 -8345
rect 11086 -8095 11096 -8079
rect 11143 -8095 11157 -8087
rect 11086 -8129 11140 -8095
rect 11154 -8129 11212 -8095
rect 14050 -8119 14052 -8085
rect 14081 -8119 14129 -8085
rect 14177 -8119 14225 -8085
rect 14273 -8119 14321 -8085
rect 14369 -8119 14417 -8085
rect 14465 -8119 14513 -8085
rect 14561 -8119 14609 -8085
rect 14657 -8119 14705 -8085
rect 14753 -8119 14801 -8085
rect 14830 -8119 14832 -8085
rect 11086 -8374 11096 -8129
rect 11542 -8130 11556 -8122
rect 11382 -8142 11396 -8131
rect 11482 -8138 11496 -8130
rect 11538 -8138 11556 -8130
rect 11337 -8144 11396 -8142
rect 11143 -8176 11157 -8165
rect 11321 -8176 11441 -8144
rect 11493 -8172 11556 -8138
rect 11154 -8210 11202 -8176
rect 11321 -8178 11369 -8176
rect 11393 -8178 11441 -8176
rect 11542 -8195 11556 -8172
rect 11382 -8210 11396 -8199
rect 11482 -8206 11496 -8195
rect 11538 -8206 11556 -8195
rect 11337 -8244 11396 -8210
rect 11493 -8240 11556 -8206
rect 11143 -8259 11157 -8248
rect 11154 -8293 11202 -8259
rect 11382 -8316 11396 -8305
rect 11542 -8309 11556 -8240
rect 11143 -8340 11157 -8329
rect 11154 -8374 11202 -8340
rect 11337 -8350 11396 -8316
rect 11482 -8320 11496 -8309
rect 11538 -8320 11556 -8309
rect 11493 -8354 11556 -8320
rect 10998 -8408 11010 -8379
rect 11052 -8408 11062 -8379
rect 11382 -8384 11396 -8373
rect 11493 -8377 11541 -8375
rect 11542 -8377 11556 -8354
rect 11337 -8418 11396 -8384
rect 11482 -8388 11556 -8377
rect 11493 -8422 11556 -8388
rect 10138 -8496 10152 -8474
rect 9514 -8567 9528 -8538
rect 9448 -8578 9467 -8567
rect 9509 -8578 9528 -8567
rect 9448 -8628 9462 -8578
rect 9464 -8612 9528 -8578
rect 9514 -8628 9528 -8612
rect 9548 -8662 9562 -8508
rect 9620 -8542 9679 -8508
rect 9609 -8581 9623 -8570
rect 9665 -8581 9679 -8570
rect 9620 -8615 9679 -8581
rect 9726 -8662 9740 -8508
rect 9760 -8567 9774 -8504
rect 9776 -8538 9840 -8504
rect 9980 -8508 9991 -8497
rect 10072 -8504 10091 -8496
rect 10133 -8504 10152 -8496
rect 9826 -8567 9840 -8538
rect 9760 -8578 9779 -8567
rect 9821 -8578 9840 -8567
rect 9760 -8628 9774 -8578
rect 9776 -8612 9840 -8578
rect 9826 -8628 9840 -8612
rect 9860 -8662 9874 -8508
rect 9932 -8542 9991 -8508
rect 9921 -8581 9935 -8570
rect 9977 -8581 9991 -8570
rect 9932 -8615 9991 -8581
rect 10038 -8662 10052 -8508
rect 10072 -8567 10086 -8504
rect 10088 -8538 10152 -8504
rect 10138 -8567 10152 -8538
rect 10072 -8578 10091 -8567
rect 10133 -8578 10152 -8567
rect 10072 -8628 10086 -8578
rect 10088 -8612 10152 -8578
rect 10138 -8628 10152 -8612
rect 10172 -8662 10186 -8508
rect 10244 -8542 10292 -8508
rect 10503 -8514 10551 -8480
rect 10571 -8514 10619 -8480
rect 10639 -8514 10687 -8480
rect 10707 -8514 10755 -8480
rect 10775 -8514 10823 -8480
rect 10843 -8514 10891 -8480
rect 10911 -8514 10959 -8480
rect 10979 -8514 11027 -8480
rect 11031 -8514 11043 -8480
rect 11065 -8548 11077 -8446
rect 10233 -8581 10247 -8570
rect 10575 -8581 10589 -8573
rect 10675 -8581 10689 -8573
rect 10731 -8581 10745 -8573
rect 10987 -8581 11001 -8573
rect 11043 -8581 11057 -8573
rect 10244 -8615 10292 -8581
rect 10530 -8615 10589 -8581
rect 10686 -8584 10745 -8581
rect 10686 -8615 10734 -8584
rect 7550 -8671 7559 -8665
rect 3219 -8718 5831 -8684
rect 5879 -8718 5927 -8684
rect 5975 -8718 6023 -8684
rect 6071 -8718 6119 -8684
rect 6167 -8718 6215 -8684
rect 6263 -8718 6311 -8684
rect 6359 -8718 6407 -8684
rect 6455 -8718 6503 -8684
rect 6551 -8718 6599 -8684
rect 6647 -8718 6695 -8684
rect 6743 -8718 6791 -8684
rect 6820 -8718 6822 -8684
rect 7727 -8702 7775 -8668
rect 7799 -8702 7847 -8668
rect 7988 -8702 8036 -8668
rect 8060 -8702 8108 -8668
rect 8132 -8702 8180 -8668
rect 8300 -8702 8348 -8668
rect 8372 -8702 8420 -8668
rect 8444 -8702 8492 -8668
rect 8612 -8702 8660 -8668
rect 8684 -8702 8732 -8668
rect 8756 -8702 8804 -8668
rect 8924 -8702 8972 -8668
rect 8996 -8702 9044 -8668
rect 9068 -8702 9116 -8668
rect 9236 -8702 9284 -8668
rect 9308 -8702 9356 -8668
rect 9380 -8702 9428 -8668
rect 9548 -8702 9596 -8668
rect 9620 -8702 9668 -8668
rect 9692 -8702 9740 -8668
rect 9860 -8702 9908 -8668
rect 9932 -8702 9980 -8668
rect 10004 -8702 10052 -8668
rect 10181 -8702 10229 -8668
rect 10253 -8702 10301 -8668
rect 10575 -8681 10589 -8670
rect 10675 -8681 10689 -8670
rect 10722 -8681 10734 -8615
rect 10530 -8715 10589 -8681
rect 10686 -8715 10734 -8681
rect 3219 -8744 5783 -8718
rect 3219 -11123 5717 -8744
rect 6874 -8761 6876 -8727
rect 6905 -8761 6953 -8727
rect 7001 -8761 7049 -8727
rect 7097 -8761 7145 -8727
rect 7193 -8761 7241 -8727
rect 7289 -8761 7337 -8727
rect 7385 -8761 7433 -8727
rect 7481 -8761 7529 -8727
rect 7577 -8761 7625 -8727
rect 7654 -8761 7656 -8727
rect 10486 -8751 10534 -8717
rect 10558 -8751 10606 -8717
rect 10722 -8731 10734 -8715
rect 10756 -8717 10768 -8620
rect 10831 -8651 10845 -8640
rect 10887 -8651 10901 -8640
rect 10842 -8685 10901 -8651
rect 10948 -8717 10960 -8620
rect 10756 -8751 10810 -8717
rect 10834 -8751 10882 -8717
rect 10906 -8751 10960 -8717
rect 10982 -8670 10994 -8586
rect 10998 -8615 11057 -8581
rect 10982 -8681 11001 -8670
rect 11043 -8681 11057 -8670
rect 10982 -8731 10994 -8681
rect 10998 -8715 11057 -8681
rect 11104 -8731 11113 -8531
rect 11138 -8573 11147 -8565
rect 11138 -8581 11157 -8573
rect 11138 -8670 11147 -8581
rect 11154 -8615 11202 -8581
rect 11542 -8582 11556 -8422
rect 11576 -8144 11590 -8122
rect 11638 -8138 11652 -8130
rect 11694 -8138 11708 -8130
rect 11649 -8144 11708 -8138
rect 11754 -8144 11768 -8122
rect 11576 -8178 11624 -8144
rect 11648 -8172 11708 -8144
rect 11648 -8178 11696 -8172
rect 11720 -8178 11768 -8144
rect 11576 -8438 11590 -8178
rect 11638 -8206 11652 -8195
rect 11694 -8206 11708 -8195
rect 11649 -8240 11708 -8206
rect 11638 -8320 11652 -8309
rect 11694 -8320 11708 -8309
rect 11649 -8354 11708 -8320
rect 11638 -8388 11652 -8377
rect 11694 -8388 11708 -8377
rect 11649 -8422 11708 -8388
rect 11754 -8438 11768 -8178
rect 11788 -8130 11802 -8122
rect 11854 -8130 11868 -8122
rect 11788 -8138 11808 -8130
rect 11850 -8138 11868 -8130
rect 11788 -8195 11802 -8138
rect 11805 -8172 11868 -8138
rect 11854 -8195 11868 -8172
rect 11788 -8206 11808 -8195
rect 11850 -8206 11868 -8195
rect 11788 -8309 11802 -8206
rect 11805 -8240 11868 -8206
rect 11854 -8309 11868 -8240
rect 11788 -8320 11808 -8309
rect 11850 -8320 11868 -8309
rect 11788 -8377 11802 -8320
rect 11805 -8354 11868 -8320
rect 11805 -8377 11853 -8375
rect 11854 -8377 11868 -8354
rect 11788 -8388 11868 -8377
rect 11576 -8560 11590 -8494
rect 11592 -8523 11640 -8510
rect 11705 -8523 11753 -8510
rect 11592 -8544 11663 -8523
rect 11615 -8557 11663 -8544
rect 11687 -8544 11753 -8523
rect 11687 -8557 11735 -8544
rect 11754 -8560 11768 -8494
rect 11381 -8594 11395 -8583
rect 11481 -8590 11495 -8582
rect 11537 -8590 11556 -8582
rect 11788 -8582 11802 -8388
rect 11805 -8422 11868 -8388
rect 11854 -8582 11868 -8422
rect 11888 -8144 11902 -8122
rect 11950 -8138 11964 -8130
rect 12006 -8138 12020 -8130
rect 11961 -8144 12020 -8138
rect 12066 -8144 12080 -8122
rect 11888 -8178 11936 -8144
rect 11960 -8172 12020 -8144
rect 11960 -8178 12008 -8172
rect 12032 -8178 12080 -8144
rect 11888 -8438 11902 -8178
rect 11950 -8206 11964 -8195
rect 12006 -8206 12020 -8195
rect 11961 -8240 12020 -8206
rect 11950 -8320 11964 -8309
rect 12006 -8320 12020 -8309
rect 11961 -8354 12020 -8320
rect 11950 -8388 11964 -8377
rect 12006 -8388 12020 -8377
rect 11961 -8422 12020 -8388
rect 12066 -8438 12080 -8178
rect 12100 -8130 12114 -8122
rect 12166 -8130 12180 -8122
rect 12100 -8138 12120 -8130
rect 12162 -8138 12180 -8130
rect 12100 -8195 12114 -8138
rect 12117 -8172 12180 -8138
rect 12166 -8195 12180 -8172
rect 12100 -8206 12120 -8195
rect 12162 -8206 12180 -8195
rect 12100 -8309 12114 -8206
rect 12117 -8240 12180 -8206
rect 12166 -8309 12180 -8240
rect 12100 -8320 12120 -8309
rect 12162 -8320 12180 -8309
rect 12100 -8377 12114 -8320
rect 12117 -8354 12180 -8320
rect 12117 -8377 12165 -8375
rect 12166 -8377 12180 -8354
rect 12100 -8388 12180 -8377
rect 11888 -8560 11902 -8494
rect 11904 -8523 11952 -8510
rect 12017 -8523 12065 -8510
rect 11904 -8544 11973 -8523
rect 11925 -8557 11973 -8544
rect 11997 -8544 12065 -8523
rect 11997 -8557 12045 -8544
rect 12066 -8560 12080 -8494
rect 11336 -8628 11395 -8594
rect 11492 -8624 11556 -8590
rect 11696 -8594 11707 -8583
rect 11788 -8590 11807 -8582
rect 11849 -8590 11868 -8582
rect 12100 -8582 12114 -8388
rect 12117 -8422 12180 -8388
rect 12166 -8582 12180 -8422
rect 12200 -8144 12214 -8122
rect 12262 -8138 12276 -8130
rect 12318 -8138 12332 -8130
rect 12273 -8144 12332 -8138
rect 12378 -8144 12392 -8122
rect 12200 -8178 12248 -8144
rect 12272 -8172 12332 -8144
rect 12272 -8178 12320 -8172
rect 12344 -8178 12392 -8144
rect 12200 -8438 12214 -8178
rect 12262 -8206 12276 -8195
rect 12318 -8206 12332 -8195
rect 12273 -8240 12332 -8206
rect 12262 -8320 12276 -8309
rect 12318 -8320 12332 -8309
rect 12273 -8354 12332 -8320
rect 12262 -8388 12276 -8377
rect 12318 -8388 12332 -8377
rect 12273 -8422 12332 -8388
rect 12378 -8438 12392 -8178
rect 12412 -8130 12426 -8122
rect 12478 -8130 12492 -8122
rect 12412 -8138 12432 -8130
rect 12474 -8138 12492 -8130
rect 12412 -8195 12426 -8138
rect 12429 -8172 12492 -8138
rect 12478 -8195 12492 -8172
rect 12412 -8206 12432 -8195
rect 12474 -8206 12492 -8195
rect 12412 -8309 12426 -8206
rect 12429 -8240 12492 -8206
rect 12478 -8309 12492 -8240
rect 12412 -8320 12432 -8309
rect 12474 -8320 12492 -8309
rect 12412 -8377 12426 -8320
rect 12429 -8354 12492 -8320
rect 12429 -8377 12477 -8375
rect 12478 -8377 12492 -8354
rect 12412 -8388 12492 -8377
rect 12200 -8560 12214 -8494
rect 12216 -8523 12264 -8510
rect 12329 -8523 12377 -8510
rect 12216 -8544 12285 -8523
rect 12237 -8557 12285 -8544
rect 12309 -8544 12377 -8523
rect 12309 -8557 12357 -8544
rect 12378 -8560 12392 -8494
rect 11542 -8653 11556 -8624
rect 11381 -8667 11395 -8656
rect 11481 -8664 11495 -8653
rect 11537 -8664 11556 -8653
rect 11138 -8681 11157 -8670
rect 11138 -8717 11147 -8681
rect 11154 -8715 11202 -8681
rect 11336 -8701 11395 -8667
rect 11492 -8698 11556 -8664
rect 11542 -8714 11556 -8698
rect 10756 -8757 10768 -8751
rect 10948 -8757 10960 -8751
rect 11138 -8751 11192 -8717
rect 11576 -8748 11590 -8594
rect 11648 -8628 11707 -8594
rect 11637 -8667 11651 -8656
rect 11693 -8667 11707 -8656
rect 11648 -8701 11707 -8667
rect 11754 -8748 11768 -8594
rect 11788 -8653 11802 -8590
rect 11804 -8624 11868 -8590
rect 12008 -8594 12019 -8583
rect 12100 -8590 12119 -8582
rect 12161 -8590 12180 -8582
rect 12412 -8582 12426 -8388
rect 12429 -8422 12492 -8388
rect 12478 -8582 12492 -8422
rect 12512 -8144 12526 -8122
rect 12574 -8138 12588 -8130
rect 12630 -8138 12644 -8130
rect 12585 -8144 12644 -8138
rect 12690 -8144 12704 -8122
rect 12512 -8178 12560 -8144
rect 12584 -8172 12644 -8144
rect 12584 -8178 12632 -8172
rect 12656 -8178 12704 -8144
rect 12512 -8438 12526 -8178
rect 12574 -8206 12588 -8195
rect 12630 -8206 12644 -8195
rect 12585 -8240 12644 -8206
rect 12574 -8320 12588 -8309
rect 12630 -8320 12644 -8309
rect 12585 -8354 12644 -8320
rect 12574 -8388 12588 -8377
rect 12630 -8388 12644 -8377
rect 12585 -8422 12644 -8388
rect 12690 -8438 12704 -8178
rect 12724 -8130 12738 -8122
rect 12790 -8130 12804 -8122
rect 12724 -8138 12744 -8130
rect 12786 -8138 12804 -8130
rect 12724 -8195 12738 -8138
rect 12741 -8172 12804 -8138
rect 12790 -8195 12804 -8172
rect 12724 -8206 12744 -8195
rect 12786 -8206 12804 -8195
rect 12724 -8309 12738 -8206
rect 12741 -8240 12804 -8206
rect 12790 -8309 12804 -8240
rect 12724 -8320 12744 -8309
rect 12786 -8320 12804 -8309
rect 12724 -8377 12738 -8320
rect 12741 -8354 12804 -8320
rect 12741 -8377 12789 -8375
rect 12790 -8377 12804 -8354
rect 12724 -8388 12804 -8377
rect 12512 -8560 12526 -8494
rect 12528 -8523 12576 -8510
rect 12641 -8523 12689 -8510
rect 12528 -8544 12597 -8523
rect 12549 -8557 12597 -8544
rect 12621 -8544 12689 -8523
rect 12621 -8557 12669 -8544
rect 12690 -8560 12704 -8494
rect 11854 -8653 11868 -8624
rect 11788 -8664 11807 -8653
rect 11849 -8664 11868 -8653
rect 11788 -8714 11802 -8664
rect 11804 -8698 11868 -8664
rect 11854 -8714 11868 -8698
rect 11888 -8748 11902 -8594
rect 11960 -8628 12019 -8594
rect 11949 -8667 11963 -8656
rect 12005 -8667 12019 -8656
rect 11960 -8701 12019 -8667
rect 12066 -8748 12080 -8594
rect 12100 -8653 12114 -8590
rect 12116 -8624 12180 -8590
rect 12320 -8594 12331 -8583
rect 12412 -8590 12431 -8582
rect 12473 -8590 12492 -8582
rect 12724 -8582 12738 -8388
rect 12741 -8422 12804 -8388
rect 12790 -8582 12804 -8422
rect 12824 -8144 12838 -8122
rect 12886 -8138 12900 -8130
rect 12942 -8138 12956 -8130
rect 12897 -8144 12956 -8138
rect 13002 -8144 13016 -8122
rect 12824 -8178 12872 -8144
rect 12896 -8172 12956 -8144
rect 12896 -8178 12944 -8172
rect 12968 -8178 13016 -8144
rect 12824 -8438 12838 -8178
rect 12886 -8206 12900 -8195
rect 12942 -8206 12956 -8195
rect 12897 -8240 12956 -8206
rect 12886 -8320 12900 -8309
rect 12942 -8320 12956 -8309
rect 12897 -8354 12956 -8320
rect 12886 -8388 12900 -8377
rect 12942 -8388 12956 -8377
rect 12897 -8422 12956 -8388
rect 13002 -8438 13016 -8178
rect 13036 -8130 13050 -8122
rect 13102 -8130 13116 -8122
rect 13036 -8138 13056 -8130
rect 13098 -8138 13116 -8130
rect 13036 -8195 13050 -8138
rect 13053 -8172 13116 -8138
rect 13102 -8195 13116 -8172
rect 13036 -8206 13056 -8195
rect 13098 -8206 13116 -8195
rect 13036 -8309 13050 -8206
rect 13053 -8240 13116 -8206
rect 13102 -8309 13116 -8240
rect 13036 -8320 13056 -8309
rect 13098 -8320 13116 -8309
rect 13036 -8377 13050 -8320
rect 13053 -8354 13116 -8320
rect 13053 -8377 13101 -8375
rect 13102 -8377 13116 -8354
rect 13036 -8388 13116 -8377
rect 12824 -8560 12838 -8494
rect 12840 -8523 12888 -8510
rect 12953 -8523 13001 -8510
rect 12840 -8544 12909 -8523
rect 12861 -8557 12909 -8544
rect 12933 -8544 13001 -8523
rect 12933 -8557 12981 -8544
rect 13002 -8560 13016 -8494
rect 12166 -8653 12180 -8624
rect 12100 -8664 12119 -8653
rect 12161 -8664 12180 -8653
rect 12100 -8714 12114 -8664
rect 12116 -8698 12180 -8664
rect 12166 -8714 12180 -8698
rect 12200 -8748 12214 -8594
rect 12272 -8628 12331 -8594
rect 12261 -8667 12275 -8656
rect 12317 -8667 12331 -8656
rect 12272 -8701 12331 -8667
rect 12378 -8748 12392 -8594
rect 12412 -8653 12426 -8590
rect 12428 -8624 12492 -8590
rect 12632 -8594 12643 -8583
rect 12724 -8590 12743 -8582
rect 12785 -8590 12804 -8582
rect 13036 -8582 13050 -8388
rect 13053 -8422 13116 -8388
rect 13102 -8582 13116 -8422
rect 13136 -8144 13150 -8122
rect 13198 -8138 13212 -8130
rect 13254 -8138 13268 -8130
rect 13209 -8144 13268 -8138
rect 13314 -8144 13328 -8122
rect 13136 -8178 13184 -8144
rect 13208 -8172 13268 -8144
rect 13208 -8178 13256 -8172
rect 13280 -8178 13328 -8144
rect 13136 -8438 13150 -8178
rect 13198 -8206 13212 -8195
rect 13254 -8206 13268 -8195
rect 13209 -8240 13268 -8206
rect 13198 -8320 13212 -8309
rect 13254 -8320 13268 -8309
rect 13209 -8354 13268 -8320
rect 13198 -8388 13212 -8377
rect 13254 -8388 13268 -8377
rect 13209 -8422 13268 -8388
rect 13314 -8438 13328 -8178
rect 13348 -8130 13362 -8122
rect 13414 -8130 13428 -8122
rect 13348 -8138 13368 -8130
rect 13410 -8138 13428 -8130
rect 13348 -8195 13362 -8138
rect 13365 -8172 13428 -8138
rect 13414 -8195 13428 -8172
rect 13348 -8206 13368 -8195
rect 13410 -8206 13428 -8195
rect 13348 -8309 13362 -8206
rect 13365 -8240 13428 -8206
rect 13414 -8309 13428 -8240
rect 13348 -8320 13368 -8309
rect 13410 -8320 13428 -8309
rect 13348 -8377 13362 -8320
rect 13365 -8354 13428 -8320
rect 13365 -8377 13413 -8375
rect 13414 -8377 13428 -8354
rect 13348 -8388 13428 -8377
rect 13136 -8560 13150 -8494
rect 13152 -8523 13200 -8510
rect 13265 -8523 13313 -8510
rect 13152 -8544 13221 -8523
rect 13173 -8557 13221 -8544
rect 13245 -8544 13313 -8523
rect 13245 -8557 13293 -8544
rect 13314 -8560 13328 -8494
rect 12478 -8653 12492 -8624
rect 12412 -8664 12431 -8653
rect 12473 -8664 12492 -8653
rect 12412 -8714 12426 -8664
rect 12428 -8698 12492 -8664
rect 12478 -8714 12492 -8698
rect 12512 -8748 12526 -8594
rect 12584 -8628 12643 -8594
rect 12573 -8667 12587 -8656
rect 12629 -8667 12643 -8656
rect 12584 -8701 12643 -8667
rect 12690 -8748 12704 -8594
rect 12724 -8653 12738 -8590
rect 12740 -8624 12804 -8590
rect 12944 -8594 12955 -8583
rect 13036 -8590 13055 -8582
rect 13097 -8590 13116 -8582
rect 13348 -8582 13362 -8388
rect 13365 -8422 13428 -8388
rect 13414 -8582 13428 -8422
rect 13448 -8144 13462 -8122
rect 13510 -8138 13524 -8130
rect 13566 -8138 13580 -8130
rect 13521 -8144 13580 -8138
rect 13626 -8144 13640 -8122
rect 13448 -8178 13496 -8144
rect 13520 -8172 13580 -8144
rect 13520 -8178 13568 -8172
rect 13592 -8178 13640 -8144
rect 13448 -8438 13462 -8178
rect 13510 -8206 13524 -8195
rect 13566 -8206 13580 -8195
rect 13521 -8240 13580 -8206
rect 13510 -8320 13524 -8309
rect 13566 -8320 13580 -8309
rect 13521 -8354 13580 -8320
rect 13510 -8388 13524 -8377
rect 13566 -8388 13580 -8377
rect 13521 -8422 13580 -8388
rect 13626 -8438 13640 -8178
rect 13660 -8130 13674 -8122
rect 13726 -8130 13740 -8122
rect 13660 -8138 13680 -8130
rect 13722 -8138 13740 -8130
rect 13660 -8195 13674 -8138
rect 13677 -8172 13740 -8138
rect 13726 -8195 13740 -8172
rect 13660 -8206 13680 -8195
rect 13722 -8206 13740 -8195
rect 13660 -8309 13674 -8206
rect 13677 -8240 13740 -8206
rect 13726 -8309 13740 -8240
rect 13660 -8320 13680 -8309
rect 13722 -8320 13740 -8309
rect 13660 -8377 13674 -8320
rect 13677 -8354 13740 -8320
rect 13677 -8377 13725 -8375
rect 13726 -8377 13740 -8354
rect 13660 -8388 13740 -8377
rect 13448 -8560 13462 -8494
rect 13464 -8523 13512 -8510
rect 13577 -8523 13625 -8510
rect 13464 -8544 13533 -8523
rect 13485 -8557 13533 -8544
rect 13557 -8544 13625 -8523
rect 13557 -8557 13605 -8544
rect 13626 -8560 13640 -8494
rect 12790 -8653 12804 -8624
rect 12724 -8664 12743 -8653
rect 12785 -8664 12804 -8653
rect 12724 -8714 12738 -8664
rect 12740 -8698 12804 -8664
rect 12790 -8714 12804 -8698
rect 12824 -8748 12838 -8594
rect 12896 -8628 12955 -8594
rect 12885 -8667 12899 -8656
rect 12941 -8667 12955 -8656
rect 12896 -8701 12955 -8667
rect 13002 -8748 13016 -8594
rect 13036 -8653 13050 -8590
rect 13052 -8624 13116 -8590
rect 13256 -8594 13267 -8583
rect 13348 -8590 13367 -8582
rect 13409 -8590 13428 -8582
rect 13660 -8582 13674 -8388
rect 13677 -8422 13740 -8388
rect 13726 -8472 13740 -8422
rect 13760 -8144 13774 -8138
rect 13822 -8142 13836 -8131
rect 13833 -8144 13881 -8142
rect 13760 -8178 13817 -8144
rect 13833 -8176 13889 -8144
rect 14884 -8162 14886 -8128
rect 14915 -8162 14963 -8128
rect 15011 -8162 15059 -8128
rect 15107 -8162 15155 -8128
rect 15203 -8162 15251 -8128
rect 15299 -8162 15347 -8128
rect 15395 -8162 15443 -8128
rect 15491 -8162 15539 -8128
rect 15587 -8162 15635 -8128
rect 15683 -8162 15731 -8128
rect 15779 -8162 15827 -8128
rect 15875 -8162 15923 -8128
rect 15971 -8162 16019 -8128
rect 16067 -8162 16115 -8128
rect 16163 -8162 16211 -8128
rect 16259 -8162 16307 -8128
rect 16355 -8162 16403 -8128
rect 16451 -8162 16499 -8128
rect 16547 -8162 16595 -8128
rect 16643 -8162 16691 -8128
rect 16739 -8162 16787 -8128
rect 16835 -8162 16883 -8128
rect 16931 -8162 16979 -8128
rect 17027 -8162 17075 -8128
rect 17123 -8162 17171 -8128
rect 17219 -8162 17267 -8128
rect 17315 -8162 17363 -8128
rect 17411 -8162 17459 -8128
rect 17507 -8162 17555 -8128
rect 14326 -8173 14338 -8165
rect 13841 -8178 13889 -8176
rect 13760 -8438 13774 -8178
rect 14163 -8181 14177 -8173
rect 14263 -8181 14277 -8173
rect 14319 -8181 14338 -8173
rect 13822 -8210 13836 -8199
rect 13833 -8244 13881 -8210
rect 14074 -8215 14194 -8181
rect 14274 -8215 14338 -8181
rect 14326 -8253 14338 -8215
rect 14163 -8264 14177 -8253
rect 14263 -8264 14277 -8253
rect 14319 -8264 14338 -8253
rect 14118 -8298 14177 -8264
rect 14274 -8298 14338 -8264
rect 13822 -8316 13836 -8305
rect 13833 -8350 13881 -8316
rect 14326 -8337 14338 -8298
rect 14163 -8348 14177 -8337
rect 14263 -8348 14277 -8337
rect 14319 -8348 14338 -8337
rect 13822 -8384 13836 -8373
rect 14118 -8382 14177 -8348
rect 14274 -8382 14338 -8348
rect 13833 -8418 13881 -8384
rect 14326 -8420 14338 -8382
rect 14163 -8431 14177 -8420
rect 14263 -8431 14277 -8420
rect 14319 -8431 14338 -8420
rect 14118 -8465 14177 -8431
rect 14274 -8465 14338 -8431
rect 14360 -8181 14372 -8165
rect 14419 -8181 14433 -8173
rect 14475 -8181 14489 -8173
rect 14552 -8181 14564 -8165
rect 14586 -8173 14598 -8165
rect 14640 -8173 14650 -8165
rect 14575 -8181 14598 -8173
rect 14631 -8181 14650 -8173
rect 14360 -8215 14414 -8181
rect 14430 -8215 14489 -8181
rect 14510 -8215 14564 -8181
rect 14360 -8460 14372 -8215
rect 14419 -8262 14433 -8251
rect 14475 -8262 14489 -8251
rect 14430 -8296 14489 -8262
rect 14419 -8345 14433 -8334
rect 14475 -8345 14489 -8334
rect 14430 -8379 14489 -8345
rect 14419 -8426 14433 -8415
rect 14475 -8426 14489 -8415
rect 14430 -8460 14489 -8426
rect 14552 -8460 14564 -8215
rect 14586 -8215 14650 -8181
rect 14586 -8253 14598 -8215
rect 14640 -8253 14650 -8215
rect 14575 -8264 14598 -8253
rect 14631 -8264 14650 -8253
rect 14586 -8298 14650 -8264
rect 14586 -8337 14598 -8298
rect 14640 -8337 14650 -8298
rect 14575 -8348 14598 -8337
rect 14631 -8348 14650 -8337
rect 14586 -8382 14650 -8348
rect 14586 -8420 14598 -8382
rect 14640 -8420 14650 -8382
rect 14575 -8431 14598 -8420
rect 14631 -8431 14650 -8420
rect 14326 -8494 14338 -8465
rect 14586 -8465 14650 -8431
rect 14674 -8181 14684 -8165
rect 14731 -8181 14745 -8173
rect 14674 -8215 14728 -8181
rect 14742 -8215 14800 -8181
rect 14674 -8460 14684 -8215
rect 15130 -8216 15144 -8208
rect 14970 -8228 14984 -8217
rect 15070 -8224 15084 -8216
rect 15126 -8224 15144 -8216
rect 14925 -8230 14984 -8228
rect 14731 -8262 14745 -8251
rect 14909 -8262 15029 -8230
rect 15081 -8258 15144 -8224
rect 14742 -8296 14790 -8262
rect 14909 -8264 14957 -8262
rect 14981 -8264 15029 -8262
rect 15130 -8281 15144 -8258
rect 14970 -8296 14984 -8285
rect 15070 -8292 15084 -8281
rect 15126 -8292 15144 -8281
rect 14925 -8330 14984 -8296
rect 15081 -8326 15144 -8292
rect 14731 -8345 14745 -8334
rect 14742 -8379 14790 -8345
rect 14970 -8402 14984 -8391
rect 15130 -8395 15144 -8326
rect 14731 -8426 14745 -8415
rect 14742 -8460 14790 -8426
rect 14925 -8436 14984 -8402
rect 15070 -8406 15084 -8395
rect 15126 -8406 15144 -8395
rect 15081 -8440 15144 -8406
rect 14586 -8494 14598 -8465
rect 14640 -8494 14650 -8465
rect 14970 -8470 14984 -8459
rect 15081 -8463 15129 -8461
rect 15130 -8463 15144 -8440
rect 14925 -8504 14984 -8470
rect 15070 -8474 15144 -8463
rect 15081 -8508 15144 -8474
rect 13726 -8582 13740 -8560
rect 13102 -8653 13116 -8624
rect 13036 -8664 13055 -8653
rect 13097 -8664 13116 -8653
rect 13036 -8714 13050 -8664
rect 13052 -8698 13116 -8664
rect 13102 -8714 13116 -8698
rect 13136 -8748 13150 -8594
rect 13208 -8628 13267 -8594
rect 13197 -8667 13211 -8656
rect 13253 -8667 13267 -8656
rect 13208 -8701 13267 -8667
rect 13314 -8748 13328 -8594
rect 13348 -8653 13362 -8590
rect 13364 -8624 13428 -8590
rect 13568 -8594 13579 -8583
rect 13660 -8590 13679 -8582
rect 13721 -8590 13740 -8582
rect 13414 -8653 13428 -8624
rect 13348 -8664 13367 -8653
rect 13409 -8664 13428 -8653
rect 13348 -8714 13362 -8664
rect 13364 -8698 13428 -8664
rect 13414 -8714 13428 -8698
rect 13448 -8748 13462 -8594
rect 13520 -8628 13579 -8594
rect 13509 -8667 13523 -8656
rect 13565 -8667 13579 -8656
rect 13520 -8701 13579 -8667
rect 13626 -8748 13640 -8594
rect 13660 -8653 13674 -8590
rect 13676 -8624 13740 -8590
rect 13726 -8653 13740 -8624
rect 13660 -8664 13679 -8653
rect 13721 -8664 13740 -8653
rect 13660 -8714 13674 -8664
rect 13676 -8698 13740 -8664
rect 13726 -8714 13740 -8698
rect 13760 -8748 13774 -8594
rect 13832 -8628 13880 -8594
rect 14091 -8600 14139 -8566
rect 14159 -8600 14207 -8566
rect 14227 -8600 14275 -8566
rect 14295 -8600 14343 -8566
rect 14363 -8600 14411 -8566
rect 14431 -8600 14479 -8566
rect 14499 -8600 14547 -8566
rect 14567 -8600 14615 -8566
rect 14619 -8600 14631 -8566
rect 14653 -8634 14665 -8532
rect 13821 -8667 13835 -8656
rect 14163 -8667 14177 -8659
rect 14263 -8667 14277 -8659
rect 14319 -8667 14333 -8659
rect 14575 -8667 14589 -8659
rect 14631 -8667 14645 -8659
rect 13832 -8701 13880 -8667
rect 14118 -8701 14177 -8667
rect 14274 -8670 14333 -8667
rect 14274 -8701 14322 -8670
rect 11138 -8757 11147 -8751
rect 7708 -8804 7710 -8770
rect 7739 -8804 7787 -8770
rect 7835 -8804 7883 -8770
rect 7931 -8804 7979 -8770
rect 8027 -8804 8075 -8770
rect 8123 -8804 8171 -8770
rect 8219 -8804 8267 -8770
rect 8315 -8804 8363 -8770
rect 8411 -8804 8459 -8770
rect 8507 -8804 8555 -8770
rect 8603 -8804 8651 -8770
rect 8699 -8804 8747 -8770
rect 8795 -8804 8843 -8770
rect 8891 -8804 8939 -8770
rect 8987 -8804 9035 -8770
rect 9083 -8804 9131 -8770
rect 9179 -8804 9227 -8770
rect 9275 -8804 9323 -8770
rect 9371 -8804 9419 -8770
rect 9467 -8804 9515 -8770
rect 9563 -8804 9611 -8770
rect 9659 -8804 9707 -8770
rect 9755 -8804 9803 -8770
rect 9851 -8804 9899 -8770
rect 9947 -8804 9995 -8770
rect 10043 -8804 10091 -8770
rect 10139 -8804 10187 -8770
rect 10235 -8804 10283 -8770
rect 10331 -8804 10379 -8770
rect 10408 -8804 10410 -8770
rect 11315 -8788 11363 -8754
rect 11387 -8788 11435 -8754
rect 11576 -8788 11624 -8754
rect 11648 -8788 11696 -8754
rect 11720 -8788 11768 -8754
rect 11888 -8788 11936 -8754
rect 11960 -8788 12008 -8754
rect 12032 -8788 12080 -8754
rect 12200 -8788 12248 -8754
rect 12272 -8788 12320 -8754
rect 12344 -8788 12392 -8754
rect 12512 -8788 12560 -8754
rect 12584 -8788 12632 -8754
rect 12656 -8788 12704 -8754
rect 12824 -8788 12872 -8754
rect 12896 -8788 12944 -8754
rect 12968 -8788 13016 -8754
rect 13136 -8788 13184 -8754
rect 13208 -8788 13256 -8754
rect 13280 -8788 13328 -8754
rect 13448 -8788 13496 -8754
rect 13520 -8788 13568 -8754
rect 13592 -8788 13640 -8754
rect 13769 -8788 13817 -8754
rect 13841 -8788 13889 -8754
rect 14163 -8767 14177 -8756
rect 14263 -8767 14277 -8756
rect 14310 -8767 14322 -8701
rect 14118 -8801 14177 -8767
rect 14274 -8801 14322 -8767
rect 10462 -8847 10464 -8813
rect 10493 -8847 10541 -8813
rect 10589 -8847 10637 -8813
rect 10685 -8847 10733 -8813
rect 10781 -8847 10829 -8813
rect 10877 -8847 10925 -8813
rect 10973 -8847 11021 -8813
rect 11069 -8847 11117 -8813
rect 11165 -8847 11213 -8813
rect 11242 -8847 11244 -8813
rect 14074 -8837 14122 -8803
rect 14146 -8837 14194 -8803
rect 14310 -8817 14322 -8801
rect 14344 -8803 14356 -8706
rect 14419 -8737 14433 -8726
rect 14475 -8737 14489 -8726
rect 14430 -8771 14489 -8737
rect 14536 -8803 14548 -8706
rect 14344 -8837 14398 -8803
rect 14422 -8837 14470 -8803
rect 14494 -8837 14548 -8803
rect 14570 -8756 14582 -8672
rect 14586 -8701 14645 -8667
rect 14570 -8767 14589 -8756
rect 14631 -8767 14645 -8756
rect 14570 -8817 14582 -8767
rect 14586 -8801 14645 -8767
rect 14692 -8817 14701 -8617
rect 14726 -8659 14735 -8651
rect 14726 -8667 14745 -8659
rect 14726 -8756 14735 -8667
rect 14742 -8701 14790 -8667
rect 15130 -8668 15144 -8508
rect 15164 -8230 15178 -8208
rect 15226 -8224 15240 -8216
rect 15282 -8224 15296 -8216
rect 15237 -8230 15296 -8224
rect 15342 -8230 15356 -8208
rect 15164 -8264 15212 -8230
rect 15236 -8258 15296 -8230
rect 15236 -8264 15284 -8258
rect 15308 -8264 15356 -8230
rect 15164 -8524 15178 -8264
rect 15226 -8292 15240 -8281
rect 15282 -8292 15296 -8281
rect 15237 -8326 15296 -8292
rect 15226 -8406 15240 -8395
rect 15282 -8406 15296 -8395
rect 15237 -8440 15296 -8406
rect 15226 -8474 15240 -8463
rect 15282 -8474 15296 -8463
rect 15237 -8508 15296 -8474
rect 15342 -8524 15356 -8264
rect 15376 -8216 15390 -8208
rect 15442 -8216 15456 -8208
rect 15376 -8224 15396 -8216
rect 15438 -8224 15456 -8216
rect 15376 -8281 15390 -8224
rect 15393 -8258 15456 -8224
rect 15442 -8281 15456 -8258
rect 15376 -8292 15396 -8281
rect 15438 -8292 15456 -8281
rect 15376 -8395 15390 -8292
rect 15393 -8326 15456 -8292
rect 15442 -8395 15456 -8326
rect 15376 -8406 15396 -8395
rect 15438 -8406 15456 -8395
rect 15376 -8463 15390 -8406
rect 15393 -8440 15456 -8406
rect 15393 -8463 15441 -8461
rect 15442 -8463 15456 -8440
rect 15376 -8474 15456 -8463
rect 15164 -8646 15178 -8580
rect 15180 -8609 15228 -8596
rect 15293 -8609 15341 -8596
rect 15180 -8630 15251 -8609
rect 15203 -8643 15251 -8630
rect 15275 -8630 15341 -8609
rect 15275 -8643 15323 -8630
rect 15342 -8646 15356 -8580
rect 14969 -8680 14983 -8669
rect 15069 -8676 15083 -8668
rect 15125 -8676 15144 -8668
rect 15376 -8668 15390 -8474
rect 15393 -8508 15456 -8474
rect 15442 -8668 15456 -8508
rect 15476 -8230 15490 -8208
rect 15538 -8224 15552 -8216
rect 15594 -8224 15608 -8216
rect 15549 -8230 15608 -8224
rect 15654 -8230 15668 -8208
rect 15476 -8264 15524 -8230
rect 15548 -8258 15608 -8230
rect 15548 -8264 15596 -8258
rect 15620 -8264 15668 -8230
rect 15476 -8524 15490 -8264
rect 15538 -8292 15552 -8281
rect 15594 -8292 15608 -8281
rect 15549 -8326 15608 -8292
rect 15538 -8406 15552 -8395
rect 15594 -8406 15608 -8395
rect 15549 -8440 15608 -8406
rect 15538 -8474 15552 -8463
rect 15594 -8474 15608 -8463
rect 15549 -8508 15608 -8474
rect 15654 -8524 15668 -8264
rect 15688 -8216 15702 -8208
rect 15754 -8216 15768 -8208
rect 15688 -8224 15708 -8216
rect 15750 -8224 15768 -8216
rect 15688 -8281 15702 -8224
rect 15705 -8258 15768 -8224
rect 15754 -8281 15768 -8258
rect 15688 -8292 15708 -8281
rect 15750 -8292 15768 -8281
rect 15688 -8395 15702 -8292
rect 15705 -8326 15768 -8292
rect 15754 -8395 15768 -8326
rect 15688 -8406 15708 -8395
rect 15750 -8406 15768 -8395
rect 15688 -8463 15702 -8406
rect 15705 -8440 15768 -8406
rect 15705 -8463 15753 -8461
rect 15754 -8463 15768 -8440
rect 15688 -8474 15768 -8463
rect 15476 -8646 15490 -8580
rect 15492 -8609 15540 -8596
rect 15605 -8609 15653 -8596
rect 15492 -8630 15561 -8609
rect 15513 -8643 15561 -8630
rect 15585 -8630 15653 -8609
rect 15585 -8643 15633 -8630
rect 15654 -8646 15668 -8580
rect 14924 -8714 14983 -8680
rect 15080 -8710 15144 -8676
rect 15284 -8680 15295 -8669
rect 15376 -8676 15395 -8668
rect 15437 -8676 15456 -8668
rect 15688 -8668 15702 -8474
rect 15705 -8508 15768 -8474
rect 15754 -8668 15768 -8508
rect 15788 -8230 15802 -8208
rect 15850 -8224 15864 -8216
rect 15906 -8224 15920 -8216
rect 15861 -8230 15920 -8224
rect 15966 -8230 15980 -8208
rect 15788 -8264 15836 -8230
rect 15860 -8258 15920 -8230
rect 15860 -8264 15908 -8258
rect 15932 -8264 15980 -8230
rect 15788 -8524 15802 -8264
rect 15850 -8292 15864 -8281
rect 15906 -8292 15920 -8281
rect 15861 -8326 15920 -8292
rect 15850 -8406 15864 -8395
rect 15906 -8406 15920 -8395
rect 15861 -8440 15920 -8406
rect 15850 -8474 15864 -8463
rect 15906 -8474 15920 -8463
rect 15861 -8508 15920 -8474
rect 15966 -8524 15980 -8264
rect 16000 -8216 16014 -8208
rect 16066 -8216 16080 -8208
rect 16000 -8224 16020 -8216
rect 16062 -8224 16080 -8216
rect 16000 -8281 16014 -8224
rect 16017 -8258 16080 -8224
rect 16066 -8281 16080 -8258
rect 16000 -8292 16020 -8281
rect 16062 -8292 16080 -8281
rect 16000 -8395 16014 -8292
rect 16017 -8326 16080 -8292
rect 16066 -8395 16080 -8326
rect 16000 -8406 16020 -8395
rect 16062 -8406 16080 -8395
rect 16000 -8463 16014 -8406
rect 16017 -8440 16080 -8406
rect 16017 -8463 16065 -8461
rect 16066 -8463 16080 -8440
rect 16000 -8474 16080 -8463
rect 15788 -8646 15802 -8580
rect 15804 -8609 15852 -8596
rect 15917 -8609 15965 -8596
rect 15804 -8630 15873 -8609
rect 15825 -8643 15873 -8630
rect 15897 -8630 15965 -8609
rect 15897 -8643 15945 -8630
rect 15966 -8646 15980 -8580
rect 15130 -8739 15144 -8710
rect 14969 -8753 14983 -8742
rect 15069 -8750 15083 -8739
rect 15125 -8750 15144 -8739
rect 14726 -8767 14745 -8756
rect 14726 -8803 14735 -8767
rect 14742 -8801 14790 -8767
rect 14924 -8787 14983 -8753
rect 15080 -8784 15144 -8750
rect 15130 -8800 15144 -8784
rect 14344 -8843 14356 -8837
rect 14536 -8843 14548 -8837
rect 14726 -8837 14780 -8803
rect 15164 -8834 15178 -8680
rect 15236 -8714 15295 -8680
rect 15225 -8753 15239 -8742
rect 15281 -8753 15295 -8742
rect 15236 -8787 15295 -8753
rect 15342 -8834 15356 -8680
rect 15376 -8739 15390 -8676
rect 15392 -8710 15456 -8676
rect 15596 -8680 15607 -8669
rect 15688 -8676 15707 -8668
rect 15749 -8676 15768 -8668
rect 16000 -8668 16014 -8474
rect 16017 -8508 16080 -8474
rect 16066 -8668 16080 -8508
rect 16100 -8230 16114 -8208
rect 16162 -8224 16176 -8216
rect 16218 -8224 16232 -8216
rect 16173 -8230 16232 -8224
rect 16278 -8230 16292 -8208
rect 16100 -8264 16148 -8230
rect 16172 -8258 16232 -8230
rect 16172 -8264 16220 -8258
rect 16244 -8264 16292 -8230
rect 16100 -8524 16114 -8264
rect 16162 -8292 16176 -8281
rect 16218 -8292 16232 -8281
rect 16173 -8326 16232 -8292
rect 16162 -8406 16176 -8395
rect 16218 -8406 16232 -8395
rect 16173 -8440 16232 -8406
rect 16162 -8474 16176 -8463
rect 16218 -8474 16232 -8463
rect 16173 -8508 16232 -8474
rect 16278 -8524 16292 -8264
rect 16312 -8216 16326 -8208
rect 16378 -8216 16392 -8208
rect 16312 -8224 16332 -8216
rect 16374 -8224 16392 -8216
rect 16312 -8281 16326 -8224
rect 16329 -8258 16392 -8224
rect 16378 -8281 16392 -8258
rect 16312 -8292 16332 -8281
rect 16374 -8292 16392 -8281
rect 16312 -8395 16326 -8292
rect 16329 -8326 16392 -8292
rect 16378 -8395 16392 -8326
rect 16312 -8406 16332 -8395
rect 16374 -8406 16392 -8395
rect 16312 -8463 16326 -8406
rect 16329 -8440 16392 -8406
rect 16329 -8463 16377 -8461
rect 16378 -8463 16392 -8440
rect 16312 -8474 16392 -8463
rect 16100 -8646 16114 -8580
rect 16116 -8609 16164 -8596
rect 16229 -8609 16277 -8596
rect 16116 -8630 16185 -8609
rect 16137 -8643 16185 -8630
rect 16209 -8630 16277 -8609
rect 16209 -8643 16257 -8630
rect 16278 -8646 16292 -8580
rect 15442 -8739 15456 -8710
rect 15376 -8750 15395 -8739
rect 15437 -8750 15456 -8739
rect 15376 -8800 15390 -8750
rect 15392 -8784 15456 -8750
rect 15442 -8800 15456 -8784
rect 15476 -8834 15490 -8680
rect 15548 -8714 15607 -8680
rect 15537 -8753 15551 -8742
rect 15593 -8753 15607 -8742
rect 15548 -8787 15607 -8753
rect 15654 -8834 15668 -8680
rect 15688 -8739 15702 -8676
rect 15704 -8710 15768 -8676
rect 15908 -8680 15919 -8669
rect 16000 -8676 16019 -8668
rect 16061 -8676 16080 -8668
rect 16312 -8668 16326 -8474
rect 16329 -8508 16392 -8474
rect 16378 -8668 16392 -8508
rect 16412 -8230 16426 -8208
rect 16474 -8224 16488 -8216
rect 16530 -8224 16544 -8216
rect 16485 -8230 16544 -8224
rect 16590 -8230 16604 -8208
rect 16412 -8264 16460 -8230
rect 16484 -8258 16544 -8230
rect 16484 -8264 16532 -8258
rect 16556 -8264 16604 -8230
rect 16412 -8524 16426 -8264
rect 16474 -8292 16488 -8281
rect 16530 -8292 16544 -8281
rect 16485 -8326 16544 -8292
rect 16474 -8406 16488 -8395
rect 16530 -8406 16544 -8395
rect 16485 -8440 16544 -8406
rect 16474 -8474 16488 -8463
rect 16530 -8474 16544 -8463
rect 16485 -8508 16544 -8474
rect 16590 -8524 16604 -8264
rect 16624 -8216 16638 -8208
rect 16690 -8216 16704 -8208
rect 16624 -8224 16644 -8216
rect 16686 -8224 16704 -8216
rect 16624 -8281 16638 -8224
rect 16641 -8258 16704 -8224
rect 16690 -8281 16704 -8258
rect 16624 -8292 16644 -8281
rect 16686 -8292 16704 -8281
rect 16624 -8395 16638 -8292
rect 16641 -8326 16704 -8292
rect 16690 -8395 16704 -8326
rect 16624 -8406 16644 -8395
rect 16686 -8406 16704 -8395
rect 16624 -8463 16638 -8406
rect 16641 -8440 16704 -8406
rect 16641 -8463 16689 -8461
rect 16690 -8463 16704 -8440
rect 16624 -8474 16704 -8463
rect 16412 -8646 16426 -8580
rect 16428 -8609 16476 -8596
rect 16541 -8609 16589 -8596
rect 16428 -8630 16497 -8609
rect 16449 -8643 16497 -8630
rect 16521 -8630 16589 -8609
rect 16521 -8643 16569 -8630
rect 16590 -8646 16604 -8580
rect 15754 -8739 15768 -8710
rect 15688 -8750 15707 -8739
rect 15749 -8750 15768 -8739
rect 15688 -8800 15702 -8750
rect 15704 -8784 15768 -8750
rect 15754 -8800 15768 -8784
rect 15788 -8834 15802 -8680
rect 15860 -8714 15919 -8680
rect 15849 -8753 15863 -8742
rect 15905 -8753 15919 -8742
rect 15860 -8787 15919 -8753
rect 15966 -8834 15980 -8680
rect 16000 -8739 16014 -8676
rect 16016 -8710 16080 -8676
rect 16220 -8680 16231 -8669
rect 16312 -8676 16331 -8668
rect 16373 -8676 16392 -8668
rect 16624 -8668 16638 -8474
rect 16641 -8508 16704 -8474
rect 16690 -8668 16704 -8508
rect 16724 -8230 16738 -8208
rect 16786 -8224 16800 -8216
rect 16842 -8224 16856 -8216
rect 16797 -8230 16856 -8224
rect 16902 -8230 16916 -8208
rect 16724 -8264 16772 -8230
rect 16796 -8258 16856 -8230
rect 16796 -8264 16844 -8258
rect 16868 -8264 16916 -8230
rect 16724 -8524 16738 -8264
rect 16786 -8292 16800 -8281
rect 16842 -8292 16856 -8281
rect 16797 -8326 16856 -8292
rect 16786 -8406 16800 -8395
rect 16842 -8406 16856 -8395
rect 16797 -8440 16856 -8406
rect 16786 -8474 16800 -8463
rect 16842 -8474 16856 -8463
rect 16797 -8508 16856 -8474
rect 16902 -8524 16916 -8264
rect 16936 -8216 16950 -8208
rect 17002 -8216 17016 -8208
rect 16936 -8224 16956 -8216
rect 16998 -8224 17016 -8216
rect 16936 -8281 16950 -8224
rect 16953 -8258 17016 -8224
rect 17002 -8281 17016 -8258
rect 16936 -8292 16956 -8281
rect 16998 -8292 17016 -8281
rect 16936 -8395 16950 -8292
rect 16953 -8326 17016 -8292
rect 17002 -8395 17016 -8326
rect 16936 -8406 16956 -8395
rect 16998 -8406 17016 -8395
rect 16936 -8463 16950 -8406
rect 16953 -8440 17016 -8406
rect 16953 -8463 17001 -8461
rect 17002 -8463 17016 -8440
rect 16936 -8474 17016 -8463
rect 16724 -8646 16738 -8580
rect 16740 -8609 16788 -8596
rect 16853 -8609 16901 -8596
rect 16740 -8630 16809 -8609
rect 16761 -8643 16809 -8630
rect 16833 -8630 16901 -8609
rect 16833 -8643 16881 -8630
rect 16902 -8646 16916 -8580
rect 16066 -8739 16080 -8710
rect 16000 -8750 16019 -8739
rect 16061 -8750 16080 -8739
rect 16000 -8800 16014 -8750
rect 16016 -8784 16080 -8750
rect 16066 -8800 16080 -8784
rect 16100 -8834 16114 -8680
rect 16172 -8714 16231 -8680
rect 16161 -8753 16175 -8742
rect 16217 -8753 16231 -8742
rect 16172 -8787 16231 -8753
rect 16278 -8834 16292 -8680
rect 16312 -8739 16326 -8676
rect 16328 -8710 16392 -8676
rect 16532 -8680 16543 -8669
rect 16624 -8676 16643 -8668
rect 16685 -8676 16704 -8668
rect 16936 -8668 16950 -8474
rect 16953 -8508 17016 -8474
rect 17002 -8668 17016 -8508
rect 17036 -8230 17050 -8208
rect 17098 -8224 17112 -8216
rect 17154 -8224 17168 -8216
rect 17109 -8230 17168 -8224
rect 17214 -8230 17228 -8208
rect 17036 -8264 17084 -8230
rect 17108 -8258 17168 -8230
rect 17108 -8264 17156 -8258
rect 17180 -8264 17228 -8230
rect 17036 -8524 17050 -8264
rect 17098 -8292 17112 -8281
rect 17154 -8292 17168 -8281
rect 17109 -8326 17168 -8292
rect 17098 -8406 17112 -8395
rect 17154 -8406 17168 -8395
rect 17109 -8440 17168 -8406
rect 17098 -8474 17112 -8463
rect 17154 -8474 17168 -8463
rect 17109 -8508 17168 -8474
rect 17214 -8524 17228 -8264
rect 17248 -8216 17262 -8208
rect 17314 -8216 17328 -8208
rect 17248 -8224 17268 -8216
rect 17310 -8224 17328 -8216
rect 17248 -8281 17262 -8224
rect 17265 -8258 17328 -8224
rect 17314 -8281 17328 -8258
rect 17248 -8292 17268 -8281
rect 17310 -8292 17328 -8281
rect 17248 -8395 17262 -8292
rect 17265 -8326 17328 -8292
rect 17314 -8395 17328 -8326
rect 17248 -8406 17268 -8395
rect 17310 -8406 17328 -8395
rect 17248 -8463 17262 -8406
rect 17265 -8440 17328 -8406
rect 17265 -8463 17313 -8461
rect 17314 -8463 17328 -8440
rect 17248 -8474 17328 -8463
rect 17036 -8646 17050 -8580
rect 17052 -8609 17100 -8596
rect 17165 -8609 17213 -8596
rect 17052 -8630 17121 -8609
rect 17073 -8643 17121 -8630
rect 17145 -8630 17213 -8609
rect 17145 -8643 17193 -8630
rect 17214 -8646 17228 -8580
rect 16378 -8739 16392 -8710
rect 16312 -8750 16331 -8739
rect 16373 -8750 16392 -8739
rect 16312 -8800 16326 -8750
rect 16328 -8784 16392 -8750
rect 16378 -8800 16392 -8784
rect 16412 -8834 16426 -8680
rect 16484 -8714 16543 -8680
rect 16473 -8753 16487 -8742
rect 16529 -8753 16543 -8742
rect 16484 -8787 16543 -8753
rect 16590 -8834 16604 -8680
rect 16624 -8739 16638 -8676
rect 16640 -8710 16704 -8676
rect 16844 -8680 16855 -8669
rect 16936 -8676 16955 -8668
rect 16997 -8676 17016 -8668
rect 17248 -8668 17262 -8474
rect 17265 -8508 17328 -8474
rect 17314 -8558 17328 -8508
rect 17348 -8230 17362 -8224
rect 17410 -8228 17424 -8217
rect 17421 -8230 17469 -8228
rect 17348 -8264 17405 -8230
rect 17421 -8262 17477 -8230
rect 17429 -8264 17477 -8262
rect 17348 -8524 17362 -8264
rect 17410 -8296 17424 -8285
rect 17421 -8330 17469 -8296
rect 17410 -8402 17424 -8391
rect 17421 -8436 17469 -8402
rect 17410 -8470 17424 -8459
rect 17421 -8504 17469 -8470
rect 17314 -8668 17328 -8646
rect 16690 -8739 16704 -8710
rect 16624 -8750 16643 -8739
rect 16685 -8750 16704 -8739
rect 16624 -8800 16638 -8750
rect 16640 -8784 16704 -8750
rect 16690 -8800 16704 -8784
rect 16724 -8834 16738 -8680
rect 16796 -8714 16855 -8680
rect 16785 -8753 16799 -8742
rect 16841 -8753 16855 -8742
rect 16796 -8787 16855 -8753
rect 16902 -8834 16916 -8680
rect 16936 -8739 16950 -8676
rect 16952 -8710 17016 -8676
rect 17156 -8680 17167 -8669
rect 17248 -8676 17267 -8668
rect 17309 -8676 17328 -8668
rect 17002 -8739 17016 -8710
rect 16936 -8750 16955 -8739
rect 16997 -8750 17016 -8739
rect 16936 -8800 16950 -8750
rect 16952 -8784 17016 -8750
rect 17002 -8800 17016 -8784
rect 17036 -8834 17050 -8680
rect 17108 -8714 17167 -8680
rect 17097 -8753 17111 -8742
rect 17153 -8753 17167 -8742
rect 17108 -8787 17167 -8753
rect 17214 -8834 17228 -8680
rect 17248 -8739 17262 -8676
rect 17264 -8710 17328 -8676
rect 17314 -8739 17328 -8710
rect 17248 -8750 17267 -8739
rect 17309 -8750 17328 -8739
rect 17248 -8800 17262 -8750
rect 17264 -8784 17328 -8750
rect 17314 -8800 17328 -8784
rect 17348 -8834 17362 -8680
rect 17420 -8714 17468 -8680
rect 17409 -8753 17423 -8742
rect 17420 -8787 17468 -8753
rect 14726 -8843 14735 -8837
rect 11296 -8890 11298 -8856
rect 11327 -8890 11375 -8856
rect 11423 -8890 11471 -8856
rect 11519 -8890 11567 -8856
rect 11615 -8890 11663 -8856
rect 11711 -8890 11759 -8856
rect 11807 -8890 11855 -8856
rect 11903 -8890 11951 -8856
rect 11999 -8890 12047 -8856
rect 12095 -8890 12143 -8856
rect 12191 -8890 12239 -8856
rect 12287 -8890 12335 -8856
rect 12383 -8890 12431 -8856
rect 12479 -8890 12527 -8856
rect 12575 -8890 12623 -8856
rect 12671 -8890 12719 -8856
rect 12767 -8890 12815 -8856
rect 12863 -8890 12911 -8856
rect 12959 -8890 13007 -8856
rect 13055 -8890 13103 -8856
rect 13151 -8890 13199 -8856
rect 13247 -8890 13295 -8856
rect 13343 -8890 13391 -8856
rect 13439 -8890 13487 -8856
rect 13535 -8890 13583 -8856
rect 13631 -8890 13679 -8856
rect 13727 -8890 13775 -8856
rect 13823 -8890 13871 -8856
rect 13919 -8890 13967 -8856
rect 13996 -8890 13998 -8856
rect 14903 -8874 14951 -8840
rect 14975 -8874 15023 -8840
rect 15164 -8874 15212 -8840
rect 15236 -8874 15284 -8840
rect 15308 -8874 15356 -8840
rect 15476 -8874 15524 -8840
rect 15548 -8874 15596 -8840
rect 15620 -8874 15668 -8840
rect 15788 -8874 15836 -8840
rect 15860 -8874 15908 -8840
rect 15932 -8874 15980 -8840
rect 16100 -8874 16148 -8840
rect 16172 -8874 16220 -8840
rect 16244 -8874 16292 -8840
rect 16412 -8874 16460 -8840
rect 16484 -8874 16532 -8840
rect 16556 -8874 16604 -8840
rect 16724 -8874 16772 -8840
rect 16796 -8874 16844 -8840
rect 16868 -8874 16916 -8840
rect 17036 -8874 17084 -8840
rect 17108 -8874 17156 -8840
rect 17180 -8874 17228 -8840
rect 17357 -8874 17405 -8840
rect 17429 -8874 17477 -8840
rect 14050 -8933 14052 -8899
rect 14081 -8933 14129 -8899
rect 14177 -8933 14225 -8899
rect 14273 -8933 14321 -8899
rect 14369 -8933 14417 -8899
rect 14465 -8933 14513 -8899
rect 14561 -8933 14609 -8899
rect 14657 -8933 14705 -8899
rect 14753 -8933 14801 -8899
rect 14830 -8933 14832 -8899
rect 14884 -8976 14886 -8942
rect 14915 -8976 14963 -8942
rect 15011 -8976 15059 -8942
rect 15107 -8976 15155 -8942
rect 15203 -8976 15251 -8942
rect 15299 -8976 15347 -8942
rect 15395 -8976 15443 -8942
rect 15491 -8976 15539 -8942
rect 15587 -8976 15635 -8942
rect 15683 -8976 15731 -8942
rect 15779 -8976 15827 -8942
rect 15875 -8976 15923 -8942
rect 15971 -8976 16019 -8942
rect 16067 -8976 16115 -8942
rect 16163 -8976 16211 -8942
rect 16259 -8976 16307 -8942
rect 16355 -8976 16403 -8942
rect 16451 -8976 16499 -8942
rect 16547 -8976 16595 -8942
rect 16643 -8976 16691 -8942
rect 16739 -8976 16787 -8942
rect 16835 -8976 16883 -8942
rect 16931 -8976 16979 -8942
rect 17027 -8976 17075 -8942
rect 17123 -8976 17171 -8942
rect 17219 -8976 17267 -8942
rect 17315 -8976 17363 -8942
rect 17411 -8976 17459 -8942
rect 17507 -8976 17555 -8942
rect 3810 -11153 5717 -11123
rect 3811 -11188 5717 -11153
rect 4401 -11248 5717 -11188
rect 4432 -11253 5717 -11248
rect 4570 -11271 5717 -11253
rect 4992 -11282 5717 -11271
rect 4992 -11318 5680 -11282
rect 5191 -11336 5680 -11318
rect 5227 -11360 5609 -11336
rect 2423 -17666 2461 -17641
rect 4889 -17709 4927 -17684
rect 7355 -17752 7393 -17727
rect 9821 -17795 9859 -17770
rect 12287 -17838 12325 -17813
rect 14753 -17881 14791 -17856
rect 17219 -17924 17257 -17899
rect 19685 -17952 19723 -17942
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
use p_ibias_mirror  x1
timestamp 1717439242
transform 1 0 5 0 1 -4800
box -95 -2270 7078 1109
use n_ibias_mirror  x2
timestamp 1717439242
transform 1 0 6 0 1 -4800
box -65 -1985 4815 721
use icell256_unary_scs  x3
timestamp 1717439242
transform 1 0 8 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x4
timestamp 1717439242
transform 1 0 9 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x5
timestamp 1717439242
transform 1 0 10 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x6
timestamp 1717439242
transform 1 0 11 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x7
timestamp 1717439242
transform 1 0 12 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x8
timestamp 1717439242
transform 1 0 13 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x9
timestamp 1717439242
transform 1 0 14 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x10
timestamp 1717439242
transform 1 0 15 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x11
timestamp 1717439242
transform 1 0 16 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x12
timestamp 1717439242
transform 1 0 17 0 1 -4800
box -66 -6638 17630 668726
use lvhvbuffc  x13
timestamp 1717439242
transform 1 0 0 0 1 -4800
box -66 -2172 6024 200
use icell256_unary_scs  x14
timestamp 1717439242
transform 1 0 18 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x15
timestamp 1717439242
transform 1 0 19 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x16
timestamp 1717439242
transform 1 0 20 0 1 -4800
box -66 -6638 17630 668726
use bin2thermo4bit_0_15  x17
timestamp 1717439242
transform 1 0 4 0 1 -4800
box -66 -11892 33912 200
use mosgsconnected  x18
timestamp 1717439242
transform 1 0 7 0 1 -4800
box -95 -495 621 2499
use icell256_unary_scs  x19
timestamp 1717439242
transform 1 0 21 0 1 -4800
box -66 -6638 17630 668726
use icell256_unary_scs  x20
timestamp 1717439242
transform 1 0 22 0 1 -4800
box -66 -6638 17630 668726
use dff15ch  x21
timestamp 1717439242
transform 1 0 23 0 1 -4800
box -66 -13845 36990 200
use lvhvbuffc  x66
timestamp 1717439242
transform 1 0 1 0 1 -4800
box -66 -2172 6024 200
use lvhvbuffc  x67
timestamp 1717439242
transform 1 0 2 0 1 -4800
box -66 -2172 6024 200
use lvhvbuffc  x68
timestamp 1717439242
transform 1 0 3 0 1 -4800
box -66 -2172 6024 200
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 dvdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 iout
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 avdd
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 dvss
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 avss
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 dlv0
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 dlv1
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 dlv2
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 dlv3
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 clk
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 iref
port 12 nsew
<< end >>
