magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< nwell >>
rect -358 -337587 358 337587
<< mvpmos >>
rect -100 334890 100 337290
rect -100 332254 100 334654
rect -100 329618 100 332018
rect -100 326982 100 329382
rect -100 324346 100 326746
rect -100 321710 100 324110
rect -100 319074 100 321474
rect -100 316438 100 318838
rect -100 313802 100 316202
rect -100 311166 100 313566
rect -100 308530 100 310930
rect -100 305894 100 308294
rect -100 303258 100 305658
rect -100 300622 100 303022
rect -100 297986 100 300386
rect -100 295350 100 297750
rect -100 292714 100 295114
rect -100 290078 100 292478
rect -100 287442 100 289842
rect -100 284806 100 287206
rect -100 282170 100 284570
rect -100 279534 100 281934
rect -100 276898 100 279298
rect -100 274262 100 276662
rect -100 271626 100 274026
rect -100 268990 100 271390
rect -100 266354 100 268754
rect -100 263718 100 266118
rect -100 261082 100 263482
rect -100 258446 100 260846
rect -100 255810 100 258210
rect -100 253174 100 255574
rect -100 250538 100 252938
rect -100 247902 100 250302
rect -100 245266 100 247666
rect -100 242630 100 245030
rect -100 239994 100 242394
rect -100 237358 100 239758
rect -100 234722 100 237122
rect -100 232086 100 234486
rect -100 229450 100 231850
rect -100 226814 100 229214
rect -100 224178 100 226578
rect -100 221542 100 223942
rect -100 218906 100 221306
rect -100 216270 100 218670
rect -100 213634 100 216034
rect -100 210998 100 213398
rect -100 208362 100 210762
rect -100 205726 100 208126
rect -100 203090 100 205490
rect -100 200454 100 202854
rect -100 197818 100 200218
rect -100 195182 100 197582
rect -100 192546 100 194946
rect -100 189910 100 192310
rect -100 187274 100 189674
rect -100 184638 100 187038
rect -100 182002 100 184402
rect -100 179366 100 181766
rect -100 176730 100 179130
rect -100 174094 100 176494
rect -100 171458 100 173858
rect -100 168822 100 171222
rect -100 166186 100 168586
rect -100 163550 100 165950
rect -100 160914 100 163314
rect -100 158278 100 160678
rect -100 155642 100 158042
rect -100 153006 100 155406
rect -100 150370 100 152770
rect -100 147734 100 150134
rect -100 145098 100 147498
rect -100 142462 100 144862
rect -100 139826 100 142226
rect -100 137190 100 139590
rect -100 134554 100 136954
rect -100 131918 100 134318
rect -100 129282 100 131682
rect -100 126646 100 129046
rect -100 124010 100 126410
rect -100 121374 100 123774
rect -100 118738 100 121138
rect -100 116102 100 118502
rect -100 113466 100 115866
rect -100 110830 100 113230
rect -100 108194 100 110594
rect -100 105558 100 107958
rect -100 102922 100 105322
rect -100 100286 100 102686
rect -100 97650 100 100050
rect -100 95014 100 97414
rect -100 92378 100 94778
rect -100 89742 100 92142
rect -100 87106 100 89506
rect -100 84470 100 86870
rect -100 81834 100 84234
rect -100 79198 100 81598
rect -100 76562 100 78962
rect -100 73926 100 76326
rect -100 71290 100 73690
rect -100 68654 100 71054
rect -100 66018 100 68418
rect -100 63382 100 65782
rect -100 60746 100 63146
rect -100 58110 100 60510
rect -100 55474 100 57874
rect -100 52838 100 55238
rect -100 50202 100 52602
rect -100 47566 100 49966
rect -100 44930 100 47330
rect -100 42294 100 44694
rect -100 39658 100 42058
rect -100 37022 100 39422
rect -100 34386 100 36786
rect -100 31750 100 34150
rect -100 29114 100 31514
rect -100 26478 100 28878
rect -100 23842 100 26242
rect -100 21206 100 23606
rect -100 18570 100 20970
rect -100 15934 100 18334
rect -100 13298 100 15698
rect -100 10662 100 13062
rect -100 8026 100 10426
rect -100 5390 100 7790
rect -100 2754 100 5154
rect -100 118 100 2518
rect -100 -2518 100 -118
rect -100 -5154 100 -2754
rect -100 -7790 100 -5390
rect -100 -10426 100 -8026
rect -100 -13062 100 -10662
rect -100 -15698 100 -13298
rect -100 -18334 100 -15934
rect -100 -20970 100 -18570
rect -100 -23606 100 -21206
rect -100 -26242 100 -23842
rect -100 -28878 100 -26478
rect -100 -31514 100 -29114
rect -100 -34150 100 -31750
rect -100 -36786 100 -34386
rect -100 -39422 100 -37022
rect -100 -42058 100 -39658
rect -100 -44694 100 -42294
rect -100 -47330 100 -44930
rect -100 -49966 100 -47566
rect -100 -52602 100 -50202
rect -100 -55238 100 -52838
rect -100 -57874 100 -55474
rect -100 -60510 100 -58110
rect -100 -63146 100 -60746
rect -100 -65782 100 -63382
rect -100 -68418 100 -66018
rect -100 -71054 100 -68654
rect -100 -73690 100 -71290
rect -100 -76326 100 -73926
rect -100 -78962 100 -76562
rect -100 -81598 100 -79198
rect -100 -84234 100 -81834
rect -100 -86870 100 -84470
rect -100 -89506 100 -87106
rect -100 -92142 100 -89742
rect -100 -94778 100 -92378
rect -100 -97414 100 -95014
rect -100 -100050 100 -97650
rect -100 -102686 100 -100286
rect -100 -105322 100 -102922
rect -100 -107958 100 -105558
rect -100 -110594 100 -108194
rect -100 -113230 100 -110830
rect -100 -115866 100 -113466
rect -100 -118502 100 -116102
rect -100 -121138 100 -118738
rect -100 -123774 100 -121374
rect -100 -126410 100 -124010
rect -100 -129046 100 -126646
rect -100 -131682 100 -129282
rect -100 -134318 100 -131918
rect -100 -136954 100 -134554
rect -100 -139590 100 -137190
rect -100 -142226 100 -139826
rect -100 -144862 100 -142462
rect -100 -147498 100 -145098
rect -100 -150134 100 -147734
rect -100 -152770 100 -150370
rect -100 -155406 100 -153006
rect -100 -158042 100 -155642
rect -100 -160678 100 -158278
rect -100 -163314 100 -160914
rect -100 -165950 100 -163550
rect -100 -168586 100 -166186
rect -100 -171222 100 -168822
rect -100 -173858 100 -171458
rect -100 -176494 100 -174094
rect -100 -179130 100 -176730
rect -100 -181766 100 -179366
rect -100 -184402 100 -182002
rect -100 -187038 100 -184638
rect -100 -189674 100 -187274
rect -100 -192310 100 -189910
rect -100 -194946 100 -192546
rect -100 -197582 100 -195182
rect -100 -200218 100 -197818
rect -100 -202854 100 -200454
rect -100 -205490 100 -203090
rect -100 -208126 100 -205726
rect -100 -210762 100 -208362
rect -100 -213398 100 -210998
rect -100 -216034 100 -213634
rect -100 -218670 100 -216270
rect -100 -221306 100 -218906
rect -100 -223942 100 -221542
rect -100 -226578 100 -224178
rect -100 -229214 100 -226814
rect -100 -231850 100 -229450
rect -100 -234486 100 -232086
rect -100 -237122 100 -234722
rect -100 -239758 100 -237358
rect -100 -242394 100 -239994
rect -100 -245030 100 -242630
rect -100 -247666 100 -245266
rect -100 -250302 100 -247902
rect -100 -252938 100 -250538
rect -100 -255574 100 -253174
rect -100 -258210 100 -255810
rect -100 -260846 100 -258446
rect -100 -263482 100 -261082
rect -100 -266118 100 -263718
rect -100 -268754 100 -266354
rect -100 -271390 100 -268990
rect -100 -274026 100 -271626
rect -100 -276662 100 -274262
rect -100 -279298 100 -276898
rect -100 -281934 100 -279534
rect -100 -284570 100 -282170
rect -100 -287206 100 -284806
rect -100 -289842 100 -287442
rect -100 -292478 100 -290078
rect -100 -295114 100 -292714
rect -100 -297750 100 -295350
rect -100 -300386 100 -297986
rect -100 -303022 100 -300622
rect -100 -305658 100 -303258
rect -100 -308294 100 -305894
rect -100 -310930 100 -308530
rect -100 -313566 100 -311166
rect -100 -316202 100 -313802
rect -100 -318838 100 -316438
rect -100 -321474 100 -319074
rect -100 -324110 100 -321710
rect -100 -326746 100 -324346
rect -100 -329382 100 -326982
rect -100 -332018 100 -329618
rect -100 -334654 100 -332254
rect -100 -337290 100 -334890
<< mvpdiff >>
rect -158 337278 -100 337290
rect -158 334902 -146 337278
rect -112 334902 -100 337278
rect -158 334890 -100 334902
rect 100 337278 158 337290
rect 100 334902 112 337278
rect 146 334902 158 337278
rect 100 334890 158 334902
rect -158 334642 -100 334654
rect -158 332266 -146 334642
rect -112 332266 -100 334642
rect -158 332254 -100 332266
rect 100 334642 158 334654
rect 100 332266 112 334642
rect 146 332266 158 334642
rect 100 332254 158 332266
rect -158 332006 -100 332018
rect -158 329630 -146 332006
rect -112 329630 -100 332006
rect -158 329618 -100 329630
rect 100 332006 158 332018
rect 100 329630 112 332006
rect 146 329630 158 332006
rect 100 329618 158 329630
rect -158 329370 -100 329382
rect -158 326994 -146 329370
rect -112 326994 -100 329370
rect -158 326982 -100 326994
rect 100 329370 158 329382
rect 100 326994 112 329370
rect 146 326994 158 329370
rect 100 326982 158 326994
rect -158 326734 -100 326746
rect -158 324358 -146 326734
rect -112 324358 -100 326734
rect -158 324346 -100 324358
rect 100 326734 158 326746
rect 100 324358 112 326734
rect 146 324358 158 326734
rect 100 324346 158 324358
rect -158 324098 -100 324110
rect -158 321722 -146 324098
rect -112 321722 -100 324098
rect -158 321710 -100 321722
rect 100 324098 158 324110
rect 100 321722 112 324098
rect 146 321722 158 324098
rect 100 321710 158 321722
rect -158 321462 -100 321474
rect -158 319086 -146 321462
rect -112 319086 -100 321462
rect -158 319074 -100 319086
rect 100 321462 158 321474
rect 100 319086 112 321462
rect 146 319086 158 321462
rect 100 319074 158 319086
rect -158 318826 -100 318838
rect -158 316450 -146 318826
rect -112 316450 -100 318826
rect -158 316438 -100 316450
rect 100 318826 158 318838
rect 100 316450 112 318826
rect 146 316450 158 318826
rect 100 316438 158 316450
rect -158 316190 -100 316202
rect -158 313814 -146 316190
rect -112 313814 -100 316190
rect -158 313802 -100 313814
rect 100 316190 158 316202
rect 100 313814 112 316190
rect 146 313814 158 316190
rect 100 313802 158 313814
rect -158 313554 -100 313566
rect -158 311178 -146 313554
rect -112 311178 -100 313554
rect -158 311166 -100 311178
rect 100 313554 158 313566
rect 100 311178 112 313554
rect 146 311178 158 313554
rect 100 311166 158 311178
rect -158 310918 -100 310930
rect -158 308542 -146 310918
rect -112 308542 -100 310918
rect -158 308530 -100 308542
rect 100 310918 158 310930
rect 100 308542 112 310918
rect 146 308542 158 310918
rect 100 308530 158 308542
rect -158 308282 -100 308294
rect -158 305906 -146 308282
rect -112 305906 -100 308282
rect -158 305894 -100 305906
rect 100 308282 158 308294
rect 100 305906 112 308282
rect 146 305906 158 308282
rect 100 305894 158 305906
rect -158 305646 -100 305658
rect -158 303270 -146 305646
rect -112 303270 -100 305646
rect -158 303258 -100 303270
rect 100 305646 158 305658
rect 100 303270 112 305646
rect 146 303270 158 305646
rect 100 303258 158 303270
rect -158 303010 -100 303022
rect -158 300634 -146 303010
rect -112 300634 -100 303010
rect -158 300622 -100 300634
rect 100 303010 158 303022
rect 100 300634 112 303010
rect 146 300634 158 303010
rect 100 300622 158 300634
rect -158 300374 -100 300386
rect -158 297998 -146 300374
rect -112 297998 -100 300374
rect -158 297986 -100 297998
rect 100 300374 158 300386
rect 100 297998 112 300374
rect 146 297998 158 300374
rect 100 297986 158 297998
rect -158 297738 -100 297750
rect -158 295362 -146 297738
rect -112 295362 -100 297738
rect -158 295350 -100 295362
rect 100 297738 158 297750
rect 100 295362 112 297738
rect 146 295362 158 297738
rect 100 295350 158 295362
rect -158 295102 -100 295114
rect -158 292726 -146 295102
rect -112 292726 -100 295102
rect -158 292714 -100 292726
rect 100 295102 158 295114
rect 100 292726 112 295102
rect 146 292726 158 295102
rect 100 292714 158 292726
rect -158 292466 -100 292478
rect -158 290090 -146 292466
rect -112 290090 -100 292466
rect -158 290078 -100 290090
rect 100 292466 158 292478
rect 100 290090 112 292466
rect 146 290090 158 292466
rect 100 290078 158 290090
rect -158 289830 -100 289842
rect -158 287454 -146 289830
rect -112 287454 -100 289830
rect -158 287442 -100 287454
rect 100 289830 158 289842
rect 100 287454 112 289830
rect 146 287454 158 289830
rect 100 287442 158 287454
rect -158 287194 -100 287206
rect -158 284818 -146 287194
rect -112 284818 -100 287194
rect -158 284806 -100 284818
rect 100 287194 158 287206
rect 100 284818 112 287194
rect 146 284818 158 287194
rect 100 284806 158 284818
rect -158 284558 -100 284570
rect -158 282182 -146 284558
rect -112 282182 -100 284558
rect -158 282170 -100 282182
rect 100 284558 158 284570
rect 100 282182 112 284558
rect 146 282182 158 284558
rect 100 282170 158 282182
rect -158 281922 -100 281934
rect -158 279546 -146 281922
rect -112 279546 -100 281922
rect -158 279534 -100 279546
rect 100 281922 158 281934
rect 100 279546 112 281922
rect 146 279546 158 281922
rect 100 279534 158 279546
rect -158 279286 -100 279298
rect -158 276910 -146 279286
rect -112 276910 -100 279286
rect -158 276898 -100 276910
rect 100 279286 158 279298
rect 100 276910 112 279286
rect 146 276910 158 279286
rect 100 276898 158 276910
rect -158 276650 -100 276662
rect -158 274274 -146 276650
rect -112 274274 -100 276650
rect -158 274262 -100 274274
rect 100 276650 158 276662
rect 100 274274 112 276650
rect 146 274274 158 276650
rect 100 274262 158 274274
rect -158 274014 -100 274026
rect -158 271638 -146 274014
rect -112 271638 -100 274014
rect -158 271626 -100 271638
rect 100 274014 158 274026
rect 100 271638 112 274014
rect 146 271638 158 274014
rect 100 271626 158 271638
rect -158 271378 -100 271390
rect -158 269002 -146 271378
rect -112 269002 -100 271378
rect -158 268990 -100 269002
rect 100 271378 158 271390
rect 100 269002 112 271378
rect 146 269002 158 271378
rect 100 268990 158 269002
rect -158 268742 -100 268754
rect -158 266366 -146 268742
rect -112 266366 -100 268742
rect -158 266354 -100 266366
rect 100 268742 158 268754
rect 100 266366 112 268742
rect 146 266366 158 268742
rect 100 266354 158 266366
rect -158 266106 -100 266118
rect -158 263730 -146 266106
rect -112 263730 -100 266106
rect -158 263718 -100 263730
rect 100 266106 158 266118
rect 100 263730 112 266106
rect 146 263730 158 266106
rect 100 263718 158 263730
rect -158 263470 -100 263482
rect -158 261094 -146 263470
rect -112 261094 -100 263470
rect -158 261082 -100 261094
rect 100 263470 158 263482
rect 100 261094 112 263470
rect 146 261094 158 263470
rect 100 261082 158 261094
rect -158 260834 -100 260846
rect -158 258458 -146 260834
rect -112 258458 -100 260834
rect -158 258446 -100 258458
rect 100 260834 158 260846
rect 100 258458 112 260834
rect 146 258458 158 260834
rect 100 258446 158 258458
rect -158 258198 -100 258210
rect -158 255822 -146 258198
rect -112 255822 -100 258198
rect -158 255810 -100 255822
rect 100 258198 158 258210
rect 100 255822 112 258198
rect 146 255822 158 258198
rect 100 255810 158 255822
rect -158 255562 -100 255574
rect -158 253186 -146 255562
rect -112 253186 -100 255562
rect -158 253174 -100 253186
rect 100 255562 158 255574
rect 100 253186 112 255562
rect 146 253186 158 255562
rect 100 253174 158 253186
rect -158 252926 -100 252938
rect -158 250550 -146 252926
rect -112 250550 -100 252926
rect -158 250538 -100 250550
rect 100 252926 158 252938
rect 100 250550 112 252926
rect 146 250550 158 252926
rect 100 250538 158 250550
rect -158 250290 -100 250302
rect -158 247914 -146 250290
rect -112 247914 -100 250290
rect -158 247902 -100 247914
rect 100 250290 158 250302
rect 100 247914 112 250290
rect 146 247914 158 250290
rect 100 247902 158 247914
rect -158 247654 -100 247666
rect -158 245278 -146 247654
rect -112 245278 -100 247654
rect -158 245266 -100 245278
rect 100 247654 158 247666
rect 100 245278 112 247654
rect 146 245278 158 247654
rect 100 245266 158 245278
rect -158 245018 -100 245030
rect -158 242642 -146 245018
rect -112 242642 -100 245018
rect -158 242630 -100 242642
rect 100 245018 158 245030
rect 100 242642 112 245018
rect 146 242642 158 245018
rect 100 242630 158 242642
rect -158 242382 -100 242394
rect -158 240006 -146 242382
rect -112 240006 -100 242382
rect -158 239994 -100 240006
rect 100 242382 158 242394
rect 100 240006 112 242382
rect 146 240006 158 242382
rect 100 239994 158 240006
rect -158 239746 -100 239758
rect -158 237370 -146 239746
rect -112 237370 -100 239746
rect -158 237358 -100 237370
rect 100 239746 158 239758
rect 100 237370 112 239746
rect 146 237370 158 239746
rect 100 237358 158 237370
rect -158 237110 -100 237122
rect -158 234734 -146 237110
rect -112 234734 -100 237110
rect -158 234722 -100 234734
rect 100 237110 158 237122
rect 100 234734 112 237110
rect 146 234734 158 237110
rect 100 234722 158 234734
rect -158 234474 -100 234486
rect -158 232098 -146 234474
rect -112 232098 -100 234474
rect -158 232086 -100 232098
rect 100 234474 158 234486
rect 100 232098 112 234474
rect 146 232098 158 234474
rect 100 232086 158 232098
rect -158 231838 -100 231850
rect -158 229462 -146 231838
rect -112 229462 -100 231838
rect -158 229450 -100 229462
rect 100 231838 158 231850
rect 100 229462 112 231838
rect 146 229462 158 231838
rect 100 229450 158 229462
rect -158 229202 -100 229214
rect -158 226826 -146 229202
rect -112 226826 -100 229202
rect -158 226814 -100 226826
rect 100 229202 158 229214
rect 100 226826 112 229202
rect 146 226826 158 229202
rect 100 226814 158 226826
rect -158 226566 -100 226578
rect -158 224190 -146 226566
rect -112 224190 -100 226566
rect -158 224178 -100 224190
rect 100 226566 158 226578
rect 100 224190 112 226566
rect 146 224190 158 226566
rect 100 224178 158 224190
rect -158 223930 -100 223942
rect -158 221554 -146 223930
rect -112 221554 -100 223930
rect -158 221542 -100 221554
rect 100 223930 158 223942
rect 100 221554 112 223930
rect 146 221554 158 223930
rect 100 221542 158 221554
rect -158 221294 -100 221306
rect -158 218918 -146 221294
rect -112 218918 -100 221294
rect -158 218906 -100 218918
rect 100 221294 158 221306
rect 100 218918 112 221294
rect 146 218918 158 221294
rect 100 218906 158 218918
rect -158 218658 -100 218670
rect -158 216282 -146 218658
rect -112 216282 -100 218658
rect -158 216270 -100 216282
rect 100 218658 158 218670
rect 100 216282 112 218658
rect 146 216282 158 218658
rect 100 216270 158 216282
rect -158 216022 -100 216034
rect -158 213646 -146 216022
rect -112 213646 -100 216022
rect -158 213634 -100 213646
rect 100 216022 158 216034
rect 100 213646 112 216022
rect 146 213646 158 216022
rect 100 213634 158 213646
rect -158 213386 -100 213398
rect -158 211010 -146 213386
rect -112 211010 -100 213386
rect -158 210998 -100 211010
rect 100 213386 158 213398
rect 100 211010 112 213386
rect 146 211010 158 213386
rect 100 210998 158 211010
rect -158 210750 -100 210762
rect -158 208374 -146 210750
rect -112 208374 -100 210750
rect -158 208362 -100 208374
rect 100 210750 158 210762
rect 100 208374 112 210750
rect 146 208374 158 210750
rect 100 208362 158 208374
rect -158 208114 -100 208126
rect -158 205738 -146 208114
rect -112 205738 -100 208114
rect -158 205726 -100 205738
rect 100 208114 158 208126
rect 100 205738 112 208114
rect 146 205738 158 208114
rect 100 205726 158 205738
rect -158 205478 -100 205490
rect -158 203102 -146 205478
rect -112 203102 -100 205478
rect -158 203090 -100 203102
rect 100 205478 158 205490
rect 100 203102 112 205478
rect 146 203102 158 205478
rect 100 203090 158 203102
rect -158 202842 -100 202854
rect -158 200466 -146 202842
rect -112 200466 -100 202842
rect -158 200454 -100 200466
rect 100 202842 158 202854
rect 100 200466 112 202842
rect 146 200466 158 202842
rect 100 200454 158 200466
rect -158 200206 -100 200218
rect -158 197830 -146 200206
rect -112 197830 -100 200206
rect -158 197818 -100 197830
rect 100 200206 158 200218
rect 100 197830 112 200206
rect 146 197830 158 200206
rect 100 197818 158 197830
rect -158 197570 -100 197582
rect -158 195194 -146 197570
rect -112 195194 -100 197570
rect -158 195182 -100 195194
rect 100 197570 158 197582
rect 100 195194 112 197570
rect 146 195194 158 197570
rect 100 195182 158 195194
rect -158 194934 -100 194946
rect -158 192558 -146 194934
rect -112 192558 -100 194934
rect -158 192546 -100 192558
rect 100 194934 158 194946
rect 100 192558 112 194934
rect 146 192558 158 194934
rect 100 192546 158 192558
rect -158 192298 -100 192310
rect -158 189922 -146 192298
rect -112 189922 -100 192298
rect -158 189910 -100 189922
rect 100 192298 158 192310
rect 100 189922 112 192298
rect 146 189922 158 192298
rect 100 189910 158 189922
rect -158 189662 -100 189674
rect -158 187286 -146 189662
rect -112 187286 -100 189662
rect -158 187274 -100 187286
rect 100 189662 158 189674
rect 100 187286 112 189662
rect 146 187286 158 189662
rect 100 187274 158 187286
rect -158 187026 -100 187038
rect -158 184650 -146 187026
rect -112 184650 -100 187026
rect -158 184638 -100 184650
rect 100 187026 158 187038
rect 100 184650 112 187026
rect 146 184650 158 187026
rect 100 184638 158 184650
rect -158 184390 -100 184402
rect -158 182014 -146 184390
rect -112 182014 -100 184390
rect -158 182002 -100 182014
rect 100 184390 158 184402
rect 100 182014 112 184390
rect 146 182014 158 184390
rect 100 182002 158 182014
rect -158 181754 -100 181766
rect -158 179378 -146 181754
rect -112 179378 -100 181754
rect -158 179366 -100 179378
rect 100 181754 158 181766
rect 100 179378 112 181754
rect 146 179378 158 181754
rect 100 179366 158 179378
rect -158 179118 -100 179130
rect -158 176742 -146 179118
rect -112 176742 -100 179118
rect -158 176730 -100 176742
rect 100 179118 158 179130
rect 100 176742 112 179118
rect 146 176742 158 179118
rect 100 176730 158 176742
rect -158 176482 -100 176494
rect -158 174106 -146 176482
rect -112 174106 -100 176482
rect -158 174094 -100 174106
rect 100 176482 158 176494
rect 100 174106 112 176482
rect 146 174106 158 176482
rect 100 174094 158 174106
rect -158 173846 -100 173858
rect -158 171470 -146 173846
rect -112 171470 -100 173846
rect -158 171458 -100 171470
rect 100 173846 158 173858
rect 100 171470 112 173846
rect 146 171470 158 173846
rect 100 171458 158 171470
rect -158 171210 -100 171222
rect -158 168834 -146 171210
rect -112 168834 -100 171210
rect -158 168822 -100 168834
rect 100 171210 158 171222
rect 100 168834 112 171210
rect 146 168834 158 171210
rect 100 168822 158 168834
rect -158 168574 -100 168586
rect -158 166198 -146 168574
rect -112 166198 -100 168574
rect -158 166186 -100 166198
rect 100 168574 158 168586
rect 100 166198 112 168574
rect 146 166198 158 168574
rect 100 166186 158 166198
rect -158 165938 -100 165950
rect -158 163562 -146 165938
rect -112 163562 -100 165938
rect -158 163550 -100 163562
rect 100 165938 158 165950
rect 100 163562 112 165938
rect 146 163562 158 165938
rect 100 163550 158 163562
rect -158 163302 -100 163314
rect -158 160926 -146 163302
rect -112 160926 -100 163302
rect -158 160914 -100 160926
rect 100 163302 158 163314
rect 100 160926 112 163302
rect 146 160926 158 163302
rect 100 160914 158 160926
rect -158 160666 -100 160678
rect -158 158290 -146 160666
rect -112 158290 -100 160666
rect -158 158278 -100 158290
rect 100 160666 158 160678
rect 100 158290 112 160666
rect 146 158290 158 160666
rect 100 158278 158 158290
rect -158 158030 -100 158042
rect -158 155654 -146 158030
rect -112 155654 -100 158030
rect -158 155642 -100 155654
rect 100 158030 158 158042
rect 100 155654 112 158030
rect 146 155654 158 158030
rect 100 155642 158 155654
rect -158 155394 -100 155406
rect -158 153018 -146 155394
rect -112 153018 -100 155394
rect -158 153006 -100 153018
rect 100 155394 158 155406
rect 100 153018 112 155394
rect 146 153018 158 155394
rect 100 153006 158 153018
rect -158 152758 -100 152770
rect -158 150382 -146 152758
rect -112 150382 -100 152758
rect -158 150370 -100 150382
rect 100 152758 158 152770
rect 100 150382 112 152758
rect 146 150382 158 152758
rect 100 150370 158 150382
rect -158 150122 -100 150134
rect -158 147746 -146 150122
rect -112 147746 -100 150122
rect -158 147734 -100 147746
rect 100 150122 158 150134
rect 100 147746 112 150122
rect 146 147746 158 150122
rect 100 147734 158 147746
rect -158 147486 -100 147498
rect -158 145110 -146 147486
rect -112 145110 -100 147486
rect -158 145098 -100 145110
rect 100 147486 158 147498
rect 100 145110 112 147486
rect 146 145110 158 147486
rect 100 145098 158 145110
rect -158 144850 -100 144862
rect -158 142474 -146 144850
rect -112 142474 -100 144850
rect -158 142462 -100 142474
rect 100 144850 158 144862
rect 100 142474 112 144850
rect 146 142474 158 144850
rect 100 142462 158 142474
rect -158 142214 -100 142226
rect -158 139838 -146 142214
rect -112 139838 -100 142214
rect -158 139826 -100 139838
rect 100 142214 158 142226
rect 100 139838 112 142214
rect 146 139838 158 142214
rect 100 139826 158 139838
rect -158 139578 -100 139590
rect -158 137202 -146 139578
rect -112 137202 -100 139578
rect -158 137190 -100 137202
rect 100 139578 158 139590
rect 100 137202 112 139578
rect 146 137202 158 139578
rect 100 137190 158 137202
rect -158 136942 -100 136954
rect -158 134566 -146 136942
rect -112 134566 -100 136942
rect -158 134554 -100 134566
rect 100 136942 158 136954
rect 100 134566 112 136942
rect 146 134566 158 136942
rect 100 134554 158 134566
rect -158 134306 -100 134318
rect -158 131930 -146 134306
rect -112 131930 -100 134306
rect -158 131918 -100 131930
rect 100 134306 158 134318
rect 100 131930 112 134306
rect 146 131930 158 134306
rect 100 131918 158 131930
rect -158 131670 -100 131682
rect -158 129294 -146 131670
rect -112 129294 -100 131670
rect -158 129282 -100 129294
rect 100 131670 158 131682
rect 100 129294 112 131670
rect 146 129294 158 131670
rect 100 129282 158 129294
rect -158 129034 -100 129046
rect -158 126658 -146 129034
rect -112 126658 -100 129034
rect -158 126646 -100 126658
rect 100 129034 158 129046
rect 100 126658 112 129034
rect 146 126658 158 129034
rect 100 126646 158 126658
rect -158 126398 -100 126410
rect -158 124022 -146 126398
rect -112 124022 -100 126398
rect -158 124010 -100 124022
rect 100 126398 158 126410
rect 100 124022 112 126398
rect 146 124022 158 126398
rect 100 124010 158 124022
rect -158 123762 -100 123774
rect -158 121386 -146 123762
rect -112 121386 -100 123762
rect -158 121374 -100 121386
rect 100 123762 158 123774
rect 100 121386 112 123762
rect 146 121386 158 123762
rect 100 121374 158 121386
rect -158 121126 -100 121138
rect -158 118750 -146 121126
rect -112 118750 -100 121126
rect -158 118738 -100 118750
rect 100 121126 158 121138
rect 100 118750 112 121126
rect 146 118750 158 121126
rect 100 118738 158 118750
rect -158 118490 -100 118502
rect -158 116114 -146 118490
rect -112 116114 -100 118490
rect -158 116102 -100 116114
rect 100 118490 158 118502
rect 100 116114 112 118490
rect 146 116114 158 118490
rect 100 116102 158 116114
rect -158 115854 -100 115866
rect -158 113478 -146 115854
rect -112 113478 -100 115854
rect -158 113466 -100 113478
rect 100 115854 158 115866
rect 100 113478 112 115854
rect 146 113478 158 115854
rect 100 113466 158 113478
rect -158 113218 -100 113230
rect -158 110842 -146 113218
rect -112 110842 -100 113218
rect -158 110830 -100 110842
rect 100 113218 158 113230
rect 100 110842 112 113218
rect 146 110842 158 113218
rect 100 110830 158 110842
rect -158 110582 -100 110594
rect -158 108206 -146 110582
rect -112 108206 -100 110582
rect -158 108194 -100 108206
rect 100 110582 158 110594
rect 100 108206 112 110582
rect 146 108206 158 110582
rect 100 108194 158 108206
rect -158 107946 -100 107958
rect -158 105570 -146 107946
rect -112 105570 -100 107946
rect -158 105558 -100 105570
rect 100 107946 158 107958
rect 100 105570 112 107946
rect 146 105570 158 107946
rect 100 105558 158 105570
rect -158 105310 -100 105322
rect -158 102934 -146 105310
rect -112 102934 -100 105310
rect -158 102922 -100 102934
rect 100 105310 158 105322
rect 100 102934 112 105310
rect 146 102934 158 105310
rect 100 102922 158 102934
rect -158 102674 -100 102686
rect -158 100298 -146 102674
rect -112 100298 -100 102674
rect -158 100286 -100 100298
rect 100 102674 158 102686
rect 100 100298 112 102674
rect 146 100298 158 102674
rect 100 100286 158 100298
rect -158 100038 -100 100050
rect -158 97662 -146 100038
rect -112 97662 -100 100038
rect -158 97650 -100 97662
rect 100 100038 158 100050
rect 100 97662 112 100038
rect 146 97662 158 100038
rect 100 97650 158 97662
rect -158 97402 -100 97414
rect -158 95026 -146 97402
rect -112 95026 -100 97402
rect -158 95014 -100 95026
rect 100 97402 158 97414
rect 100 95026 112 97402
rect 146 95026 158 97402
rect 100 95014 158 95026
rect -158 94766 -100 94778
rect -158 92390 -146 94766
rect -112 92390 -100 94766
rect -158 92378 -100 92390
rect 100 94766 158 94778
rect 100 92390 112 94766
rect 146 92390 158 94766
rect 100 92378 158 92390
rect -158 92130 -100 92142
rect -158 89754 -146 92130
rect -112 89754 -100 92130
rect -158 89742 -100 89754
rect 100 92130 158 92142
rect 100 89754 112 92130
rect 146 89754 158 92130
rect 100 89742 158 89754
rect -158 89494 -100 89506
rect -158 87118 -146 89494
rect -112 87118 -100 89494
rect -158 87106 -100 87118
rect 100 89494 158 89506
rect 100 87118 112 89494
rect 146 87118 158 89494
rect 100 87106 158 87118
rect -158 86858 -100 86870
rect -158 84482 -146 86858
rect -112 84482 -100 86858
rect -158 84470 -100 84482
rect 100 86858 158 86870
rect 100 84482 112 86858
rect 146 84482 158 86858
rect 100 84470 158 84482
rect -158 84222 -100 84234
rect -158 81846 -146 84222
rect -112 81846 -100 84222
rect -158 81834 -100 81846
rect 100 84222 158 84234
rect 100 81846 112 84222
rect 146 81846 158 84222
rect 100 81834 158 81846
rect -158 81586 -100 81598
rect -158 79210 -146 81586
rect -112 79210 -100 81586
rect -158 79198 -100 79210
rect 100 81586 158 81598
rect 100 79210 112 81586
rect 146 79210 158 81586
rect 100 79198 158 79210
rect -158 78950 -100 78962
rect -158 76574 -146 78950
rect -112 76574 -100 78950
rect -158 76562 -100 76574
rect 100 78950 158 78962
rect 100 76574 112 78950
rect 146 76574 158 78950
rect 100 76562 158 76574
rect -158 76314 -100 76326
rect -158 73938 -146 76314
rect -112 73938 -100 76314
rect -158 73926 -100 73938
rect 100 76314 158 76326
rect 100 73938 112 76314
rect 146 73938 158 76314
rect 100 73926 158 73938
rect -158 73678 -100 73690
rect -158 71302 -146 73678
rect -112 71302 -100 73678
rect -158 71290 -100 71302
rect 100 73678 158 73690
rect 100 71302 112 73678
rect 146 71302 158 73678
rect 100 71290 158 71302
rect -158 71042 -100 71054
rect -158 68666 -146 71042
rect -112 68666 -100 71042
rect -158 68654 -100 68666
rect 100 71042 158 71054
rect 100 68666 112 71042
rect 146 68666 158 71042
rect 100 68654 158 68666
rect -158 68406 -100 68418
rect -158 66030 -146 68406
rect -112 66030 -100 68406
rect -158 66018 -100 66030
rect 100 68406 158 68418
rect 100 66030 112 68406
rect 146 66030 158 68406
rect 100 66018 158 66030
rect -158 65770 -100 65782
rect -158 63394 -146 65770
rect -112 63394 -100 65770
rect -158 63382 -100 63394
rect 100 65770 158 65782
rect 100 63394 112 65770
rect 146 63394 158 65770
rect 100 63382 158 63394
rect -158 63134 -100 63146
rect -158 60758 -146 63134
rect -112 60758 -100 63134
rect -158 60746 -100 60758
rect 100 63134 158 63146
rect 100 60758 112 63134
rect 146 60758 158 63134
rect 100 60746 158 60758
rect -158 60498 -100 60510
rect -158 58122 -146 60498
rect -112 58122 -100 60498
rect -158 58110 -100 58122
rect 100 60498 158 60510
rect 100 58122 112 60498
rect 146 58122 158 60498
rect 100 58110 158 58122
rect -158 57862 -100 57874
rect -158 55486 -146 57862
rect -112 55486 -100 57862
rect -158 55474 -100 55486
rect 100 57862 158 57874
rect 100 55486 112 57862
rect 146 55486 158 57862
rect 100 55474 158 55486
rect -158 55226 -100 55238
rect -158 52850 -146 55226
rect -112 52850 -100 55226
rect -158 52838 -100 52850
rect 100 55226 158 55238
rect 100 52850 112 55226
rect 146 52850 158 55226
rect 100 52838 158 52850
rect -158 52590 -100 52602
rect -158 50214 -146 52590
rect -112 50214 -100 52590
rect -158 50202 -100 50214
rect 100 52590 158 52602
rect 100 50214 112 52590
rect 146 50214 158 52590
rect 100 50202 158 50214
rect -158 49954 -100 49966
rect -158 47578 -146 49954
rect -112 47578 -100 49954
rect -158 47566 -100 47578
rect 100 49954 158 49966
rect 100 47578 112 49954
rect 146 47578 158 49954
rect 100 47566 158 47578
rect -158 47318 -100 47330
rect -158 44942 -146 47318
rect -112 44942 -100 47318
rect -158 44930 -100 44942
rect 100 47318 158 47330
rect 100 44942 112 47318
rect 146 44942 158 47318
rect 100 44930 158 44942
rect -158 44682 -100 44694
rect -158 42306 -146 44682
rect -112 42306 -100 44682
rect -158 42294 -100 42306
rect 100 44682 158 44694
rect 100 42306 112 44682
rect 146 42306 158 44682
rect 100 42294 158 42306
rect -158 42046 -100 42058
rect -158 39670 -146 42046
rect -112 39670 -100 42046
rect -158 39658 -100 39670
rect 100 42046 158 42058
rect 100 39670 112 42046
rect 146 39670 158 42046
rect 100 39658 158 39670
rect -158 39410 -100 39422
rect -158 37034 -146 39410
rect -112 37034 -100 39410
rect -158 37022 -100 37034
rect 100 39410 158 39422
rect 100 37034 112 39410
rect 146 37034 158 39410
rect 100 37022 158 37034
rect -158 36774 -100 36786
rect -158 34398 -146 36774
rect -112 34398 -100 36774
rect -158 34386 -100 34398
rect 100 36774 158 36786
rect 100 34398 112 36774
rect 146 34398 158 36774
rect 100 34386 158 34398
rect -158 34138 -100 34150
rect -158 31762 -146 34138
rect -112 31762 -100 34138
rect -158 31750 -100 31762
rect 100 34138 158 34150
rect 100 31762 112 34138
rect 146 31762 158 34138
rect 100 31750 158 31762
rect -158 31502 -100 31514
rect -158 29126 -146 31502
rect -112 29126 -100 31502
rect -158 29114 -100 29126
rect 100 31502 158 31514
rect 100 29126 112 31502
rect 146 29126 158 31502
rect 100 29114 158 29126
rect -158 28866 -100 28878
rect -158 26490 -146 28866
rect -112 26490 -100 28866
rect -158 26478 -100 26490
rect 100 28866 158 28878
rect 100 26490 112 28866
rect 146 26490 158 28866
rect 100 26478 158 26490
rect -158 26230 -100 26242
rect -158 23854 -146 26230
rect -112 23854 -100 26230
rect -158 23842 -100 23854
rect 100 26230 158 26242
rect 100 23854 112 26230
rect 146 23854 158 26230
rect 100 23842 158 23854
rect -158 23594 -100 23606
rect -158 21218 -146 23594
rect -112 21218 -100 23594
rect -158 21206 -100 21218
rect 100 23594 158 23606
rect 100 21218 112 23594
rect 146 21218 158 23594
rect 100 21206 158 21218
rect -158 20958 -100 20970
rect -158 18582 -146 20958
rect -112 18582 -100 20958
rect -158 18570 -100 18582
rect 100 20958 158 20970
rect 100 18582 112 20958
rect 146 18582 158 20958
rect 100 18570 158 18582
rect -158 18322 -100 18334
rect -158 15946 -146 18322
rect -112 15946 -100 18322
rect -158 15934 -100 15946
rect 100 18322 158 18334
rect 100 15946 112 18322
rect 146 15946 158 18322
rect 100 15934 158 15946
rect -158 15686 -100 15698
rect -158 13310 -146 15686
rect -112 13310 -100 15686
rect -158 13298 -100 13310
rect 100 15686 158 15698
rect 100 13310 112 15686
rect 146 13310 158 15686
rect 100 13298 158 13310
rect -158 13050 -100 13062
rect -158 10674 -146 13050
rect -112 10674 -100 13050
rect -158 10662 -100 10674
rect 100 13050 158 13062
rect 100 10674 112 13050
rect 146 10674 158 13050
rect 100 10662 158 10674
rect -158 10414 -100 10426
rect -158 8038 -146 10414
rect -112 8038 -100 10414
rect -158 8026 -100 8038
rect 100 10414 158 10426
rect 100 8038 112 10414
rect 146 8038 158 10414
rect 100 8026 158 8038
rect -158 7778 -100 7790
rect -158 5402 -146 7778
rect -112 5402 -100 7778
rect -158 5390 -100 5402
rect 100 7778 158 7790
rect 100 5402 112 7778
rect 146 5402 158 7778
rect 100 5390 158 5402
rect -158 5142 -100 5154
rect -158 2766 -146 5142
rect -112 2766 -100 5142
rect -158 2754 -100 2766
rect 100 5142 158 5154
rect 100 2766 112 5142
rect 146 2766 158 5142
rect 100 2754 158 2766
rect -158 2506 -100 2518
rect -158 130 -146 2506
rect -112 130 -100 2506
rect -158 118 -100 130
rect 100 2506 158 2518
rect 100 130 112 2506
rect 146 130 158 2506
rect 100 118 158 130
rect -158 -130 -100 -118
rect -158 -2506 -146 -130
rect -112 -2506 -100 -130
rect -158 -2518 -100 -2506
rect 100 -130 158 -118
rect 100 -2506 112 -130
rect 146 -2506 158 -130
rect 100 -2518 158 -2506
rect -158 -2766 -100 -2754
rect -158 -5142 -146 -2766
rect -112 -5142 -100 -2766
rect -158 -5154 -100 -5142
rect 100 -2766 158 -2754
rect 100 -5142 112 -2766
rect 146 -5142 158 -2766
rect 100 -5154 158 -5142
rect -158 -5402 -100 -5390
rect -158 -7778 -146 -5402
rect -112 -7778 -100 -5402
rect -158 -7790 -100 -7778
rect 100 -5402 158 -5390
rect 100 -7778 112 -5402
rect 146 -7778 158 -5402
rect 100 -7790 158 -7778
rect -158 -8038 -100 -8026
rect -158 -10414 -146 -8038
rect -112 -10414 -100 -8038
rect -158 -10426 -100 -10414
rect 100 -8038 158 -8026
rect 100 -10414 112 -8038
rect 146 -10414 158 -8038
rect 100 -10426 158 -10414
rect -158 -10674 -100 -10662
rect -158 -13050 -146 -10674
rect -112 -13050 -100 -10674
rect -158 -13062 -100 -13050
rect 100 -10674 158 -10662
rect 100 -13050 112 -10674
rect 146 -13050 158 -10674
rect 100 -13062 158 -13050
rect -158 -13310 -100 -13298
rect -158 -15686 -146 -13310
rect -112 -15686 -100 -13310
rect -158 -15698 -100 -15686
rect 100 -13310 158 -13298
rect 100 -15686 112 -13310
rect 146 -15686 158 -13310
rect 100 -15698 158 -15686
rect -158 -15946 -100 -15934
rect -158 -18322 -146 -15946
rect -112 -18322 -100 -15946
rect -158 -18334 -100 -18322
rect 100 -15946 158 -15934
rect 100 -18322 112 -15946
rect 146 -18322 158 -15946
rect 100 -18334 158 -18322
rect -158 -18582 -100 -18570
rect -158 -20958 -146 -18582
rect -112 -20958 -100 -18582
rect -158 -20970 -100 -20958
rect 100 -18582 158 -18570
rect 100 -20958 112 -18582
rect 146 -20958 158 -18582
rect 100 -20970 158 -20958
rect -158 -21218 -100 -21206
rect -158 -23594 -146 -21218
rect -112 -23594 -100 -21218
rect -158 -23606 -100 -23594
rect 100 -21218 158 -21206
rect 100 -23594 112 -21218
rect 146 -23594 158 -21218
rect 100 -23606 158 -23594
rect -158 -23854 -100 -23842
rect -158 -26230 -146 -23854
rect -112 -26230 -100 -23854
rect -158 -26242 -100 -26230
rect 100 -23854 158 -23842
rect 100 -26230 112 -23854
rect 146 -26230 158 -23854
rect 100 -26242 158 -26230
rect -158 -26490 -100 -26478
rect -158 -28866 -146 -26490
rect -112 -28866 -100 -26490
rect -158 -28878 -100 -28866
rect 100 -26490 158 -26478
rect 100 -28866 112 -26490
rect 146 -28866 158 -26490
rect 100 -28878 158 -28866
rect -158 -29126 -100 -29114
rect -158 -31502 -146 -29126
rect -112 -31502 -100 -29126
rect -158 -31514 -100 -31502
rect 100 -29126 158 -29114
rect 100 -31502 112 -29126
rect 146 -31502 158 -29126
rect 100 -31514 158 -31502
rect -158 -31762 -100 -31750
rect -158 -34138 -146 -31762
rect -112 -34138 -100 -31762
rect -158 -34150 -100 -34138
rect 100 -31762 158 -31750
rect 100 -34138 112 -31762
rect 146 -34138 158 -31762
rect 100 -34150 158 -34138
rect -158 -34398 -100 -34386
rect -158 -36774 -146 -34398
rect -112 -36774 -100 -34398
rect -158 -36786 -100 -36774
rect 100 -34398 158 -34386
rect 100 -36774 112 -34398
rect 146 -36774 158 -34398
rect 100 -36786 158 -36774
rect -158 -37034 -100 -37022
rect -158 -39410 -146 -37034
rect -112 -39410 -100 -37034
rect -158 -39422 -100 -39410
rect 100 -37034 158 -37022
rect 100 -39410 112 -37034
rect 146 -39410 158 -37034
rect 100 -39422 158 -39410
rect -158 -39670 -100 -39658
rect -158 -42046 -146 -39670
rect -112 -42046 -100 -39670
rect -158 -42058 -100 -42046
rect 100 -39670 158 -39658
rect 100 -42046 112 -39670
rect 146 -42046 158 -39670
rect 100 -42058 158 -42046
rect -158 -42306 -100 -42294
rect -158 -44682 -146 -42306
rect -112 -44682 -100 -42306
rect -158 -44694 -100 -44682
rect 100 -42306 158 -42294
rect 100 -44682 112 -42306
rect 146 -44682 158 -42306
rect 100 -44694 158 -44682
rect -158 -44942 -100 -44930
rect -158 -47318 -146 -44942
rect -112 -47318 -100 -44942
rect -158 -47330 -100 -47318
rect 100 -44942 158 -44930
rect 100 -47318 112 -44942
rect 146 -47318 158 -44942
rect 100 -47330 158 -47318
rect -158 -47578 -100 -47566
rect -158 -49954 -146 -47578
rect -112 -49954 -100 -47578
rect -158 -49966 -100 -49954
rect 100 -47578 158 -47566
rect 100 -49954 112 -47578
rect 146 -49954 158 -47578
rect 100 -49966 158 -49954
rect -158 -50214 -100 -50202
rect -158 -52590 -146 -50214
rect -112 -52590 -100 -50214
rect -158 -52602 -100 -52590
rect 100 -50214 158 -50202
rect 100 -52590 112 -50214
rect 146 -52590 158 -50214
rect 100 -52602 158 -52590
rect -158 -52850 -100 -52838
rect -158 -55226 -146 -52850
rect -112 -55226 -100 -52850
rect -158 -55238 -100 -55226
rect 100 -52850 158 -52838
rect 100 -55226 112 -52850
rect 146 -55226 158 -52850
rect 100 -55238 158 -55226
rect -158 -55486 -100 -55474
rect -158 -57862 -146 -55486
rect -112 -57862 -100 -55486
rect -158 -57874 -100 -57862
rect 100 -55486 158 -55474
rect 100 -57862 112 -55486
rect 146 -57862 158 -55486
rect 100 -57874 158 -57862
rect -158 -58122 -100 -58110
rect -158 -60498 -146 -58122
rect -112 -60498 -100 -58122
rect -158 -60510 -100 -60498
rect 100 -58122 158 -58110
rect 100 -60498 112 -58122
rect 146 -60498 158 -58122
rect 100 -60510 158 -60498
rect -158 -60758 -100 -60746
rect -158 -63134 -146 -60758
rect -112 -63134 -100 -60758
rect -158 -63146 -100 -63134
rect 100 -60758 158 -60746
rect 100 -63134 112 -60758
rect 146 -63134 158 -60758
rect 100 -63146 158 -63134
rect -158 -63394 -100 -63382
rect -158 -65770 -146 -63394
rect -112 -65770 -100 -63394
rect -158 -65782 -100 -65770
rect 100 -63394 158 -63382
rect 100 -65770 112 -63394
rect 146 -65770 158 -63394
rect 100 -65782 158 -65770
rect -158 -66030 -100 -66018
rect -158 -68406 -146 -66030
rect -112 -68406 -100 -66030
rect -158 -68418 -100 -68406
rect 100 -66030 158 -66018
rect 100 -68406 112 -66030
rect 146 -68406 158 -66030
rect 100 -68418 158 -68406
rect -158 -68666 -100 -68654
rect -158 -71042 -146 -68666
rect -112 -71042 -100 -68666
rect -158 -71054 -100 -71042
rect 100 -68666 158 -68654
rect 100 -71042 112 -68666
rect 146 -71042 158 -68666
rect 100 -71054 158 -71042
rect -158 -71302 -100 -71290
rect -158 -73678 -146 -71302
rect -112 -73678 -100 -71302
rect -158 -73690 -100 -73678
rect 100 -71302 158 -71290
rect 100 -73678 112 -71302
rect 146 -73678 158 -71302
rect 100 -73690 158 -73678
rect -158 -73938 -100 -73926
rect -158 -76314 -146 -73938
rect -112 -76314 -100 -73938
rect -158 -76326 -100 -76314
rect 100 -73938 158 -73926
rect 100 -76314 112 -73938
rect 146 -76314 158 -73938
rect 100 -76326 158 -76314
rect -158 -76574 -100 -76562
rect -158 -78950 -146 -76574
rect -112 -78950 -100 -76574
rect -158 -78962 -100 -78950
rect 100 -76574 158 -76562
rect 100 -78950 112 -76574
rect 146 -78950 158 -76574
rect 100 -78962 158 -78950
rect -158 -79210 -100 -79198
rect -158 -81586 -146 -79210
rect -112 -81586 -100 -79210
rect -158 -81598 -100 -81586
rect 100 -79210 158 -79198
rect 100 -81586 112 -79210
rect 146 -81586 158 -79210
rect 100 -81598 158 -81586
rect -158 -81846 -100 -81834
rect -158 -84222 -146 -81846
rect -112 -84222 -100 -81846
rect -158 -84234 -100 -84222
rect 100 -81846 158 -81834
rect 100 -84222 112 -81846
rect 146 -84222 158 -81846
rect 100 -84234 158 -84222
rect -158 -84482 -100 -84470
rect -158 -86858 -146 -84482
rect -112 -86858 -100 -84482
rect -158 -86870 -100 -86858
rect 100 -84482 158 -84470
rect 100 -86858 112 -84482
rect 146 -86858 158 -84482
rect 100 -86870 158 -86858
rect -158 -87118 -100 -87106
rect -158 -89494 -146 -87118
rect -112 -89494 -100 -87118
rect -158 -89506 -100 -89494
rect 100 -87118 158 -87106
rect 100 -89494 112 -87118
rect 146 -89494 158 -87118
rect 100 -89506 158 -89494
rect -158 -89754 -100 -89742
rect -158 -92130 -146 -89754
rect -112 -92130 -100 -89754
rect -158 -92142 -100 -92130
rect 100 -89754 158 -89742
rect 100 -92130 112 -89754
rect 146 -92130 158 -89754
rect 100 -92142 158 -92130
rect -158 -92390 -100 -92378
rect -158 -94766 -146 -92390
rect -112 -94766 -100 -92390
rect -158 -94778 -100 -94766
rect 100 -92390 158 -92378
rect 100 -94766 112 -92390
rect 146 -94766 158 -92390
rect 100 -94778 158 -94766
rect -158 -95026 -100 -95014
rect -158 -97402 -146 -95026
rect -112 -97402 -100 -95026
rect -158 -97414 -100 -97402
rect 100 -95026 158 -95014
rect 100 -97402 112 -95026
rect 146 -97402 158 -95026
rect 100 -97414 158 -97402
rect -158 -97662 -100 -97650
rect -158 -100038 -146 -97662
rect -112 -100038 -100 -97662
rect -158 -100050 -100 -100038
rect 100 -97662 158 -97650
rect 100 -100038 112 -97662
rect 146 -100038 158 -97662
rect 100 -100050 158 -100038
rect -158 -100298 -100 -100286
rect -158 -102674 -146 -100298
rect -112 -102674 -100 -100298
rect -158 -102686 -100 -102674
rect 100 -100298 158 -100286
rect 100 -102674 112 -100298
rect 146 -102674 158 -100298
rect 100 -102686 158 -102674
rect -158 -102934 -100 -102922
rect -158 -105310 -146 -102934
rect -112 -105310 -100 -102934
rect -158 -105322 -100 -105310
rect 100 -102934 158 -102922
rect 100 -105310 112 -102934
rect 146 -105310 158 -102934
rect 100 -105322 158 -105310
rect -158 -105570 -100 -105558
rect -158 -107946 -146 -105570
rect -112 -107946 -100 -105570
rect -158 -107958 -100 -107946
rect 100 -105570 158 -105558
rect 100 -107946 112 -105570
rect 146 -107946 158 -105570
rect 100 -107958 158 -107946
rect -158 -108206 -100 -108194
rect -158 -110582 -146 -108206
rect -112 -110582 -100 -108206
rect -158 -110594 -100 -110582
rect 100 -108206 158 -108194
rect 100 -110582 112 -108206
rect 146 -110582 158 -108206
rect 100 -110594 158 -110582
rect -158 -110842 -100 -110830
rect -158 -113218 -146 -110842
rect -112 -113218 -100 -110842
rect -158 -113230 -100 -113218
rect 100 -110842 158 -110830
rect 100 -113218 112 -110842
rect 146 -113218 158 -110842
rect 100 -113230 158 -113218
rect -158 -113478 -100 -113466
rect -158 -115854 -146 -113478
rect -112 -115854 -100 -113478
rect -158 -115866 -100 -115854
rect 100 -113478 158 -113466
rect 100 -115854 112 -113478
rect 146 -115854 158 -113478
rect 100 -115866 158 -115854
rect -158 -116114 -100 -116102
rect -158 -118490 -146 -116114
rect -112 -118490 -100 -116114
rect -158 -118502 -100 -118490
rect 100 -116114 158 -116102
rect 100 -118490 112 -116114
rect 146 -118490 158 -116114
rect 100 -118502 158 -118490
rect -158 -118750 -100 -118738
rect -158 -121126 -146 -118750
rect -112 -121126 -100 -118750
rect -158 -121138 -100 -121126
rect 100 -118750 158 -118738
rect 100 -121126 112 -118750
rect 146 -121126 158 -118750
rect 100 -121138 158 -121126
rect -158 -121386 -100 -121374
rect -158 -123762 -146 -121386
rect -112 -123762 -100 -121386
rect -158 -123774 -100 -123762
rect 100 -121386 158 -121374
rect 100 -123762 112 -121386
rect 146 -123762 158 -121386
rect 100 -123774 158 -123762
rect -158 -124022 -100 -124010
rect -158 -126398 -146 -124022
rect -112 -126398 -100 -124022
rect -158 -126410 -100 -126398
rect 100 -124022 158 -124010
rect 100 -126398 112 -124022
rect 146 -126398 158 -124022
rect 100 -126410 158 -126398
rect -158 -126658 -100 -126646
rect -158 -129034 -146 -126658
rect -112 -129034 -100 -126658
rect -158 -129046 -100 -129034
rect 100 -126658 158 -126646
rect 100 -129034 112 -126658
rect 146 -129034 158 -126658
rect 100 -129046 158 -129034
rect -158 -129294 -100 -129282
rect -158 -131670 -146 -129294
rect -112 -131670 -100 -129294
rect -158 -131682 -100 -131670
rect 100 -129294 158 -129282
rect 100 -131670 112 -129294
rect 146 -131670 158 -129294
rect 100 -131682 158 -131670
rect -158 -131930 -100 -131918
rect -158 -134306 -146 -131930
rect -112 -134306 -100 -131930
rect -158 -134318 -100 -134306
rect 100 -131930 158 -131918
rect 100 -134306 112 -131930
rect 146 -134306 158 -131930
rect 100 -134318 158 -134306
rect -158 -134566 -100 -134554
rect -158 -136942 -146 -134566
rect -112 -136942 -100 -134566
rect -158 -136954 -100 -136942
rect 100 -134566 158 -134554
rect 100 -136942 112 -134566
rect 146 -136942 158 -134566
rect 100 -136954 158 -136942
rect -158 -137202 -100 -137190
rect -158 -139578 -146 -137202
rect -112 -139578 -100 -137202
rect -158 -139590 -100 -139578
rect 100 -137202 158 -137190
rect 100 -139578 112 -137202
rect 146 -139578 158 -137202
rect 100 -139590 158 -139578
rect -158 -139838 -100 -139826
rect -158 -142214 -146 -139838
rect -112 -142214 -100 -139838
rect -158 -142226 -100 -142214
rect 100 -139838 158 -139826
rect 100 -142214 112 -139838
rect 146 -142214 158 -139838
rect 100 -142226 158 -142214
rect -158 -142474 -100 -142462
rect -158 -144850 -146 -142474
rect -112 -144850 -100 -142474
rect -158 -144862 -100 -144850
rect 100 -142474 158 -142462
rect 100 -144850 112 -142474
rect 146 -144850 158 -142474
rect 100 -144862 158 -144850
rect -158 -145110 -100 -145098
rect -158 -147486 -146 -145110
rect -112 -147486 -100 -145110
rect -158 -147498 -100 -147486
rect 100 -145110 158 -145098
rect 100 -147486 112 -145110
rect 146 -147486 158 -145110
rect 100 -147498 158 -147486
rect -158 -147746 -100 -147734
rect -158 -150122 -146 -147746
rect -112 -150122 -100 -147746
rect -158 -150134 -100 -150122
rect 100 -147746 158 -147734
rect 100 -150122 112 -147746
rect 146 -150122 158 -147746
rect 100 -150134 158 -150122
rect -158 -150382 -100 -150370
rect -158 -152758 -146 -150382
rect -112 -152758 -100 -150382
rect -158 -152770 -100 -152758
rect 100 -150382 158 -150370
rect 100 -152758 112 -150382
rect 146 -152758 158 -150382
rect 100 -152770 158 -152758
rect -158 -153018 -100 -153006
rect -158 -155394 -146 -153018
rect -112 -155394 -100 -153018
rect -158 -155406 -100 -155394
rect 100 -153018 158 -153006
rect 100 -155394 112 -153018
rect 146 -155394 158 -153018
rect 100 -155406 158 -155394
rect -158 -155654 -100 -155642
rect -158 -158030 -146 -155654
rect -112 -158030 -100 -155654
rect -158 -158042 -100 -158030
rect 100 -155654 158 -155642
rect 100 -158030 112 -155654
rect 146 -158030 158 -155654
rect 100 -158042 158 -158030
rect -158 -158290 -100 -158278
rect -158 -160666 -146 -158290
rect -112 -160666 -100 -158290
rect -158 -160678 -100 -160666
rect 100 -158290 158 -158278
rect 100 -160666 112 -158290
rect 146 -160666 158 -158290
rect 100 -160678 158 -160666
rect -158 -160926 -100 -160914
rect -158 -163302 -146 -160926
rect -112 -163302 -100 -160926
rect -158 -163314 -100 -163302
rect 100 -160926 158 -160914
rect 100 -163302 112 -160926
rect 146 -163302 158 -160926
rect 100 -163314 158 -163302
rect -158 -163562 -100 -163550
rect -158 -165938 -146 -163562
rect -112 -165938 -100 -163562
rect -158 -165950 -100 -165938
rect 100 -163562 158 -163550
rect 100 -165938 112 -163562
rect 146 -165938 158 -163562
rect 100 -165950 158 -165938
rect -158 -166198 -100 -166186
rect -158 -168574 -146 -166198
rect -112 -168574 -100 -166198
rect -158 -168586 -100 -168574
rect 100 -166198 158 -166186
rect 100 -168574 112 -166198
rect 146 -168574 158 -166198
rect 100 -168586 158 -168574
rect -158 -168834 -100 -168822
rect -158 -171210 -146 -168834
rect -112 -171210 -100 -168834
rect -158 -171222 -100 -171210
rect 100 -168834 158 -168822
rect 100 -171210 112 -168834
rect 146 -171210 158 -168834
rect 100 -171222 158 -171210
rect -158 -171470 -100 -171458
rect -158 -173846 -146 -171470
rect -112 -173846 -100 -171470
rect -158 -173858 -100 -173846
rect 100 -171470 158 -171458
rect 100 -173846 112 -171470
rect 146 -173846 158 -171470
rect 100 -173858 158 -173846
rect -158 -174106 -100 -174094
rect -158 -176482 -146 -174106
rect -112 -176482 -100 -174106
rect -158 -176494 -100 -176482
rect 100 -174106 158 -174094
rect 100 -176482 112 -174106
rect 146 -176482 158 -174106
rect 100 -176494 158 -176482
rect -158 -176742 -100 -176730
rect -158 -179118 -146 -176742
rect -112 -179118 -100 -176742
rect -158 -179130 -100 -179118
rect 100 -176742 158 -176730
rect 100 -179118 112 -176742
rect 146 -179118 158 -176742
rect 100 -179130 158 -179118
rect -158 -179378 -100 -179366
rect -158 -181754 -146 -179378
rect -112 -181754 -100 -179378
rect -158 -181766 -100 -181754
rect 100 -179378 158 -179366
rect 100 -181754 112 -179378
rect 146 -181754 158 -179378
rect 100 -181766 158 -181754
rect -158 -182014 -100 -182002
rect -158 -184390 -146 -182014
rect -112 -184390 -100 -182014
rect -158 -184402 -100 -184390
rect 100 -182014 158 -182002
rect 100 -184390 112 -182014
rect 146 -184390 158 -182014
rect 100 -184402 158 -184390
rect -158 -184650 -100 -184638
rect -158 -187026 -146 -184650
rect -112 -187026 -100 -184650
rect -158 -187038 -100 -187026
rect 100 -184650 158 -184638
rect 100 -187026 112 -184650
rect 146 -187026 158 -184650
rect 100 -187038 158 -187026
rect -158 -187286 -100 -187274
rect -158 -189662 -146 -187286
rect -112 -189662 -100 -187286
rect -158 -189674 -100 -189662
rect 100 -187286 158 -187274
rect 100 -189662 112 -187286
rect 146 -189662 158 -187286
rect 100 -189674 158 -189662
rect -158 -189922 -100 -189910
rect -158 -192298 -146 -189922
rect -112 -192298 -100 -189922
rect -158 -192310 -100 -192298
rect 100 -189922 158 -189910
rect 100 -192298 112 -189922
rect 146 -192298 158 -189922
rect 100 -192310 158 -192298
rect -158 -192558 -100 -192546
rect -158 -194934 -146 -192558
rect -112 -194934 -100 -192558
rect -158 -194946 -100 -194934
rect 100 -192558 158 -192546
rect 100 -194934 112 -192558
rect 146 -194934 158 -192558
rect 100 -194946 158 -194934
rect -158 -195194 -100 -195182
rect -158 -197570 -146 -195194
rect -112 -197570 -100 -195194
rect -158 -197582 -100 -197570
rect 100 -195194 158 -195182
rect 100 -197570 112 -195194
rect 146 -197570 158 -195194
rect 100 -197582 158 -197570
rect -158 -197830 -100 -197818
rect -158 -200206 -146 -197830
rect -112 -200206 -100 -197830
rect -158 -200218 -100 -200206
rect 100 -197830 158 -197818
rect 100 -200206 112 -197830
rect 146 -200206 158 -197830
rect 100 -200218 158 -200206
rect -158 -200466 -100 -200454
rect -158 -202842 -146 -200466
rect -112 -202842 -100 -200466
rect -158 -202854 -100 -202842
rect 100 -200466 158 -200454
rect 100 -202842 112 -200466
rect 146 -202842 158 -200466
rect 100 -202854 158 -202842
rect -158 -203102 -100 -203090
rect -158 -205478 -146 -203102
rect -112 -205478 -100 -203102
rect -158 -205490 -100 -205478
rect 100 -203102 158 -203090
rect 100 -205478 112 -203102
rect 146 -205478 158 -203102
rect 100 -205490 158 -205478
rect -158 -205738 -100 -205726
rect -158 -208114 -146 -205738
rect -112 -208114 -100 -205738
rect -158 -208126 -100 -208114
rect 100 -205738 158 -205726
rect 100 -208114 112 -205738
rect 146 -208114 158 -205738
rect 100 -208126 158 -208114
rect -158 -208374 -100 -208362
rect -158 -210750 -146 -208374
rect -112 -210750 -100 -208374
rect -158 -210762 -100 -210750
rect 100 -208374 158 -208362
rect 100 -210750 112 -208374
rect 146 -210750 158 -208374
rect 100 -210762 158 -210750
rect -158 -211010 -100 -210998
rect -158 -213386 -146 -211010
rect -112 -213386 -100 -211010
rect -158 -213398 -100 -213386
rect 100 -211010 158 -210998
rect 100 -213386 112 -211010
rect 146 -213386 158 -211010
rect 100 -213398 158 -213386
rect -158 -213646 -100 -213634
rect -158 -216022 -146 -213646
rect -112 -216022 -100 -213646
rect -158 -216034 -100 -216022
rect 100 -213646 158 -213634
rect 100 -216022 112 -213646
rect 146 -216022 158 -213646
rect 100 -216034 158 -216022
rect -158 -216282 -100 -216270
rect -158 -218658 -146 -216282
rect -112 -218658 -100 -216282
rect -158 -218670 -100 -218658
rect 100 -216282 158 -216270
rect 100 -218658 112 -216282
rect 146 -218658 158 -216282
rect 100 -218670 158 -218658
rect -158 -218918 -100 -218906
rect -158 -221294 -146 -218918
rect -112 -221294 -100 -218918
rect -158 -221306 -100 -221294
rect 100 -218918 158 -218906
rect 100 -221294 112 -218918
rect 146 -221294 158 -218918
rect 100 -221306 158 -221294
rect -158 -221554 -100 -221542
rect -158 -223930 -146 -221554
rect -112 -223930 -100 -221554
rect -158 -223942 -100 -223930
rect 100 -221554 158 -221542
rect 100 -223930 112 -221554
rect 146 -223930 158 -221554
rect 100 -223942 158 -223930
rect -158 -224190 -100 -224178
rect -158 -226566 -146 -224190
rect -112 -226566 -100 -224190
rect -158 -226578 -100 -226566
rect 100 -224190 158 -224178
rect 100 -226566 112 -224190
rect 146 -226566 158 -224190
rect 100 -226578 158 -226566
rect -158 -226826 -100 -226814
rect -158 -229202 -146 -226826
rect -112 -229202 -100 -226826
rect -158 -229214 -100 -229202
rect 100 -226826 158 -226814
rect 100 -229202 112 -226826
rect 146 -229202 158 -226826
rect 100 -229214 158 -229202
rect -158 -229462 -100 -229450
rect -158 -231838 -146 -229462
rect -112 -231838 -100 -229462
rect -158 -231850 -100 -231838
rect 100 -229462 158 -229450
rect 100 -231838 112 -229462
rect 146 -231838 158 -229462
rect 100 -231850 158 -231838
rect -158 -232098 -100 -232086
rect -158 -234474 -146 -232098
rect -112 -234474 -100 -232098
rect -158 -234486 -100 -234474
rect 100 -232098 158 -232086
rect 100 -234474 112 -232098
rect 146 -234474 158 -232098
rect 100 -234486 158 -234474
rect -158 -234734 -100 -234722
rect -158 -237110 -146 -234734
rect -112 -237110 -100 -234734
rect -158 -237122 -100 -237110
rect 100 -234734 158 -234722
rect 100 -237110 112 -234734
rect 146 -237110 158 -234734
rect 100 -237122 158 -237110
rect -158 -237370 -100 -237358
rect -158 -239746 -146 -237370
rect -112 -239746 -100 -237370
rect -158 -239758 -100 -239746
rect 100 -237370 158 -237358
rect 100 -239746 112 -237370
rect 146 -239746 158 -237370
rect 100 -239758 158 -239746
rect -158 -240006 -100 -239994
rect -158 -242382 -146 -240006
rect -112 -242382 -100 -240006
rect -158 -242394 -100 -242382
rect 100 -240006 158 -239994
rect 100 -242382 112 -240006
rect 146 -242382 158 -240006
rect 100 -242394 158 -242382
rect -158 -242642 -100 -242630
rect -158 -245018 -146 -242642
rect -112 -245018 -100 -242642
rect -158 -245030 -100 -245018
rect 100 -242642 158 -242630
rect 100 -245018 112 -242642
rect 146 -245018 158 -242642
rect 100 -245030 158 -245018
rect -158 -245278 -100 -245266
rect -158 -247654 -146 -245278
rect -112 -247654 -100 -245278
rect -158 -247666 -100 -247654
rect 100 -245278 158 -245266
rect 100 -247654 112 -245278
rect 146 -247654 158 -245278
rect 100 -247666 158 -247654
rect -158 -247914 -100 -247902
rect -158 -250290 -146 -247914
rect -112 -250290 -100 -247914
rect -158 -250302 -100 -250290
rect 100 -247914 158 -247902
rect 100 -250290 112 -247914
rect 146 -250290 158 -247914
rect 100 -250302 158 -250290
rect -158 -250550 -100 -250538
rect -158 -252926 -146 -250550
rect -112 -252926 -100 -250550
rect -158 -252938 -100 -252926
rect 100 -250550 158 -250538
rect 100 -252926 112 -250550
rect 146 -252926 158 -250550
rect 100 -252938 158 -252926
rect -158 -253186 -100 -253174
rect -158 -255562 -146 -253186
rect -112 -255562 -100 -253186
rect -158 -255574 -100 -255562
rect 100 -253186 158 -253174
rect 100 -255562 112 -253186
rect 146 -255562 158 -253186
rect 100 -255574 158 -255562
rect -158 -255822 -100 -255810
rect -158 -258198 -146 -255822
rect -112 -258198 -100 -255822
rect -158 -258210 -100 -258198
rect 100 -255822 158 -255810
rect 100 -258198 112 -255822
rect 146 -258198 158 -255822
rect 100 -258210 158 -258198
rect -158 -258458 -100 -258446
rect -158 -260834 -146 -258458
rect -112 -260834 -100 -258458
rect -158 -260846 -100 -260834
rect 100 -258458 158 -258446
rect 100 -260834 112 -258458
rect 146 -260834 158 -258458
rect 100 -260846 158 -260834
rect -158 -261094 -100 -261082
rect -158 -263470 -146 -261094
rect -112 -263470 -100 -261094
rect -158 -263482 -100 -263470
rect 100 -261094 158 -261082
rect 100 -263470 112 -261094
rect 146 -263470 158 -261094
rect 100 -263482 158 -263470
rect -158 -263730 -100 -263718
rect -158 -266106 -146 -263730
rect -112 -266106 -100 -263730
rect -158 -266118 -100 -266106
rect 100 -263730 158 -263718
rect 100 -266106 112 -263730
rect 146 -266106 158 -263730
rect 100 -266118 158 -266106
rect -158 -266366 -100 -266354
rect -158 -268742 -146 -266366
rect -112 -268742 -100 -266366
rect -158 -268754 -100 -268742
rect 100 -266366 158 -266354
rect 100 -268742 112 -266366
rect 146 -268742 158 -266366
rect 100 -268754 158 -268742
rect -158 -269002 -100 -268990
rect -158 -271378 -146 -269002
rect -112 -271378 -100 -269002
rect -158 -271390 -100 -271378
rect 100 -269002 158 -268990
rect 100 -271378 112 -269002
rect 146 -271378 158 -269002
rect 100 -271390 158 -271378
rect -158 -271638 -100 -271626
rect -158 -274014 -146 -271638
rect -112 -274014 -100 -271638
rect -158 -274026 -100 -274014
rect 100 -271638 158 -271626
rect 100 -274014 112 -271638
rect 146 -274014 158 -271638
rect 100 -274026 158 -274014
rect -158 -274274 -100 -274262
rect -158 -276650 -146 -274274
rect -112 -276650 -100 -274274
rect -158 -276662 -100 -276650
rect 100 -274274 158 -274262
rect 100 -276650 112 -274274
rect 146 -276650 158 -274274
rect 100 -276662 158 -276650
rect -158 -276910 -100 -276898
rect -158 -279286 -146 -276910
rect -112 -279286 -100 -276910
rect -158 -279298 -100 -279286
rect 100 -276910 158 -276898
rect 100 -279286 112 -276910
rect 146 -279286 158 -276910
rect 100 -279298 158 -279286
rect -158 -279546 -100 -279534
rect -158 -281922 -146 -279546
rect -112 -281922 -100 -279546
rect -158 -281934 -100 -281922
rect 100 -279546 158 -279534
rect 100 -281922 112 -279546
rect 146 -281922 158 -279546
rect 100 -281934 158 -281922
rect -158 -282182 -100 -282170
rect -158 -284558 -146 -282182
rect -112 -284558 -100 -282182
rect -158 -284570 -100 -284558
rect 100 -282182 158 -282170
rect 100 -284558 112 -282182
rect 146 -284558 158 -282182
rect 100 -284570 158 -284558
rect -158 -284818 -100 -284806
rect -158 -287194 -146 -284818
rect -112 -287194 -100 -284818
rect -158 -287206 -100 -287194
rect 100 -284818 158 -284806
rect 100 -287194 112 -284818
rect 146 -287194 158 -284818
rect 100 -287206 158 -287194
rect -158 -287454 -100 -287442
rect -158 -289830 -146 -287454
rect -112 -289830 -100 -287454
rect -158 -289842 -100 -289830
rect 100 -287454 158 -287442
rect 100 -289830 112 -287454
rect 146 -289830 158 -287454
rect 100 -289842 158 -289830
rect -158 -290090 -100 -290078
rect -158 -292466 -146 -290090
rect -112 -292466 -100 -290090
rect -158 -292478 -100 -292466
rect 100 -290090 158 -290078
rect 100 -292466 112 -290090
rect 146 -292466 158 -290090
rect 100 -292478 158 -292466
rect -158 -292726 -100 -292714
rect -158 -295102 -146 -292726
rect -112 -295102 -100 -292726
rect -158 -295114 -100 -295102
rect 100 -292726 158 -292714
rect 100 -295102 112 -292726
rect 146 -295102 158 -292726
rect 100 -295114 158 -295102
rect -158 -295362 -100 -295350
rect -158 -297738 -146 -295362
rect -112 -297738 -100 -295362
rect -158 -297750 -100 -297738
rect 100 -295362 158 -295350
rect 100 -297738 112 -295362
rect 146 -297738 158 -295362
rect 100 -297750 158 -297738
rect -158 -297998 -100 -297986
rect -158 -300374 -146 -297998
rect -112 -300374 -100 -297998
rect -158 -300386 -100 -300374
rect 100 -297998 158 -297986
rect 100 -300374 112 -297998
rect 146 -300374 158 -297998
rect 100 -300386 158 -300374
rect -158 -300634 -100 -300622
rect -158 -303010 -146 -300634
rect -112 -303010 -100 -300634
rect -158 -303022 -100 -303010
rect 100 -300634 158 -300622
rect 100 -303010 112 -300634
rect 146 -303010 158 -300634
rect 100 -303022 158 -303010
rect -158 -303270 -100 -303258
rect -158 -305646 -146 -303270
rect -112 -305646 -100 -303270
rect -158 -305658 -100 -305646
rect 100 -303270 158 -303258
rect 100 -305646 112 -303270
rect 146 -305646 158 -303270
rect 100 -305658 158 -305646
rect -158 -305906 -100 -305894
rect -158 -308282 -146 -305906
rect -112 -308282 -100 -305906
rect -158 -308294 -100 -308282
rect 100 -305906 158 -305894
rect 100 -308282 112 -305906
rect 146 -308282 158 -305906
rect 100 -308294 158 -308282
rect -158 -308542 -100 -308530
rect -158 -310918 -146 -308542
rect -112 -310918 -100 -308542
rect -158 -310930 -100 -310918
rect 100 -308542 158 -308530
rect 100 -310918 112 -308542
rect 146 -310918 158 -308542
rect 100 -310930 158 -310918
rect -158 -311178 -100 -311166
rect -158 -313554 -146 -311178
rect -112 -313554 -100 -311178
rect -158 -313566 -100 -313554
rect 100 -311178 158 -311166
rect 100 -313554 112 -311178
rect 146 -313554 158 -311178
rect 100 -313566 158 -313554
rect -158 -313814 -100 -313802
rect -158 -316190 -146 -313814
rect -112 -316190 -100 -313814
rect -158 -316202 -100 -316190
rect 100 -313814 158 -313802
rect 100 -316190 112 -313814
rect 146 -316190 158 -313814
rect 100 -316202 158 -316190
rect -158 -316450 -100 -316438
rect -158 -318826 -146 -316450
rect -112 -318826 -100 -316450
rect -158 -318838 -100 -318826
rect 100 -316450 158 -316438
rect 100 -318826 112 -316450
rect 146 -318826 158 -316450
rect 100 -318838 158 -318826
rect -158 -319086 -100 -319074
rect -158 -321462 -146 -319086
rect -112 -321462 -100 -319086
rect -158 -321474 -100 -321462
rect 100 -319086 158 -319074
rect 100 -321462 112 -319086
rect 146 -321462 158 -319086
rect 100 -321474 158 -321462
rect -158 -321722 -100 -321710
rect -158 -324098 -146 -321722
rect -112 -324098 -100 -321722
rect -158 -324110 -100 -324098
rect 100 -321722 158 -321710
rect 100 -324098 112 -321722
rect 146 -324098 158 -321722
rect 100 -324110 158 -324098
rect -158 -324358 -100 -324346
rect -158 -326734 -146 -324358
rect -112 -326734 -100 -324358
rect -158 -326746 -100 -326734
rect 100 -324358 158 -324346
rect 100 -326734 112 -324358
rect 146 -326734 158 -324358
rect 100 -326746 158 -326734
rect -158 -326994 -100 -326982
rect -158 -329370 -146 -326994
rect -112 -329370 -100 -326994
rect -158 -329382 -100 -329370
rect 100 -326994 158 -326982
rect 100 -329370 112 -326994
rect 146 -329370 158 -326994
rect 100 -329382 158 -329370
rect -158 -329630 -100 -329618
rect -158 -332006 -146 -329630
rect -112 -332006 -100 -329630
rect -158 -332018 -100 -332006
rect 100 -329630 158 -329618
rect 100 -332006 112 -329630
rect 146 -332006 158 -329630
rect 100 -332018 158 -332006
rect -158 -332266 -100 -332254
rect -158 -334642 -146 -332266
rect -112 -334642 -100 -332266
rect -158 -334654 -100 -334642
rect 100 -332266 158 -332254
rect 100 -334642 112 -332266
rect 146 -334642 158 -332266
rect 100 -334654 158 -334642
rect -158 -334902 -100 -334890
rect -158 -337278 -146 -334902
rect -112 -337278 -100 -334902
rect -158 -337290 -100 -337278
rect 100 -334902 158 -334890
rect 100 -337278 112 -334902
rect 146 -337278 158 -334902
rect 100 -337290 158 -337278
<< mvpdiffc >>
rect -146 334902 -112 337278
rect 112 334902 146 337278
rect -146 332266 -112 334642
rect 112 332266 146 334642
rect -146 329630 -112 332006
rect 112 329630 146 332006
rect -146 326994 -112 329370
rect 112 326994 146 329370
rect -146 324358 -112 326734
rect 112 324358 146 326734
rect -146 321722 -112 324098
rect 112 321722 146 324098
rect -146 319086 -112 321462
rect 112 319086 146 321462
rect -146 316450 -112 318826
rect 112 316450 146 318826
rect -146 313814 -112 316190
rect 112 313814 146 316190
rect -146 311178 -112 313554
rect 112 311178 146 313554
rect -146 308542 -112 310918
rect 112 308542 146 310918
rect -146 305906 -112 308282
rect 112 305906 146 308282
rect -146 303270 -112 305646
rect 112 303270 146 305646
rect -146 300634 -112 303010
rect 112 300634 146 303010
rect -146 297998 -112 300374
rect 112 297998 146 300374
rect -146 295362 -112 297738
rect 112 295362 146 297738
rect -146 292726 -112 295102
rect 112 292726 146 295102
rect -146 290090 -112 292466
rect 112 290090 146 292466
rect -146 287454 -112 289830
rect 112 287454 146 289830
rect -146 284818 -112 287194
rect 112 284818 146 287194
rect -146 282182 -112 284558
rect 112 282182 146 284558
rect -146 279546 -112 281922
rect 112 279546 146 281922
rect -146 276910 -112 279286
rect 112 276910 146 279286
rect -146 274274 -112 276650
rect 112 274274 146 276650
rect -146 271638 -112 274014
rect 112 271638 146 274014
rect -146 269002 -112 271378
rect 112 269002 146 271378
rect -146 266366 -112 268742
rect 112 266366 146 268742
rect -146 263730 -112 266106
rect 112 263730 146 266106
rect -146 261094 -112 263470
rect 112 261094 146 263470
rect -146 258458 -112 260834
rect 112 258458 146 260834
rect -146 255822 -112 258198
rect 112 255822 146 258198
rect -146 253186 -112 255562
rect 112 253186 146 255562
rect -146 250550 -112 252926
rect 112 250550 146 252926
rect -146 247914 -112 250290
rect 112 247914 146 250290
rect -146 245278 -112 247654
rect 112 245278 146 247654
rect -146 242642 -112 245018
rect 112 242642 146 245018
rect -146 240006 -112 242382
rect 112 240006 146 242382
rect -146 237370 -112 239746
rect 112 237370 146 239746
rect -146 234734 -112 237110
rect 112 234734 146 237110
rect -146 232098 -112 234474
rect 112 232098 146 234474
rect -146 229462 -112 231838
rect 112 229462 146 231838
rect -146 226826 -112 229202
rect 112 226826 146 229202
rect -146 224190 -112 226566
rect 112 224190 146 226566
rect -146 221554 -112 223930
rect 112 221554 146 223930
rect -146 218918 -112 221294
rect 112 218918 146 221294
rect -146 216282 -112 218658
rect 112 216282 146 218658
rect -146 213646 -112 216022
rect 112 213646 146 216022
rect -146 211010 -112 213386
rect 112 211010 146 213386
rect -146 208374 -112 210750
rect 112 208374 146 210750
rect -146 205738 -112 208114
rect 112 205738 146 208114
rect -146 203102 -112 205478
rect 112 203102 146 205478
rect -146 200466 -112 202842
rect 112 200466 146 202842
rect -146 197830 -112 200206
rect 112 197830 146 200206
rect -146 195194 -112 197570
rect 112 195194 146 197570
rect -146 192558 -112 194934
rect 112 192558 146 194934
rect -146 189922 -112 192298
rect 112 189922 146 192298
rect -146 187286 -112 189662
rect 112 187286 146 189662
rect -146 184650 -112 187026
rect 112 184650 146 187026
rect -146 182014 -112 184390
rect 112 182014 146 184390
rect -146 179378 -112 181754
rect 112 179378 146 181754
rect -146 176742 -112 179118
rect 112 176742 146 179118
rect -146 174106 -112 176482
rect 112 174106 146 176482
rect -146 171470 -112 173846
rect 112 171470 146 173846
rect -146 168834 -112 171210
rect 112 168834 146 171210
rect -146 166198 -112 168574
rect 112 166198 146 168574
rect -146 163562 -112 165938
rect 112 163562 146 165938
rect -146 160926 -112 163302
rect 112 160926 146 163302
rect -146 158290 -112 160666
rect 112 158290 146 160666
rect -146 155654 -112 158030
rect 112 155654 146 158030
rect -146 153018 -112 155394
rect 112 153018 146 155394
rect -146 150382 -112 152758
rect 112 150382 146 152758
rect -146 147746 -112 150122
rect 112 147746 146 150122
rect -146 145110 -112 147486
rect 112 145110 146 147486
rect -146 142474 -112 144850
rect 112 142474 146 144850
rect -146 139838 -112 142214
rect 112 139838 146 142214
rect -146 137202 -112 139578
rect 112 137202 146 139578
rect -146 134566 -112 136942
rect 112 134566 146 136942
rect -146 131930 -112 134306
rect 112 131930 146 134306
rect -146 129294 -112 131670
rect 112 129294 146 131670
rect -146 126658 -112 129034
rect 112 126658 146 129034
rect -146 124022 -112 126398
rect 112 124022 146 126398
rect -146 121386 -112 123762
rect 112 121386 146 123762
rect -146 118750 -112 121126
rect 112 118750 146 121126
rect -146 116114 -112 118490
rect 112 116114 146 118490
rect -146 113478 -112 115854
rect 112 113478 146 115854
rect -146 110842 -112 113218
rect 112 110842 146 113218
rect -146 108206 -112 110582
rect 112 108206 146 110582
rect -146 105570 -112 107946
rect 112 105570 146 107946
rect -146 102934 -112 105310
rect 112 102934 146 105310
rect -146 100298 -112 102674
rect 112 100298 146 102674
rect -146 97662 -112 100038
rect 112 97662 146 100038
rect -146 95026 -112 97402
rect 112 95026 146 97402
rect -146 92390 -112 94766
rect 112 92390 146 94766
rect -146 89754 -112 92130
rect 112 89754 146 92130
rect -146 87118 -112 89494
rect 112 87118 146 89494
rect -146 84482 -112 86858
rect 112 84482 146 86858
rect -146 81846 -112 84222
rect 112 81846 146 84222
rect -146 79210 -112 81586
rect 112 79210 146 81586
rect -146 76574 -112 78950
rect 112 76574 146 78950
rect -146 73938 -112 76314
rect 112 73938 146 76314
rect -146 71302 -112 73678
rect 112 71302 146 73678
rect -146 68666 -112 71042
rect 112 68666 146 71042
rect -146 66030 -112 68406
rect 112 66030 146 68406
rect -146 63394 -112 65770
rect 112 63394 146 65770
rect -146 60758 -112 63134
rect 112 60758 146 63134
rect -146 58122 -112 60498
rect 112 58122 146 60498
rect -146 55486 -112 57862
rect 112 55486 146 57862
rect -146 52850 -112 55226
rect 112 52850 146 55226
rect -146 50214 -112 52590
rect 112 50214 146 52590
rect -146 47578 -112 49954
rect 112 47578 146 49954
rect -146 44942 -112 47318
rect 112 44942 146 47318
rect -146 42306 -112 44682
rect 112 42306 146 44682
rect -146 39670 -112 42046
rect 112 39670 146 42046
rect -146 37034 -112 39410
rect 112 37034 146 39410
rect -146 34398 -112 36774
rect 112 34398 146 36774
rect -146 31762 -112 34138
rect 112 31762 146 34138
rect -146 29126 -112 31502
rect 112 29126 146 31502
rect -146 26490 -112 28866
rect 112 26490 146 28866
rect -146 23854 -112 26230
rect 112 23854 146 26230
rect -146 21218 -112 23594
rect 112 21218 146 23594
rect -146 18582 -112 20958
rect 112 18582 146 20958
rect -146 15946 -112 18322
rect 112 15946 146 18322
rect -146 13310 -112 15686
rect 112 13310 146 15686
rect -146 10674 -112 13050
rect 112 10674 146 13050
rect -146 8038 -112 10414
rect 112 8038 146 10414
rect -146 5402 -112 7778
rect 112 5402 146 7778
rect -146 2766 -112 5142
rect 112 2766 146 5142
rect -146 130 -112 2506
rect 112 130 146 2506
rect -146 -2506 -112 -130
rect 112 -2506 146 -130
rect -146 -5142 -112 -2766
rect 112 -5142 146 -2766
rect -146 -7778 -112 -5402
rect 112 -7778 146 -5402
rect -146 -10414 -112 -8038
rect 112 -10414 146 -8038
rect -146 -13050 -112 -10674
rect 112 -13050 146 -10674
rect -146 -15686 -112 -13310
rect 112 -15686 146 -13310
rect -146 -18322 -112 -15946
rect 112 -18322 146 -15946
rect -146 -20958 -112 -18582
rect 112 -20958 146 -18582
rect -146 -23594 -112 -21218
rect 112 -23594 146 -21218
rect -146 -26230 -112 -23854
rect 112 -26230 146 -23854
rect -146 -28866 -112 -26490
rect 112 -28866 146 -26490
rect -146 -31502 -112 -29126
rect 112 -31502 146 -29126
rect -146 -34138 -112 -31762
rect 112 -34138 146 -31762
rect -146 -36774 -112 -34398
rect 112 -36774 146 -34398
rect -146 -39410 -112 -37034
rect 112 -39410 146 -37034
rect -146 -42046 -112 -39670
rect 112 -42046 146 -39670
rect -146 -44682 -112 -42306
rect 112 -44682 146 -42306
rect -146 -47318 -112 -44942
rect 112 -47318 146 -44942
rect -146 -49954 -112 -47578
rect 112 -49954 146 -47578
rect -146 -52590 -112 -50214
rect 112 -52590 146 -50214
rect -146 -55226 -112 -52850
rect 112 -55226 146 -52850
rect -146 -57862 -112 -55486
rect 112 -57862 146 -55486
rect -146 -60498 -112 -58122
rect 112 -60498 146 -58122
rect -146 -63134 -112 -60758
rect 112 -63134 146 -60758
rect -146 -65770 -112 -63394
rect 112 -65770 146 -63394
rect -146 -68406 -112 -66030
rect 112 -68406 146 -66030
rect -146 -71042 -112 -68666
rect 112 -71042 146 -68666
rect -146 -73678 -112 -71302
rect 112 -73678 146 -71302
rect -146 -76314 -112 -73938
rect 112 -76314 146 -73938
rect -146 -78950 -112 -76574
rect 112 -78950 146 -76574
rect -146 -81586 -112 -79210
rect 112 -81586 146 -79210
rect -146 -84222 -112 -81846
rect 112 -84222 146 -81846
rect -146 -86858 -112 -84482
rect 112 -86858 146 -84482
rect -146 -89494 -112 -87118
rect 112 -89494 146 -87118
rect -146 -92130 -112 -89754
rect 112 -92130 146 -89754
rect -146 -94766 -112 -92390
rect 112 -94766 146 -92390
rect -146 -97402 -112 -95026
rect 112 -97402 146 -95026
rect -146 -100038 -112 -97662
rect 112 -100038 146 -97662
rect -146 -102674 -112 -100298
rect 112 -102674 146 -100298
rect -146 -105310 -112 -102934
rect 112 -105310 146 -102934
rect -146 -107946 -112 -105570
rect 112 -107946 146 -105570
rect -146 -110582 -112 -108206
rect 112 -110582 146 -108206
rect -146 -113218 -112 -110842
rect 112 -113218 146 -110842
rect -146 -115854 -112 -113478
rect 112 -115854 146 -113478
rect -146 -118490 -112 -116114
rect 112 -118490 146 -116114
rect -146 -121126 -112 -118750
rect 112 -121126 146 -118750
rect -146 -123762 -112 -121386
rect 112 -123762 146 -121386
rect -146 -126398 -112 -124022
rect 112 -126398 146 -124022
rect -146 -129034 -112 -126658
rect 112 -129034 146 -126658
rect -146 -131670 -112 -129294
rect 112 -131670 146 -129294
rect -146 -134306 -112 -131930
rect 112 -134306 146 -131930
rect -146 -136942 -112 -134566
rect 112 -136942 146 -134566
rect -146 -139578 -112 -137202
rect 112 -139578 146 -137202
rect -146 -142214 -112 -139838
rect 112 -142214 146 -139838
rect -146 -144850 -112 -142474
rect 112 -144850 146 -142474
rect -146 -147486 -112 -145110
rect 112 -147486 146 -145110
rect -146 -150122 -112 -147746
rect 112 -150122 146 -147746
rect -146 -152758 -112 -150382
rect 112 -152758 146 -150382
rect -146 -155394 -112 -153018
rect 112 -155394 146 -153018
rect -146 -158030 -112 -155654
rect 112 -158030 146 -155654
rect -146 -160666 -112 -158290
rect 112 -160666 146 -158290
rect -146 -163302 -112 -160926
rect 112 -163302 146 -160926
rect -146 -165938 -112 -163562
rect 112 -165938 146 -163562
rect -146 -168574 -112 -166198
rect 112 -168574 146 -166198
rect -146 -171210 -112 -168834
rect 112 -171210 146 -168834
rect -146 -173846 -112 -171470
rect 112 -173846 146 -171470
rect -146 -176482 -112 -174106
rect 112 -176482 146 -174106
rect -146 -179118 -112 -176742
rect 112 -179118 146 -176742
rect -146 -181754 -112 -179378
rect 112 -181754 146 -179378
rect -146 -184390 -112 -182014
rect 112 -184390 146 -182014
rect -146 -187026 -112 -184650
rect 112 -187026 146 -184650
rect -146 -189662 -112 -187286
rect 112 -189662 146 -187286
rect -146 -192298 -112 -189922
rect 112 -192298 146 -189922
rect -146 -194934 -112 -192558
rect 112 -194934 146 -192558
rect -146 -197570 -112 -195194
rect 112 -197570 146 -195194
rect -146 -200206 -112 -197830
rect 112 -200206 146 -197830
rect -146 -202842 -112 -200466
rect 112 -202842 146 -200466
rect -146 -205478 -112 -203102
rect 112 -205478 146 -203102
rect -146 -208114 -112 -205738
rect 112 -208114 146 -205738
rect -146 -210750 -112 -208374
rect 112 -210750 146 -208374
rect -146 -213386 -112 -211010
rect 112 -213386 146 -211010
rect -146 -216022 -112 -213646
rect 112 -216022 146 -213646
rect -146 -218658 -112 -216282
rect 112 -218658 146 -216282
rect -146 -221294 -112 -218918
rect 112 -221294 146 -218918
rect -146 -223930 -112 -221554
rect 112 -223930 146 -221554
rect -146 -226566 -112 -224190
rect 112 -226566 146 -224190
rect -146 -229202 -112 -226826
rect 112 -229202 146 -226826
rect -146 -231838 -112 -229462
rect 112 -231838 146 -229462
rect -146 -234474 -112 -232098
rect 112 -234474 146 -232098
rect -146 -237110 -112 -234734
rect 112 -237110 146 -234734
rect -146 -239746 -112 -237370
rect 112 -239746 146 -237370
rect -146 -242382 -112 -240006
rect 112 -242382 146 -240006
rect -146 -245018 -112 -242642
rect 112 -245018 146 -242642
rect -146 -247654 -112 -245278
rect 112 -247654 146 -245278
rect -146 -250290 -112 -247914
rect 112 -250290 146 -247914
rect -146 -252926 -112 -250550
rect 112 -252926 146 -250550
rect -146 -255562 -112 -253186
rect 112 -255562 146 -253186
rect -146 -258198 -112 -255822
rect 112 -258198 146 -255822
rect -146 -260834 -112 -258458
rect 112 -260834 146 -258458
rect -146 -263470 -112 -261094
rect 112 -263470 146 -261094
rect -146 -266106 -112 -263730
rect 112 -266106 146 -263730
rect -146 -268742 -112 -266366
rect 112 -268742 146 -266366
rect -146 -271378 -112 -269002
rect 112 -271378 146 -269002
rect -146 -274014 -112 -271638
rect 112 -274014 146 -271638
rect -146 -276650 -112 -274274
rect 112 -276650 146 -274274
rect -146 -279286 -112 -276910
rect 112 -279286 146 -276910
rect -146 -281922 -112 -279546
rect 112 -281922 146 -279546
rect -146 -284558 -112 -282182
rect 112 -284558 146 -282182
rect -146 -287194 -112 -284818
rect 112 -287194 146 -284818
rect -146 -289830 -112 -287454
rect 112 -289830 146 -287454
rect -146 -292466 -112 -290090
rect 112 -292466 146 -290090
rect -146 -295102 -112 -292726
rect 112 -295102 146 -292726
rect -146 -297738 -112 -295362
rect 112 -297738 146 -295362
rect -146 -300374 -112 -297998
rect 112 -300374 146 -297998
rect -146 -303010 -112 -300634
rect 112 -303010 146 -300634
rect -146 -305646 -112 -303270
rect 112 -305646 146 -303270
rect -146 -308282 -112 -305906
rect 112 -308282 146 -305906
rect -146 -310918 -112 -308542
rect 112 -310918 146 -308542
rect -146 -313554 -112 -311178
rect 112 -313554 146 -311178
rect -146 -316190 -112 -313814
rect 112 -316190 146 -313814
rect -146 -318826 -112 -316450
rect 112 -318826 146 -316450
rect -146 -321462 -112 -319086
rect 112 -321462 146 -319086
rect -146 -324098 -112 -321722
rect 112 -324098 146 -321722
rect -146 -326734 -112 -324358
rect 112 -326734 146 -324358
rect -146 -329370 -112 -326994
rect 112 -329370 146 -326994
rect -146 -332006 -112 -329630
rect 112 -332006 146 -329630
rect -146 -334642 -112 -332266
rect 112 -334642 146 -332266
rect -146 -337278 -112 -334902
rect 112 -337278 146 -334902
<< mvnsubdiff >>
rect -292 337509 292 337521
rect -292 337475 -184 337509
rect 184 337475 292 337509
rect -292 337463 292 337475
rect -292 337413 -234 337463
rect -292 -337413 -280 337413
rect -246 -337413 -234 337413
rect 234 337413 292 337463
rect -292 -337463 -234 -337413
rect 234 -337413 246 337413
rect 280 -337413 292 337413
rect 234 -337463 292 -337413
rect -292 -337475 292 -337463
rect -292 -337509 -184 -337475
rect 184 -337509 292 -337475
rect -292 -337521 292 -337509
<< mvnsubdiffcont >>
rect -184 337475 184 337509
rect -280 -337413 -246 337413
rect 246 -337413 280 337413
rect -184 -337509 184 -337475
<< poly >>
rect -100 337371 100 337387
rect -100 337337 -84 337371
rect 84 337337 100 337371
rect -100 337290 100 337337
rect -100 334843 100 334890
rect -100 334809 -84 334843
rect 84 334809 100 334843
rect -100 334793 100 334809
rect -100 334735 100 334751
rect -100 334701 -84 334735
rect 84 334701 100 334735
rect -100 334654 100 334701
rect -100 332207 100 332254
rect -100 332173 -84 332207
rect 84 332173 100 332207
rect -100 332157 100 332173
rect -100 332099 100 332115
rect -100 332065 -84 332099
rect 84 332065 100 332099
rect -100 332018 100 332065
rect -100 329571 100 329618
rect -100 329537 -84 329571
rect 84 329537 100 329571
rect -100 329521 100 329537
rect -100 329463 100 329479
rect -100 329429 -84 329463
rect 84 329429 100 329463
rect -100 329382 100 329429
rect -100 326935 100 326982
rect -100 326901 -84 326935
rect 84 326901 100 326935
rect -100 326885 100 326901
rect -100 326827 100 326843
rect -100 326793 -84 326827
rect 84 326793 100 326827
rect -100 326746 100 326793
rect -100 324299 100 324346
rect -100 324265 -84 324299
rect 84 324265 100 324299
rect -100 324249 100 324265
rect -100 324191 100 324207
rect -100 324157 -84 324191
rect 84 324157 100 324191
rect -100 324110 100 324157
rect -100 321663 100 321710
rect -100 321629 -84 321663
rect 84 321629 100 321663
rect -100 321613 100 321629
rect -100 321555 100 321571
rect -100 321521 -84 321555
rect 84 321521 100 321555
rect -100 321474 100 321521
rect -100 319027 100 319074
rect -100 318993 -84 319027
rect 84 318993 100 319027
rect -100 318977 100 318993
rect -100 318919 100 318935
rect -100 318885 -84 318919
rect 84 318885 100 318919
rect -100 318838 100 318885
rect -100 316391 100 316438
rect -100 316357 -84 316391
rect 84 316357 100 316391
rect -100 316341 100 316357
rect -100 316283 100 316299
rect -100 316249 -84 316283
rect 84 316249 100 316283
rect -100 316202 100 316249
rect -100 313755 100 313802
rect -100 313721 -84 313755
rect 84 313721 100 313755
rect -100 313705 100 313721
rect -100 313647 100 313663
rect -100 313613 -84 313647
rect 84 313613 100 313647
rect -100 313566 100 313613
rect -100 311119 100 311166
rect -100 311085 -84 311119
rect 84 311085 100 311119
rect -100 311069 100 311085
rect -100 311011 100 311027
rect -100 310977 -84 311011
rect 84 310977 100 311011
rect -100 310930 100 310977
rect -100 308483 100 308530
rect -100 308449 -84 308483
rect 84 308449 100 308483
rect -100 308433 100 308449
rect -100 308375 100 308391
rect -100 308341 -84 308375
rect 84 308341 100 308375
rect -100 308294 100 308341
rect -100 305847 100 305894
rect -100 305813 -84 305847
rect 84 305813 100 305847
rect -100 305797 100 305813
rect -100 305739 100 305755
rect -100 305705 -84 305739
rect 84 305705 100 305739
rect -100 305658 100 305705
rect -100 303211 100 303258
rect -100 303177 -84 303211
rect 84 303177 100 303211
rect -100 303161 100 303177
rect -100 303103 100 303119
rect -100 303069 -84 303103
rect 84 303069 100 303103
rect -100 303022 100 303069
rect -100 300575 100 300622
rect -100 300541 -84 300575
rect 84 300541 100 300575
rect -100 300525 100 300541
rect -100 300467 100 300483
rect -100 300433 -84 300467
rect 84 300433 100 300467
rect -100 300386 100 300433
rect -100 297939 100 297986
rect -100 297905 -84 297939
rect 84 297905 100 297939
rect -100 297889 100 297905
rect -100 297831 100 297847
rect -100 297797 -84 297831
rect 84 297797 100 297831
rect -100 297750 100 297797
rect -100 295303 100 295350
rect -100 295269 -84 295303
rect 84 295269 100 295303
rect -100 295253 100 295269
rect -100 295195 100 295211
rect -100 295161 -84 295195
rect 84 295161 100 295195
rect -100 295114 100 295161
rect -100 292667 100 292714
rect -100 292633 -84 292667
rect 84 292633 100 292667
rect -100 292617 100 292633
rect -100 292559 100 292575
rect -100 292525 -84 292559
rect 84 292525 100 292559
rect -100 292478 100 292525
rect -100 290031 100 290078
rect -100 289997 -84 290031
rect 84 289997 100 290031
rect -100 289981 100 289997
rect -100 289923 100 289939
rect -100 289889 -84 289923
rect 84 289889 100 289923
rect -100 289842 100 289889
rect -100 287395 100 287442
rect -100 287361 -84 287395
rect 84 287361 100 287395
rect -100 287345 100 287361
rect -100 287287 100 287303
rect -100 287253 -84 287287
rect 84 287253 100 287287
rect -100 287206 100 287253
rect -100 284759 100 284806
rect -100 284725 -84 284759
rect 84 284725 100 284759
rect -100 284709 100 284725
rect -100 284651 100 284667
rect -100 284617 -84 284651
rect 84 284617 100 284651
rect -100 284570 100 284617
rect -100 282123 100 282170
rect -100 282089 -84 282123
rect 84 282089 100 282123
rect -100 282073 100 282089
rect -100 282015 100 282031
rect -100 281981 -84 282015
rect 84 281981 100 282015
rect -100 281934 100 281981
rect -100 279487 100 279534
rect -100 279453 -84 279487
rect 84 279453 100 279487
rect -100 279437 100 279453
rect -100 279379 100 279395
rect -100 279345 -84 279379
rect 84 279345 100 279379
rect -100 279298 100 279345
rect -100 276851 100 276898
rect -100 276817 -84 276851
rect 84 276817 100 276851
rect -100 276801 100 276817
rect -100 276743 100 276759
rect -100 276709 -84 276743
rect 84 276709 100 276743
rect -100 276662 100 276709
rect -100 274215 100 274262
rect -100 274181 -84 274215
rect 84 274181 100 274215
rect -100 274165 100 274181
rect -100 274107 100 274123
rect -100 274073 -84 274107
rect 84 274073 100 274107
rect -100 274026 100 274073
rect -100 271579 100 271626
rect -100 271545 -84 271579
rect 84 271545 100 271579
rect -100 271529 100 271545
rect -100 271471 100 271487
rect -100 271437 -84 271471
rect 84 271437 100 271471
rect -100 271390 100 271437
rect -100 268943 100 268990
rect -100 268909 -84 268943
rect 84 268909 100 268943
rect -100 268893 100 268909
rect -100 268835 100 268851
rect -100 268801 -84 268835
rect 84 268801 100 268835
rect -100 268754 100 268801
rect -100 266307 100 266354
rect -100 266273 -84 266307
rect 84 266273 100 266307
rect -100 266257 100 266273
rect -100 266199 100 266215
rect -100 266165 -84 266199
rect 84 266165 100 266199
rect -100 266118 100 266165
rect -100 263671 100 263718
rect -100 263637 -84 263671
rect 84 263637 100 263671
rect -100 263621 100 263637
rect -100 263563 100 263579
rect -100 263529 -84 263563
rect 84 263529 100 263563
rect -100 263482 100 263529
rect -100 261035 100 261082
rect -100 261001 -84 261035
rect 84 261001 100 261035
rect -100 260985 100 261001
rect -100 260927 100 260943
rect -100 260893 -84 260927
rect 84 260893 100 260927
rect -100 260846 100 260893
rect -100 258399 100 258446
rect -100 258365 -84 258399
rect 84 258365 100 258399
rect -100 258349 100 258365
rect -100 258291 100 258307
rect -100 258257 -84 258291
rect 84 258257 100 258291
rect -100 258210 100 258257
rect -100 255763 100 255810
rect -100 255729 -84 255763
rect 84 255729 100 255763
rect -100 255713 100 255729
rect -100 255655 100 255671
rect -100 255621 -84 255655
rect 84 255621 100 255655
rect -100 255574 100 255621
rect -100 253127 100 253174
rect -100 253093 -84 253127
rect 84 253093 100 253127
rect -100 253077 100 253093
rect -100 253019 100 253035
rect -100 252985 -84 253019
rect 84 252985 100 253019
rect -100 252938 100 252985
rect -100 250491 100 250538
rect -100 250457 -84 250491
rect 84 250457 100 250491
rect -100 250441 100 250457
rect -100 250383 100 250399
rect -100 250349 -84 250383
rect 84 250349 100 250383
rect -100 250302 100 250349
rect -100 247855 100 247902
rect -100 247821 -84 247855
rect 84 247821 100 247855
rect -100 247805 100 247821
rect -100 247747 100 247763
rect -100 247713 -84 247747
rect 84 247713 100 247747
rect -100 247666 100 247713
rect -100 245219 100 245266
rect -100 245185 -84 245219
rect 84 245185 100 245219
rect -100 245169 100 245185
rect -100 245111 100 245127
rect -100 245077 -84 245111
rect 84 245077 100 245111
rect -100 245030 100 245077
rect -100 242583 100 242630
rect -100 242549 -84 242583
rect 84 242549 100 242583
rect -100 242533 100 242549
rect -100 242475 100 242491
rect -100 242441 -84 242475
rect 84 242441 100 242475
rect -100 242394 100 242441
rect -100 239947 100 239994
rect -100 239913 -84 239947
rect 84 239913 100 239947
rect -100 239897 100 239913
rect -100 239839 100 239855
rect -100 239805 -84 239839
rect 84 239805 100 239839
rect -100 239758 100 239805
rect -100 237311 100 237358
rect -100 237277 -84 237311
rect 84 237277 100 237311
rect -100 237261 100 237277
rect -100 237203 100 237219
rect -100 237169 -84 237203
rect 84 237169 100 237203
rect -100 237122 100 237169
rect -100 234675 100 234722
rect -100 234641 -84 234675
rect 84 234641 100 234675
rect -100 234625 100 234641
rect -100 234567 100 234583
rect -100 234533 -84 234567
rect 84 234533 100 234567
rect -100 234486 100 234533
rect -100 232039 100 232086
rect -100 232005 -84 232039
rect 84 232005 100 232039
rect -100 231989 100 232005
rect -100 231931 100 231947
rect -100 231897 -84 231931
rect 84 231897 100 231931
rect -100 231850 100 231897
rect -100 229403 100 229450
rect -100 229369 -84 229403
rect 84 229369 100 229403
rect -100 229353 100 229369
rect -100 229295 100 229311
rect -100 229261 -84 229295
rect 84 229261 100 229295
rect -100 229214 100 229261
rect -100 226767 100 226814
rect -100 226733 -84 226767
rect 84 226733 100 226767
rect -100 226717 100 226733
rect -100 226659 100 226675
rect -100 226625 -84 226659
rect 84 226625 100 226659
rect -100 226578 100 226625
rect -100 224131 100 224178
rect -100 224097 -84 224131
rect 84 224097 100 224131
rect -100 224081 100 224097
rect -100 224023 100 224039
rect -100 223989 -84 224023
rect 84 223989 100 224023
rect -100 223942 100 223989
rect -100 221495 100 221542
rect -100 221461 -84 221495
rect 84 221461 100 221495
rect -100 221445 100 221461
rect -100 221387 100 221403
rect -100 221353 -84 221387
rect 84 221353 100 221387
rect -100 221306 100 221353
rect -100 218859 100 218906
rect -100 218825 -84 218859
rect 84 218825 100 218859
rect -100 218809 100 218825
rect -100 218751 100 218767
rect -100 218717 -84 218751
rect 84 218717 100 218751
rect -100 218670 100 218717
rect -100 216223 100 216270
rect -100 216189 -84 216223
rect 84 216189 100 216223
rect -100 216173 100 216189
rect -100 216115 100 216131
rect -100 216081 -84 216115
rect 84 216081 100 216115
rect -100 216034 100 216081
rect -100 213587 100 213634
rect -100 213553 -84 213587
rect 84 213553 100 213587
rect -100 213537 100 213553
rect -100 213479 100 213495
rect -100 213445 -84 213479
rect 84 213445 100 213479
rect -100 213398 100 213445
rect -100 210951 100 210998
rect -100 210917 -84 210951
rect 84 210917 100 210951
rect -100 210901 100 210917
rect -100 210843 100 210859
rect -100 210809 -84 210843
rect 84 210809 100 210843
rect -100 210762 100 210809
rect -100 208315 100 208362
rect -100 208281 -84 208315
rect 84 208281 100 208315
rect -100 208265 100 208281
rect -100 208207 100 208223
rect -100 208173 -84 208207
rect 84 208173 100 208207
rect -100 208126 100 208173
rect -100 205679 100 205726
rect -100 205645 -84 205679
rect 84 205645 100 205679
rect -100 205629 100 205645
rect -100 205571 100 205587
rect -100 205537 -84 205571
rect 84 205537 100 205571
rect -100 205490 100 205537
rect -100 203043 100 203090
rect -100 203009 -84 203043
rect 84 203009 100 203043
rect -100 202993 100 203009
rect -100 202935 100 202951
rect -100 202901 -84 202935
rect 84 202901 100 202935
rect -100 202854 100 202901
rect -100 200407 100 200454
rect -100 200373 -84 200407
rect 84 200373 100 200407
rect -100 200357 100 200373
rect -100 200299 100 200315
rect -100 200265 -84 200299
rect 84 200265 100 200299
rect -100 200218 100 200265
rect -100 197771 100 197818
rect -100 197737 -84 197771
rect 84 197737 100 197771
rect -100 197721 100 197737
rect -100 197663 100 197679
rect -100 197629 -84 197663
rect 84 197629 100 197663
rect -100 197582 100 197629
rect -100 195135 100 195182
rect -100 195101 -84 195135
rect 84 195101 100 195135
rect -100 195085 100 195101
rect -100 195027 100 195043
rect -100 194993 -84 195027
rect 84 194993 100 195027
rect -100 194946 100 194993
rect -100 192499 100 192546
rect -100 192465 -84 192499
rect 84 192465 100 192499
rect -100 192449 100 192465
rect -100 192391 100 192407
rect -100 192357 -84 192391
rect 84 192357 100 192391
rect -100 192310 100 192357
rect -100 189863 100 189910
rect -100 189829 -84 189863
rect 84 189829 100 189863
rect -100 189813 100 189829
rect -100 189755 100 189771
rect -100 189721 -84 189755
rect 84 189721 100 189755
rect -100 189674 100 189721
rect -100 187227 100 187274
rect -100 187193 -84 187227
rect 84 187193 100 187227
rect -100 187177 100 187193
rect -100 187119 100 187135
rect -100 187085 -84 187119
rect 84 187085 100 187119
rect -100 187038 100 187085
rect -100 184591 100 184638
rect -100 184557 -84 184591
rect 84 184557 100 184591
rect -100 184541 100 184557
rect -100 184483 100 184499
rect -100 184449 -84 184483
rect 84 184449 100 184483
rect -100 184402 100 184449
rect -100 181955 100 182002
rect -100 181921 -84 181955
rect 84 181921 100 181955
rect -100 181905 100 181921
rect -100 181847 100 181863
rect -100 181813 -84 181847
rect 84 181813 100 181847
rect -100 181766 100 181813
rect -100 179319 100 179366
rect -100 179285 -84 179319
rect 84 179285 100 179319
rect -100 179269 100 179285
rect -100 179211 100 179227
rect -100 179177 -84 179211
rect 84 179177 100 179211
rect -100 179130 100 179177
rect -100 176683 100 176730
rect -100 176649 -84 176683
rect 84 176649 100 176683
rect -100 176633 100 176649
rect -100 176575 100 176591
rect -100 176541 -84 176575
rect 84 176541 100 176575
rect -100 176494 100 176541
rect -100 174047 100 174094
rect -100 174013 -84 174047
rect 84 174013 100 174047
rect -100 173997 100 174013
rect -100 173939 100 173955
rect -100 173905 -84 173939
rect 84 173905 100 173939
rect -100 173858 100 173905
rect -100 171411 100 171458
rect -100 171377 -84 171411
rect 84 171377 100 171411
rect -100 171361 100 171377
rect -100 171303 100 171319
rect -100 171269 -84 171303
rect 84 171269 100 171303
rect -100 171222 100 171269
rect -100 168775 100 168822
rect -100 168741 -84 168775
rect 84 168741 100 168775
rect -100 168725 100 168741
rect -100 168667 100 168683
rect -100 168633 -84 168667
rect 84 168633 100 168667
rect -100 168586 100 168633
rect -100 166139 100 166186
rect -100 166105 -84 166139
rect 84 166105 100 166139
rect -100 166089 100 166105
rect -100 166031 100 166047
rect -100 165997 -84 166031
rect 84 165997 100 166031
rect -100 165950 100 165997
rect -100 163503 100 163550
rect -100 163469 -84 163503
rect 84 163469 100 163503
rect -100 163453 100 163469
rect -100 163395 100 163411
rect -100 163361 -84 163395
rect 84 163361 100 163395
rect -100 163314 100 163361
rect -100 160867 100 160914
rect -100 160833 -84 160867
rect 84 160833 100 160867
rect -100 160817 100 160833
rect -100 160759 100 160775
rect -100 160725 -84 160759
rect 84 160725 100 160759
rect -100 160678 100 160725
rect -100 158231 100 158278
rect -100 158197 -84 158231
rect 84 158197 100 158231
rect -100 158181 100 158197
rect -100 158123 100 158139
rect -100 158089 -84 158123
rect 84 158089 100 158123
rect -100 158042 100 158089
rect -100 155595 100 155642
rect -100 155561 -84 155595
rect 84 155561 100 155595
rect -100 155545 100 155561
rect -100 155487 100 155503
rect -100 155453 -84 155487
rect 84 155453 100 155487
rect -100 155406 100 155453
rect -100 152959 100 153006
rect -100 152925 -84 152959
rect 84 152925 100 152959
rect -100 152909 100 152925
rect -100 152851 100 152867
rect -100 152817 -84 152851
rect 84 152817 100 152851
rect -100 152770 100 152817
rect -100 150323 100 150370
rect -100 150289 -84 150323
rect 84 150289 100 150323
rect -100 150273 100 150289
rect -100 150215 100 150231
rect -100 150181 -84 150215
rect 84 150181 100 150215
rect -100 150134 100 150181
rect -100 147687 100 147734
rect -100 147653 -84 147687
rect 84 147653 100 147687
rect -100 147637 100 147653
rect -100 147579 100 147595
rect -100 147545 -84 147579
rect 84 147545 100 147579
rect -100 147498 100 147545
rect -100 145051 100 145098
rect -100 145017 -84 145051
rect 84 145017 100 145051
rect -100 145001 100 145017
rect -100 144943 100 144959
rect -100 144909 -84 144943
rect 84 144909 100 144943
rect -100 144862 100 144909
rect -100 142415 100 142462
rect -100 142381 -84 142415
rect 84 142381 100 142415
rect -100 142365 100 142381
rect -100 142307 100 142323
rect -100 142273 -84 142307
rect 84 142273 100 142307
rect -100 142226 100 142273
rect -100 139779 100 139826
rect -100 139745 -84 139779
rect 84 139745 100 139779
rect -100 139729 100 139745
rect -100 139671 100 139687
rect -100 139637 -84 139671
rect 84 139637 100 139671
rect -100 139590 100 139637
rect -100 137143 100 137190
rect -100 137109 -84 137143
rect 84 137109 100 137143
rect -100 137093 100 137109
rect -100 137035 100 137051
rect -100 137001 -84 137035
rect 84 137001 100 137035
rect -100 136954 100 137001
rect -100 134507 100 134554
rect -100 134473 -84 134507
rect 84 134473 100 134507
rect -100 134457 100 134473
rect -100 134399 100 134415
rect -100 134365 -84 134399
rect 84 134365 100 134399
rect -100 134318 100 134365
rect -100 131871 100 131918
rect -100 131837 -84 131871
rect 84 131837 100 131871
rect -100 131821 100 131837
rect -100 131763 100 131779
rect -100 131729 -84 131763
rect 84 131729 100 131763
rect -100 131682 100 131729
rect -100 129235 100 129282
rect -100 129201 -84 129235
rect 84 129201 100 129235
rect -100 129185 100 129201
rect -100 129127 100 129143
rect -100 129093 -84 129127
rect 84 129093 100 129127
rect -100 129046 100 129093
rect -100 126599 100 126646
rect -100 126565 -84 126599
rect 84 126565 100 126599
rect -100 126549 100 126565
rect -100 126491 100 126507
rect -100 126457 -84 126491
rect 84 126457 100 126491
rect -100 126410 100 126457
rect -100 123963 100 124010
rect -100 123929 -84 123963
rect 84 123929 100 123963
rect -100 123913 100 123929
rect -100 123855 100 123871
rect -100 123821 -84 123855
rect 84 123821 100 123855
rect -100 123774 100 123821
rect -100 121327 100 121374
rect -100 121293 -84 121327
rect 84 121293 100 121327
rect -100 121277 100 121293
rect -100 121219 100 121235
rect -100 121185 -84 121219
rect 84 121185 100 121219
rect -100 121138 100 121185
rect -100 118691 100 118738
rect -100 118657 -84 118691
rect 84 118657 100 118691
rect -100 118641 100 118657
rect -100 118583 100 118599
rect -100 118549 -84 118583
rect 84 118549 100 118583
rect -100 118502 100 118549
rect -100 116055 100 116102
rect -100 116021 -84 116055
rect 84 116021 100 116055
rect -100 116005 100 116021
rect -100 115947 100 115963
rect -100 115913 -84 115947
rect 84 115913 100 115947
rect -100 115866 100 115913
rect -100 113419 100 113466
rect -100 113385 -84 113419
rect 84 113385 100 113419
rect -100 113369 100 113385
rect -100 113311 100 113327
rect -100 113277 -84 113311
rect 84 113277 100 113311
rect -100 113230 100 113277
rect -100 110783 100 110830
rect -100 110749 -84 110783
rect 84 110749 100 110783
rect -100 110733 100 110749
rect -100 110675 100 110691
rect -100 110641 -84 110675
rect 84 110641 100 110675
rect -100 110594 100 110641
rect -100 108147 100 108194
rect -100 108113 -84 108147
rect 84 108113 100 108147
rect -100 108097 100 108113
rect -100 108039 100 108055
rect -100 108005 -84 108039
rect 84 108005 100 108039
rect -100 107958 100 108005
rect -100 105511 100 105558
rect -100 105477 -84 105511
rect 84 105477 100 105511
rect -100 105461 100 105477
rect -100 105403 100 105419
rect -100 105369 -84 105403
rect 84 105369 100 105403
rect -100 105322 100 105369
rect -100 102875 100 102922
rect -100 102841 -84 102875
rect 84 102841 100 102875
rect -100 102825 100 102841
rect -100 102767 100 102783
rect -100 102733 -84 102767
rect 84 102733 100 102767
rect -100 102686 100 102733
rect -100 100239 100 100286
rect -100 100205 -84 100239
rect 84 100205 100 100239
rect -100 100189 100 100205
rect -100 100131 100 100147
rect -100 100097 -84 100131
rect 84 100097 100 100131
rect -100 100050 100 100097
rect -100 97603 100 97650
rect -100 97569 -84 97603
rect 84 97569 100 97603
rect -100 97553 100 97569
rect -100 97495 100 97511
rect -100 97461 -84 97495
rect 84 97461 100 97495
rect -100 97414 100 97461
rect -100 94967 100 95014
rect -100 94933 -84 94967
rect 84 94933 100 94967
rect -100 94917 100 94933
rect -100 94859 100 94875
rect -100 94825 -84 94859
rect 84 94825 100 94859
rect -100 94778 100 94825
rect -100 92331 100 92378
rect -100 92297 -84 92331
rect 84 92297 100 92331
rect -100 92281 100 92297
rect -100 92223 100 92239
rect -100 92189 -84 92223
rect 84 92189 100 92223
rect -100 92142 100 92189
rect -100 89695 100 89742
rect -100 89661 -84 89695
rect 84 89661 100 89695
rect -100 89645 100 89661
rect -100 89587 100 89603
rect -100 89553 -84 89587
rect 84 89553 100 89587
rect -100 89506 100 89553
rect -100 87059 100 87106
rect -100 87025 -84 87059
rect 84 87025 100 87059
rect -100 87009 100 87025
rect -100 86951 100 86967
rect -100 86917 -84 86951
rect 84 86917 100 86951
rect -100 86870 100 86917
rect -100 84423 100 84470
rect -100 84389 -84 84423
rect 84 84389 100 84423
rect -100 84373 100 84389
rect -100 84315 100 84331
rect -100 84281 -84 84315
rect 84 84281 100 84315
rect -100 84234 100 84281
rect -100 81787 100 81834
rect -100 81753 -84 81787
rect 84 81753 100 81787
rect -100 81737 100 81753
rect -100 81679 100 81695
rect -100 81645 -84 81679
rect 84 81645 100 81679
rect -100 81598 100 81645
rect -100 79151 100 79198
rect -100 79117 -84 79151
rect 84 79117 100 79151
rect -100 79101 100 79117
rect -100 79043 100 79059
rect -100 79009 -84 79043
rect 84 79009 100 79043
rect -100 78962 100 79009
rect -100 76515 100 76562
rect -100 76481 -84 76515
rect 84 76481 100 76515
rect -100 76465 100 76481
rect -100 76407 100 76423
rect -100 76373 -84 76407
rect 84 76373 100 76407
rect -100 76326 100 76373
rect -100 73879 100 73926
rect -100 73845 -84 73879
rect 84 73845 100 73879
rect -100 73829 100 73845
rect -100 73771 100 73787
rect -100 73737 -84 73771
rect 84 73737 100 73771
rect -100 73690 100 73737
rect -100 71243 100 71290
rect -100 71209 -84 71243
rect 84 71209 100 71243
rect -100 71193 100 71209
rect -100 71135 100 71151
rect -100 71101 -84 71135
rect 84 71101 100 71135
rect -100 71054 100 71101
rect -100 68607 100 68654
rect -100 68573 -84 68607
rect 84 68573 100 68607
rect -100 68557 100 68573
rect -100 68499 100 68515
rect -100 68465 -84 68499
rect 84 68465 100 68499
rect -100 68418 100 68465
rect -100 65971 100 66018
rect -100 65937 -84 65971
rect 84 65937 100 65971
rect -100 65921 100 65937
rect -100 65863 100 65879
rect -100 65829 -84 65863
rect 84 65829 100 65863
rect -100 65782 100 65829
rect -100 63335 100 63382
rect -100 63301 -84 63335
rect 84 63301 100 63335
rect -100 63285 100 63301
rect -100 63227 100 63243
rect -100 63193 -84 63227
rect 84 63193 100 63227
rect -100 63146 100 63193
rect -100 60699 100 60746
rect -100 60665 -84 60699
rect 84 60665 100 60699
rect -100 60649 100 60665
rect -100 60591 100 60607
rect -100 60557 -84 60591
rect 84 60557 100 60591
rect -100 60510 100 60557
rect -100 58063 100 58110
rect -100 58029 -84 58063
rect 84 58029 100 58063
rect -100 58013 100 58029
rect -100 57955 100 57971
rect -100 57921 -84 57955
rect 84 57921 100 57955
rect -100 57874 100 57921
rect -100 55427 100 55474
rect -100 55393 -84 55427
rect 84 55393 100 55427
rect -100 55377 100 55393
rect -100 55319 100 55335
rect -100 55285 -84 55319
rect 84 55285 100 55319
rect -100 55238 100 55285
rect -100 52791 100 52838
rect -100 52757 -84 52791
rect 84 52757 100 52791
rect -100 52741 100 52757
rect -100 52683 100 52699
rect -100 52649 -84 52683
rect 84 52649 100 52683
rect -100 52602 100 52649
rect -100 50155 100 50202
rect -100 50121 -84 50155
rect 84 50121 100 50155
rect -100 50105 100 50121
rect -100 50047 100 50063
rect -100 50013 -84 50047
rect 84 50013 100 50047
rect -100 49966 100 50013
rect -100 47519 100 47566
rect -100 47485 -84 47519
rect 84 47485 100 47519
rect -100 47469 100 47485
rect -100 47411 100 47427
rect -100 47377 -84 47411
rect 84 47377 100 47411
rect -100 47330 100 47377
rect -100 44883 100 44930
rect -100 44849 -84 44883
rect 84 44849 100 44883
rect -100 44833 100 44849
rect -100 44775 100 44791
rect -100 44741 -84 44775
rect 84 44741 100 44775
rect -100 44694 100 44741
rect -100 42247 100 42294
rect -100 42213 -84 42247
rect 84 42213 100 42247
rect -100 42197 100 42213
rect -100 42139 100 42155
rect -100 42105 -84 42139
rect 84 42105 100 42139
rect -100 42058 100 42105
rect -100 39611 100 39658
rect -100 39577 -84 39611
rect 84 39577 100 39611
rect -100 39561 100 39577
rect -100 39503 100 39519
rect -100 39469 -84 39503
rect 84 39469 100 39503
rect -100 39422 100 39469
rect -100 36975 100 37022
rect -100 36941 -84 36975
rect 84 36941 100 36975
rect -100 36925 100 36941
rect -100 36867 100 36883
rect -100 36833 -84 36867
rect 84 36833 100 36867
rect -100 36786 100 36833
rect -100 34339 100 34386
rect -100 34305 -84 34339
rect 84 34305 100 34339
rect -100 34289 100 34305
rect -100 34231 100 34247
rect -100 34197 -84 34231
rect 84 34197 100 34231
rect -100 34150 100 34197
rect -100 31703 100 31750
rect -100 31669 -84 31703
rect 84 31669 100 31703
rect -100 31653 100 31669
rect -100 31595 100 31611
rect -100 31561 -84 31595
rect 84 31561 100 31595
rect -100 31514 100 31561
rect -100 29067 100 29114
rect -100 29033 -84 29067
rect 84 29033 100 29067
rect -100 29017 100 29033
rect -100 28959 100 28975
rect -100 28925 -84 28959
rect 84 28925 100 28959
rect -100 28878 100 28925
rect -100 26431 100 26478
rect -100 26397 -84 26431
rect 84 26397 100 26431
rect -100 26381 100 26397
rect -100 26323 100 26339
rect -100 26289 -84 26323
rect 84 26289 100 26323
rect -100 26242 100 26289
rect -100 23795 100 23842
rect -100 23761 -84 23795
rect 84 23761 100 23795
rect -100 23745 100 23761
rect -100 23687 100 23703
rect -100 23653 -84 23687
rect 84 23653 100 23687
rect -100 23606 100 23653
rect -100 21159 100 21206
rect -100 21125 -84 21159
rect 84 21125 100 21159
rect -100 21109 100 21125
rect -100 21051 100 21067
rect -100 21017 -84 21051
rect 84 21017 100 21051
rect -100 20970 100 21017
rect -100 18523 100 18570
rect -100 18489 -84 18523
rect 84 18489 100 18523
rect -100 18473 100 18489
rect -100 18415 100 18431
rect -100 18381 -84 18415
rect 84 18381 100 18415
rect -100 18334 100 18381
rect -100 15887 100 15934
rect -100 15853 -84 15887
rect 84 15853 100 15887
rect -100 15837 100 15853
rect -100 15779 100 15795
rect -100 15745 -84 15779
rect 84 15745 100 15779
rect -100 15698 100 15745
rect -100 13251 100 13298
rect -100 13217 -84 13251
rect 84 13217 100 13251
rect -100 13201 100 13217
rect -100 13143 100 13159
rect -100 13109 -84 13143
rect 84 13109 100 13143
rect -100 13062 100 13109
rect -100 10615 100 10662
rect -100 10581 -84 10615
rect 84 10581 100 10615
rect -100 10565 100 10581
rect -100 10507 100 10523
rect -100 10473 -84 10507
rect 84 10473 100 10507
rect -100 10426 100 10473
rect -100 7979 100 8026
rect -100 7945 -84 7979
rect 84 7945 100 7979
rect -100 7929 100 7945
rect -100 7871 100 7887
rect -100 7837 -84 7871
rect 84 7837 100 7871
rect -100 7790 100 7837
rect -100 5343 100 5390
rect -100 5309 -84 5343
rect 84 5309 100 5343
rect -100 5293 100 5309
rect -100 5235 100 5251
rect -100 5201 -84 5235
rect 84 5201 100 5235
rect -100 5154 100 5201
rect -100 2707 100 2754
rect -100 2673 -84 2707
rect 84 2673 100 2707
rect -100 2657 100 2673
rect -100 2599 100 2615
rect -100 2565 -84 2599
rect 84 2565 100 2599
rect -100 2518 100 2565
rect -100 71 100 118
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -118 100 -71
rect -100 -2565 100 -2518
rect -100 -2599 -84 -2565
rect 84 -2599 100 -2565
rect -100 -2615 100 -2599
rect -100 -2673 100 -2657
rect -100 -2707 -84 -2673
rect 84 -2707 100 -2673
rect -100 -2754 100 -2707
rect -100 -5201 100 -5154
rect -100 -5235 -84 -5201
rect 84 -5235 100 -5201
rect -100 -5251 100 -5235
rect -100 -5309 100 -5293
rect -100 -5343 -84 -5309
rect 84 -5343 100 -5309
rect -100 -5390 100 -5343
rect -100 -7837 100 -7790
rect -100 -7871 -84 -7837
rect 84 -7871 100 -7837
rect -100 -7887 100 -7871
rect -100 -7945 100 -7929
rect -100 -7979 -84 -7945
rect 84 -7979 100 -7945
rect -100 -8026 100 -7979
rect -100 -10473 100 -10426
rect -100 -10507 -84 -10473
rect 84 -10507 100 -10473
rect -100 -10523 100 -10507
rect -100 -10581 100 -10565
rect -100 -10615 -84 -10581
rect 84 -10615 100 -10581
rect -100 -10662 100 -10615
rect -100 -13109 100 -13062
rect -100 -13143 -84 -13109
rect 84 -13143 100 -13109
rect -100 -13159 100 -13143
rect -100 -13217 100 -13201
rect -100 -13251 -84 -13217
rect 84 -13251 100 -13217
rect -100 -13298 100 -13251
rect -100 -15745 100 -15698
rect -100 -15779 -84 -15745
rect 84 -15779 100 -15745
rect -100 -15795 100 -15779
rect -100 -15853 100 -15837
rect -100 -15887 -84 -15853
rect 84 -15887 100 -15853
rect -100 -15934 100 -15887
rect -100 -18381 100 -18334
rect -100 -18415 -84 -18381
rect 84 -18415 100 -18381
rect -100 -18431 100 -18415
rect -100 -18489 100 -18473
rect -100 -18523 -84 -18489
rect 84 -18523 100 -18489
rect -100 -18570 100 -18523
rect -100 -21017 100 -20970
rect -100 -21051 -84 -21017
rect 84 -21051 100 -21017
rect -100 -21067 100 -21051
rect -100 -21125 100 -21109
rect -100 -21159 -84 -21125
rect 84 -21159 100 -21125
rect -100 -21206 100 -21159
rect -100 -23653 100 -23606
rect -100 -23687 -84 -23653
rect 84 -23687 100 -23653
rect -100 -23703 100 -23687
rect -100 -23761 100 -23745
rect -100 -23795 -84 -23761
rect 84 -23795 100 -23761
rect -100 -23842 100 -23795
rect -100 -26289 100 -26242
rect -100 -26323 -84 -26289
rect 84 -26323 100 -26289
rect -100 -26339 100 -26323
rect -100 -26397 100 -26381
rect -100 -26431 -84 -26397
rect 84 -26431 100 -26397
rect -100 -26478 100 -26431
rect -100 -28925 100 -28878
rect -100 -28959 -84 -28925
rect 84 -28959 100 -28925
rect -100 -28975 100 -28959
rect -100 -29033 100 -29017
rect -100 -29067 -84 -29033
rect 84 -29067 100 -29033
rect -100 -29114 100 -29067
rect -100 -31561 100 -31514
rect -100 -31595 -84 -31561
rect 84 -31595 100 -31561
rect -100 -31611 100 -31595
rect -100 -31669 100 -31653
rect -100 -31703 -84 -31669
rect 84 -31703 100 -31669
rect -100 -31750 100 -31703
rect -100 -34197 100 -34150
rect -100 -34231 -84 -34197
rect 84 -34231 100 -34197
rect -100 -34247 100 -34231
rect -100 -34305 100 -34289
rect -100 -34339 -84 -34305
rect 84 -34339 100 -34305
rect -100 -34386 100 -34339
rect -100 -36833 100 -36786
rect -100 -36867 -84 -36833
rect 84 -36867 100 -36833
rect -100 -36883 100 -36867
rect -100 -36941 100 -36925
rect -100 -36975 -84 -36941
rect 84 -36975 100 -36941
rect -100 -37022 100 -36975
rect -100 -39469 100 -39422
rect -100 -39503 -84 -39469
rect 84 -39503 100 -39469
rect -100 -39519 100 -39503
rect -100 -39577 100 -39561
rect -100 -39611 -84 -39577
rect 84 -39611 100 -39577
rect -100 -39658 100 -39611
rect -100 -42105 100 -42058
rect -100 -42139 -84 -42105
rect 84 -42139 100 -42105
rect -100 -42155 100 -42139
rect -100 -42213 100 -42197
rect -100 -42247 -84 -42213
rect 84 -42247 100 -42213
rect -100 -42294 100 -42247
rect -100 -44741 100 -44694
rect -100 -44775 -84 -44741
rect 84 -44775 100 -44741
rect -100 -44791 100 -44775
rect -100 -44849 100 -44833
rect -100 -44883 -84 -44849
rect 84 -44883 100 -44849
rect -100 -44930 100 -44883
rect -100 -47377 100 -47330
rect -100 -47411 -84 -47377
rect 84 -47411 100 -47377
rect -100 -47427 100 -47411
rect -100 -47485 100 -47469
rect -100 -47519 -84 -47485
rect 84 -47519 100 -47485
rect -100 -47566 100 -47519
rect -100 -50013 100 -49966
rect -100 -50047 -84 -50013
rect 84 -50047 100 -50013
rect -100 -50063 100 -50047
rect -100 -50121 100 -50105
rect -100 -50155 -84 -50121
rect 84 -50155 100 -50121
rect -100 -50202 100 -50155
rect -100 -52649 100 -52602
rect -100 -52683 -84 -52649
rect 84 -52683 100 -52649
rect -100 -52699 100 -52683
rect -100 -52757 100 -52741
rect -100 -52791 -84 -52757
rect 84 -52791 100 -52757
rect -100 -52838 100 -52791
rect -100 -55285 100 -55238
rect -100 -55319 -84 -55285
rect 84 -55319 100 -55285
rect -100 -55335 100 -55319
rect -100 -55393 100 -55377
rect -100 -55427 -84 -55393
rect 84 -55427 100 -55393
rect -100 -55474 100 -55427
rect -100 -57921 100 -57874
rect -100 -57955 -84 -57921
rect 84 -57955 100 -57921
rect -100 -57971 100 -57955
rect -100 -58029 100 -58013
rect -100 -58063 -84 -58029
rect 84 -58063 100 -58029
rect -100 -58110 100 -58063
rect -100 -60557 100 -60510
rect -100 -60591 -84 -60557
rect 84 -60591 100 -60557
rect -100 -60607 100 -60591
rect -100 -60665 100 -60649
rect -100 -60699 -84 -60665
rect 84 -60699 100 -60665
rect -100 -60746 100 -60699
rect -100 -63193 100 -63146
rect -100 -63227 -84 -63193
rect 84 -63227 100 -63193
rect -100 -63243 100 -63227
rect -100 -63301 100 -63285
rect -100 -63335 -84 -63301
rect 84 -63335 100 -63301
rect -100 -63382 100 -63335
rect -100 -65829 100 -65782
rect -100 -65863 -84 -65829
rect 84 -65863 100 -65829
rect -100 -65879 100 -65863
rect -100 -65937 100 -65921
rect -100 -65971 -84 -65937
rect 84 -65971 100 -65937
rect -100 -66018 100 -65971
rect -100 -68465 100 -68418
rect -100 -68499 -84 -68465
rect 84 -68499 100 -68465
rect -100 -68515 100 -68499
rect -100 -68573 100 -68557
rect -100 -68607 -84 -68573
rect 84 -68607 100 -68573
rect -100 -68654 100 -68607
rect -100 -71101 100 -71054
rect -100 -71135 -84 -71101
rect 84 -71135 100 -71101
rect -100 -71151 100 -71135
rect -100 -71209 100 -71193
rect -100 -71243 -84 -71209
rect 84 -71243 100 -71209
rect -100 -71290 100 -71243
rect -100 -73737 100 -73690
rect -100 -73771 -84 -73737
rect 84 -73771 100 -73737
rect -100 -73787 100 -73771
rect -100 -73845 100 -73829
rect -100 -73879 -84 -73845
rect 84 -73879 100 -73845
rect -100 -73926 100 -73879
rect -100 -76373 100 -76326
rect -100 -76407 -84 -76373
rect 84 -76407 100 -76373
rect -100 -76423 100 -76407
rect -100 -76481 100 -76465
rect -100 -76515 -84 -76481
rect 84 -76515 100 -76481
rect -100 -76562 100 -76515
rect -100 -79009 100 -78962
rect -100 -79043 -84 -79009
rect 84 -79043 100 -79009
rect -100 -79059 100 -79043
rect -100 -79117 100 -79101
rect -100 -79151 -84 -79117
rect 84 -79151 100 -79117
rect -100 -79198 100 -79151
rect -100 -81645 100 -81598
rect -100 -81679 -84 -81645
rect 84 -81679 100 -81645
rect -100 -81695 100 -81679
rect -100 -81753 100 -81737
rect -100 -81787 -84 -81753
rect 84 -81787 100 -81753
rect -100 -81834 100 -81787
rect -100 -84281 100 -84234
rect -100 -84315 -84 -84281
rect 84 -84315 100 -84281
rect -100 -84331 100 -84315
rect -100 -84389 100 -84373
rect -100 -84423 -84 -84389
rect 84 -84423 100 -84389
rect -100 -84470 100 -84423
rect -100 -86917 100 -86870
rect -100 -86951 -84 -86917
rect 84 -86951 100 -86917
rect -100 -86967 100 -86951
rect -100 -87025 100 -87009
rect -100 -87059 -84 -87025
rect 84 -87059 100 -87025
rect -100 -87106 100 -87059
rect -100 -89553 100 -89506
rect -100 -89587 -84 -89553
rect 84 -89587 100 -89553
rect -100 -89603 100 -89587
rect -100 -89661 100 -89645
rect -100 -89695 -84 -89661
rect 84 -89695 100 -89661
rect -100 -89742 100 -89695
rect -100 -92189 100 -92142
rect -100 -92223 -84 -92189
rect 84 -92223 100 -92189
rect -100 -92239 100 -92223
rect -100 -92297 100 -92281
rect -100 -92331 -84 -92297
rect 84 -92331 100 -92297
rect -100 -92378 100 -92331
rect -100 -94825 100 -94778
rect -100 -94859 -84 -94825
rect 84 -94859 100 -94825
rect -100 -94875 100 -94859
rect -100 -94933 100 -94917
rect -100 -94967 -84 -94933
rect 84 -94967 100 -94933
rect -100 -95014 100 -94967
rect -100 -97461 100 -97414
rect -100 -97495 -84 -97461
rect 84 -97495 100 -97461
rect -100 -97511 100 -97495
rect -100 -97569 100 -97553
rect -100 -97603 -84 -97569
rect 84 -97603 100 -97569
rect -100 -97650 100 -97603
rect -100 -100097 100 -100050
rect -100 -100131 -84 -100097
rect 84 -100131 100 -100097
rect -100 -100147 100 -100131
rect -100 -100205 100 -100189
rect -100 -100239 -84 -100205
rect 84 -100239 100 -100205
rect -100 -100286 100 -100239
rect -100 -102733 100 -102686
rect -100 -102767 -84 -102733
rect 84 -102767 100 -102733
rect -100 -102783 100 -102767
rect -100 -102841 100 -102825
rect -100 -102875 -84 -102841
rect 84 -102875 100 -102841
rect -100 -102922 100 -102875
rect -100 -105369 100 -105322
rect -100 -105403 -84 -105369
rect 84 -105403 100 -105369
rect -100 -105419 100 -105403
rect -100 -105477 100 -105461
rect -100 -105511 -84 -105477
rect 84 -105511 100 -105477
rect -100 -105558 100 -105511
rect -100 -108005 100 -107958
rect -100 -108039 -84 -108005
rect 84 -108039 100 -108005
rect -100 -108055 100 -108039
rect -100 -108113 100 -108097
rect -100 -108147 -84 -108113
rect 84 -108147 100 -108113
rect -100 -108194 100 -108147
rect -100 -110641 100 -110594
rect -100 -110675 -84 -110641
rect 84 -110675 100 -110641
rect -100 -110691 100 -110675
rect -100 -110749 100 -110733
rect -100 -110783 -84 -110749
rect 84 -110783 100 -110749
rect -100 -110830 100 -110783
rect -100 -113277 100 -113230
rect -100 -113311 -84 -113277
rect 84 -113311 100 -113277
rect -100 -113327 100 -113311
rect -100 -113385 100 -113369
rect -100 -113419 -84 -113385
rect 84 -113419 100 -113385
rect -100 -113466 100 -113419
rect -100 -115913 100 -115866
rect -100 -115947 -84 -115913
rect 84 -115947 100 -115913
rect -100 -115963 100 -115947
rect -100 -116021 100 -116005
rect -100 -116055 -84 -116021
rect 84 -116055 100 -116021
rect -100 -116102 100 -116055
rect -100 -118549 100 -118502
rect -100 -118583 -84 -118549
rect 84 -118583 100 -118549
rect -100 -118599 100 -118583
rect -100 -118657 100 -118641
rect -100 -118691 -84 -118657
rect 84 -118691 100 -118657
rect -100 -118738 100 -118691
rect -100 -121185 100 -121138
rect -100 -121219 -84 -121185
rect 84 -121219 100 -121185
rect -100 -121235 100 -121219
rect -100 -121293 100 -121277
rect -100 -121327 -84 -121293
rect 84 -121327 100 -121293
rect -100 -121374 100 -121327
rect -100 -123821 100 -123774
rect -100 -123855 -84 -123821
rect 84 -123855 100 -123821
rect -100 -123871 100 -123855
rect -100 -123929 100 -123913
rect -100 -123963 -84 -123929
rect 84 -123963 100 -123929
rect -100 -124010 100 -123963
rect -100 -126457 100 -126410
rect -100 -126491 -84 -126457
rect 84 -126491 100 -126457
rect -100 -126507 100 -126491
rect -100 -126565 100 -126549
rect -100 -126599 -84 -126565
rect 84 -126599 100 -126565
rect -100 -126646 100 -126599
rect -100 -129093 100 -129046
rect -100 -129127 -84 -129093
rect 84 -129127 100 -129093
rect -100 -129143 100 -129127
rect -100 -129201 100 -129185
rect -100 -129235 -84 -129201
rect 84 -129235 100 -129201
rect -100 -129282 100 -129235
rect -100 -131729 100 -131682
rect -100 -131763 -84 -131729
rect 84 -131763 100 -131729
rect -100 -131779 100 -131763
rect -100 -131837 100 -131821
rect -100 -131871 -84 -131837
rect 84 -131871 100 -131837
rect -100 -131918 100 -131871
rect -100 -134365 100 -134318
rect -100 -134399 -84 -134365
rect 84 -134399 100 -134365
rect -100 -134415 100 -134399
rect -100 -134473 100 -134457
rect -100 -134507 -84 -134473
rect 84 -134507 100 -134473
rect -100 -134554 100 -134507
rect -100 -137001 100 -136954
rect -100 -137035 -84 -137001
rect 84 -137035 100 -137001
rect -100 -137051 100 -137035
rect -100 -137109 100 -137093
rect -100 -137143 -84 -137109
rect 84 -137143 100 -137109
rect -100 -137190 100 -137143
rect -100 -139637 100 -139590
rect -100 -139671 -84 -139637
rect 84 -139671 100 -139637
rect -100 -139687 100 -139671
rect -100 -139745 100 -139729
rect -100 -139779 -84 -139745
rect 84 -139779 100 -139745
rect -100 -139826 100 -139779
rect -100 -142273 100 -142226
rect -100 -142307 -84 -142273
rect 84 -142307 100 -142273
rect -100 -142323 100 -142307
rect -100 -142381 100 -142365
rect -100 -142415 -84 -142381
rect 84 -142415 100 -142381
rect -100 -142462 100 -142415
rect -100 -144909 100 -144862
rect -100 -144943 -84 -144909
rect 84 -144943 100 -144909
rect -100 -144959 100 -144943
rect -100 -145017 100 -145001
rect -100 -145051 -84 -145017
rect 84 -145051 100 -145017
rect -100 -145098 100 -145051
rect -100 -147545 100 -147498
rect -100 -147579 -84 -147545
rect 84 -147579 100 -147545
rect -100 -147595 100 -147579
rect -100 -147653 100 -147637
rect -100 -147687 -84 -147653
rect 84 -147687 100 -147653
rect -100 -147734 100 -147687
rect -100 -150181 100 -150134
rect -100 -150215 -84 -150181
rect 84 -150215 100 -150181
rect -100 -150231 100 -150215
rect -100 -150289 100 -150273
rect -100 -150323 -84 -150289
rect 84 -150323 100 -150289
rect -100 -150370 100 -150323
rect -100 -152817 100 -152770
rect -100 -152851 -84 -152817
rect 84 -152851 100 -152817
rect -100 -152867 100 -152851
rect -100 -152925 100 -152909
rect -100 -152959 -84 -152925
rect 84 -152959 100 -152925
rect -100 -153006 100 -152959
rect -100 -155453 100 -155406
rect -100 -155487 -84 -155453
rect 84 -155487 100 -155453
rect -100 -155503 100 -155487
rect -100 -155561 100 -155545
rect -100 -155595 -84 -155561
rect 84 -155595 100 -155561
rect -100 -155642 100 -155595
rect -100 -158089 100 -158042
rect -100 -158123 -84 -158089
rect 84 -158123 100 -158089
rect -100 -158139 100 -158123
rect -100 -158197 100 -158181
rect -100 -158231 -84 -158197
rect 84 -158231 100 -158197
rect -100 -158278 100 -158231
rect -100 -160725 100 -160678
rect -100 -160759 -84 -160725
rect 84 -160759 100 -160725
rect -100 -160775 100 -160759
rect -100 -160833 100 -160817
rect -100 -160867 -84 -160833
rect 84 -160867 100 -160833
rect -100 -160914 100 -160867
rect -100 -163361 100 -163314
rect -100 -163395 -84 -163361
rect 84 -163395 100 -163361
rect -100 -163411 100 -163395
rect -100 -163469 100 -163453
rect -100 -163503 -84 -163469
rect 84 -163503 100 -163469
rect -100 -163550 100 -163503
rect -100 -165997 100 -165950
rect -100 -166031 -84 -165997
rect 84 -166031 100 -165997
rect -100 -166047 100 -166031
rect -100 -166105 100 -166089
rect -100 -166139 -84 -166105
rect 84 -166139 100 -166105
rect -100 -166186 100 -166139
rect -100 -168633 100 -168586
rect -100 -168667 -84 -168633
rect 84 -168667 100 -168633
rect -100 -168683 100 -168667
rect -100 -168741 100 -168725
rect -100 -168775 -84 -168741
rect 84 -168775 100 -168741
rect -100 -168822 100 -168775
rect -100 -171269 100 -171222
rect -100 -171303 -84 -171269
rect 84 -171303 100 -171269
rect -100 -171319 100 -171303
rect -100 -171377 100 -171361
rect -100 -171411 -84 -171377
rect 84 -171411 100 -171377
rect -100 -171458 100 -171411
rect -100 -173905 100 -173858
rect -100 -173939 -84 -173905
rect 84 -173939 100 -173905
rect -100 -173955 100 -173939
rect -100 -174013 100 -173997
rect -100 -174047 -84 -174013
rect 84 -174047 100 -174013
rect -100 -174094 100 -174047
rect -100 -176541 100 -176494
rect -100 -176575 -84 -176541
rect 84 -176575 100 -176541
rect -100 -176591 100 -176575
rect -100 -176649 100 -176633
rect -100 -176683 -84 -176649
rect 84 -176683 100 -176649
rect -100 -176730 100 -176683
rect -100 -179177 100 -179130
rect -100 -179211 -84 -179177
rect 84 -179211 100 -179177
rect -100 -179227 100 -179211
rect -100 -179285 100 -179269
rect -100 -179319 -84 -179285
rect 84 -179319 100 -179285
rect -100 -179366 100 -179319
rect -100 -181813 100 -181766
rect -100 -181847 -84 -181813
rect 84 -181847 100 -181813
rect -100 -181863 100 -181847
rect -100 -181921 100 -181905
rect -100 -181955 -84 -181921
rect 84 -181955 100 -181921
rect -100 -182002 100 -181955
rect -100 -184449 100 -184402
rect -100 -184483 -84 -184449
rect 84 -184483 100 -184449
rect -100 -184499 100 -184483
rect -100 -184557 100 -184541
rect -100 -184591 -84 -184557
rect 84 -184591 100 -184557
rect -100 -184638 100 -184591
rect -100 -187085 100 -187038
rect -100 -187119 -84 -187085
rect 84 -187119 100 -187085
rect -100 -187135 100 -187119
rect -100 -187193 100 -187177
rect -100 -187227 -84 -187193
rect 84 -187227 100 -187193
rect -100 -187274 100 -187227
rect -100 -189721 100 -189674
rect -100 -189755 -84 -189721
rect 84 -189755 100 -189721
rect -100 -189771 100 -189755
rect -100 -189829 100 -189813
rect -100 -189863 -84 -189829
rect 84 -189863 100 -189829
rect -100 -189910 100 -189863
rect -100 -192357 100 -192310
rect -100 -192391 -84 -192357
rect 84 -192391 100 -192357
rect -100 -192407 100 -192391
rect -100 -192465 100 -192449
rect -100 -192499 -84 -192465
rect 84 -192499 100 -192465
rect -100 -192546 100 -192499
rect -100 -194993 100 -194946
rect -100 -195027 -84 -194993
rect 84 -195027 100 -194993
rect -100 -195043 100 -195027
rect -100 -195101 100 -195085
rect -100 -195135 -84 -195101
rect 84 -195135 100 -195101
rect -100 -195182 100 -195135
rect -100 -197629 100 -197582
rect -100 -197663 -84 -197629
rect 84 -197663 100 -197629
rect -100 -197679 100 -197663
rect -100 -197737 100 -197721
rect -100 -197771 -84 -197737
rect 84 -197771 100 -197737
rect -100 -197818 100 -197771
rect -100 -200265 100 -200218
rect -100 -200299 -84 -200265
rect 84 -200299 100 -200265
rect -100 -200315 100 -200299
rect -100 -200373 100 -200357
rect -100 -200407 -84 -200373
rect 84 -200407 100 -200373
rect -100 -200454 100 -200407
rect -100 -202901 100 -202854
rect -100 -202935 -84 -202901
rect 84 -202935 100 -202901
rect -100 -202951 100 -202935
rect -100 -203009 100 -202993
rect -100 -203043 -84 -203009
rect 84 -203043 100 -203009
rect -100 -203090 100 -203043
rect -100 -205537 100 -205490
rect -100 -205571 -84 -205537
rect 84 -205571 100 -205537
rect -100 -205587 100 -205571
rect -100 -205645 100 -205629
rect -100 -205679 -84 -205645
rect 84 -205679 100 -205645
rect -100 -205726 100 -205679
rect -100 -208173 100 -208126
rect -100 -208207 -84 -208173
rect 84 -208207 100 -208173
rect -100 -208223 100 -208207
rect -100 -208281 100 -208265
rect -100 -208315 -84 -208281
rect 84 -208315 100 -208281
rect -100 -208362 100 -208315
rect -100 -210809 100 -210762
rect -100 -210843 -84 -210809
rect 84 -210843 100 -210809
rect -100 -210859 100 -210843
rect -100 -210917 100 -210901
rect -100 -210951 -84 -210917
rect 84 -210951 100 -210917
rect -100 -210998 100 -210951
rect -100 -213445 100 -213398
rect -100 -213479 -84 -213445
rect 84 -213479 100 -213445
rect -100 -213495 100 -213479
rect -100 -213553 100 -213537
rect -100 -213587 -84 -213553
rect 84 -213587 100 -213553
rect -100 -213634 100 -213587
rect -100 -216081 100 -216034
rect -100 -216115 -84 -216081
rect 84 -216115 100 -216081
rect -100 -216131 100 -216115
rect -100 -216189 100 -216173
rect -100 -216223 -84 -216189
rect 84 -216223 100 -216189
rect -100 -216270 100 -216223
rect -100 -218717 100 -218670
rect -100 -218751 -84 -218717
rect 84 -218751 100 -218717
rect -100 -218767 100 -218751
rect -100 -218825 100 -218809
rect -100 -218859 -84 -218825
rect 84 -218859 100 -218825
rect -100 -218906 100 -218859
rect -100 -221353 100 -221306
rect -100 -221387 -84 -221353
rect 84 -221387 100 -221353
rect -100 -221403 100 -221387
rect -100 -221461 100 -221445
rect -100 -221495 -84 -221461
rect 84 -221495 100 -221461
rect -100 -221542 100 -221495
rect -100 -223989 100 -223942
rect -100 -224023 -84 -223989
rect 84 -224023 100 -223989
rect -100 -224039 100 -224023
rect -100 -224097 100 -224081
rect -100 -224131 -84 -224097
rect 84 -224131 100 -224097
rect -100 -224178 100 -224131
rect -100 -226625 100 -226578
rect -100 -226659 -84 -226625
rect 84 -226659 100 -226625
rect -100 -226675 100 -226659
rect -100 -226733 100 -226717
rect -100 -226767 -84 -226733
rect 84 -226767 100 -226733
rect -100 -226814 100 -226767
rect -100 -229261 100 -229214
rect -100 -229295 -84 -229261
rect 84 -229295 100 -229261
rect -100 -229311 100 -229295
rect -100 -229369 100 -229353
rect -100 -229403 -84 -229369
rect 84 -229403 100 -229369
rect -100 -229450 100 -229403
rect -100 -231897 100 -231850
rect -100 -231931 -84 -231897
rect 84 -231931 100 -231897
rect -100 -231947 100 -231931
rect -100 -232005 100 -231989
rect -100 -232039 -84 -232005
rect 84 -232039 100 -232005
rect -100 -232086 100 -232039
rect -100 -234533 100 -234486
rect -100 -234567 -84 -234533
rect 84 -234567 100 -234533
rect -100 -234583 100 -234567
rect -100 -234641 100 -234625
rect -100 -234675 -84 -234641
rect 84 -234675 100 -234641
rect -100 -234722 100 -234675
rect -100 -237169 100 -237122
rect -100 -237203 -84 -237169
rect 84 -237203 100 -237169
rect -100 -237219 100 -237203
rect -100 -237277 100 -237261
rect -100 -237311 -84 -237277
rect 84 -237311 100 -237277
rect -100 -237358 100 -237311
rect -100 -239805 100 -239758
rect -100 -239839 -84 -239805
rect 84 -239839 100 -239805
rect -100 -239855 100 -239839
rect -100 -239913 100 -239897
rect -100 -239947 -84 -239913
rect 84 -239947 100 -239913
rect -100 -239994 100 -239947
rect -100 -242441 100 -242394
rect -100 -242475 -84 -242441
rect 84 -242475 100 -242441
rect -100 -242491 100 -242475
rect -100 -242549 100 -242533
rect -100 -242583 -84 -242549
rect 84 -242583 100 -242549
rect -100 -242630 100 -242583
rect -100 -245077 100 -245030
rect -100 -245111 -84 -245077
rect 84 -245111 100 -245077
rect -100 -245127 100 -245111
rect -100 -245185 100 -245169
rect -100 -245219 -84 -245185
rect 84 -245219 100 -245185
rect -100 -245266 100 -245219
rect -100 -247713 100 -247666
rect -100 -247747 -84 -247713
rect 84 -247747 100 -247713
rect -100 -247763 100 -247747
rect -100 -247821 100 -247805
rect -100 -247855 -84 -247821
rect 84 -247855 100 -247821
rect -100 -247902 100 -247855
rect -100 -250349 100 -250302
rect -100 -250383 -84 -250349
rect 84 -250383 100 -250349
rect -100 -250399 100 -250383
rect -100 -250457 100 -250441
rect -100 -250491 -84 -250457
rect 84 -250491 100 -250457
rect -100 -250538 100 -250491
rect -100 -252985 100 -252938
rect -100 -253019 -84 -252985
rect 84 -253019 100 -252985
rect -100 -253035 100 -253019
rect -100 -253093 100 -253077
rect -100 -253127 -84 -253093
rect 84 -253127 100 -253093
rect -100 -253174 100 -253127
rect -100 -255621 100 -255574
rect -100 -255655 -84 -255621
rect 84 -255655 100 -255621
rect -100 -255671 100 -255655
rect -100 -255729 100 -255713
rect -100 -255763 -84 -255729
rect 84 -255763 100 -255729
rect -100 -255810 100 -255763
rect -100 -258257 100 -258210
rect -100 -258291 -84 -258257
rect 84 -258291 100 -258257
rect -100 -258307 100 -258291
rect -100 -258365 100 -258349
rect -100 -258399 -84 -258365
rect 84 -258399 100 -258365
rect -100 -258446 100 -258399
rect -100 -260893 100 -260846
rect -100 -260927 -84 -260893
rect 84 -260927 100 -260893
rect -100 -260943 100 -260927
rect -100 -261001 100 -260985
rect -100 -261035 -84 -261001
rect 84 -261035 100 -261001
rect -100 -261082 100 -261035
rect -100 -263529 100 -263482
rect -100 -263563 -84 -263529
rect 84 -263563 100 -263529
rect -100 -263579 100 -263563
rect -100 -263637 100 -263621
rect -100 -263671 -84 -263637
rect 84 -263671 100 -263637
rect -100 -263718 100 -263671
rect -100 -266165 100 -266118
rect -100 -266199 -84 -266165
rect 84 -266199 100 -266165
rect -100 -266215 100 -266199
rect -100 -266273 100 -266257
rect -100 -266307 -84 -266273
rect 84 -266307 100 -266273
rect -100 -266354 100 -266307
rect -100 -268801 100 -268754
rect -100 -268835 -84 -268801
rect 84 -268835 100 -268801
rect -100 -268851 100 -268835
rect -100 -268909 100 -268893
rect -100 -268943 -84 -268909
rect 84 -268943 100 -268909
rect -100 -268990 100 -268943
rect -100 -271437 100 -271390
rect -100 -271471 -84 -271437
rect 84 -271471 100 -271437
rect -100 -271487 100 -271471
rect -100 -271545 100 -271529
rect -100 -271579 -84 -271545
rect 84 -271579 100 -271545
rect -100 -271626 100 -271579
rect -100 -274073 100 -274026
rect -100 -274107 -84 -274073
rect 84 -274107 100 -274073
rect -100 -274123 100 -274107
rect -100 -274181 100 -274165
rect -100 -274215 -84 -274181
rect 84 -274215 100 -274181
rect -100 -274262 100 -274215
rect -100 -276709 100 -276662
rect -100 -276743 -84 -276709
rect 84 -276743 100 -276709
rect -100 -276759 100 -276743
rect -100 -276817 100 -276801
rect -100 -276851 -84 -276817
rect 84 -276851 100 -276817
rect -100 -276898 100 -276851
rect -100 -279345 100 -279298
rect -100 -279379 -84 -279345
rect 84 -279379 100 -279345
rect -100 -279395 100 -279379
rect -100 -279453 100 -279437
rect -100 -279487 -84 -279453
rect 84 -279487 100 -279453
rect -100 -279534 100 -279487
rect -100 -281981 100 -281934
rect -100 -282015 -84 -281981
rect 84 -282015 100 -281981
rect -100 -282031 100 -282015
rect -100 -282089 100 -282073
rect -100 -282123 -84 -282089
rect 84 -282123 100 -282089
rect -100 -282170 100 -282123
rect -100 -284617 100 -284570
rect -100 -284651 -84 -284617
rect 84 -284651 100 -284617
rect -100 -284667 100 -284651
rect -100 -284725 100 -284709
rect -100 -284759 -84 -284725
rect 84 -284759 100 -284725
rect -100 -284806 100 -284759
rect -100 -287253 100 -287206
rect -100 -287287 -84 -287253
rect 84 -287287 100 -287253
rect -100 -287303 100 -287287
rect -100 -287361 100 -287345
rect -100 -287395 -84 -287361
rect 84 -287395 100 -287361
rect -100 -287442 100 -287395
rect -100 -289889 100 -289842
rect -100 -289923 -84 -289889
rect 84 -289923 100 -289889
rect -100 -289939 100 -289923
rect -100 -289997 100 -289981
rect -100 -290031 -84 -289997
rect 84 -290031 100 -289997
rect -100 -290078 100 -290031
rect -100 -292525 100 -292478
rect -100 -292559 -84 -292525
rect 84 -292559 100 -292525
rect -100 -292575 100 -292559
rect -100 -292633 100 -292617
rect -100 -292667 -84 -292633
rect 84 -292667 100 -292633
rect -100 -292714 100 -292667
rect -100 -295161 100 -295114
rect -100 -295195 -84 -295161
rect 84 -295195 100 -295161
rect -100 -295211 100 -295195
rect -100 -295269 100 -295253
rect -100 -295303 -84 -295269
rect 84 -295303 100 -295269
rect -100 -295350 100 -295303
rect -100 -297797 100 -297750
rect -100 -297831 -84 -297797
rect 84 -297831 100 -297797
rect -100 -297847 100 -297831
rect -100 -297905 100 -297889
rect -100 -297939 -84 -297905
rect 84 -297939 100 -297905
rect -100 -297986 100 -297939
rect -100 -300433 100 -300386
rect -100 -300467 -84 -300433
rect 84 -300467 100 -300433
rect -100 -300483 100 -300467
rect -100 -300541 100 -300525
rect -100 -300575 -84 -300541
rect 84 -300575 100 -300541
rect -100 -300622 100 -300575
rect -100 -303069 100 -303022
rect -100 -303103 -84 -303069
rect 84 -303103 100 -303069
rect -100 -303119 100 -303103
rect -100 -303177 100 -303161
rect -100 -303211 -84 -303177
rect 84 -303211 100 -303177
rect -100 -303258 100 -303211
rect -100 -305705 100 -305658
rect -100 -305739 -84 -305705
rect 84 -305739 100 -305705
rect -100 -305755 100 -305739
rect -100 -305813 100 -305797
rect -100 -305847 -84 -305813
rect 84 -305847 100 -305813
rect -100 -305894 100 -305847
rect -100 -308341 100 -308294
rect -100 -308375 -84 -308341
rect 84 -308375 100 -308341
rect -100 -308391 100 -308375
rect -100 -308449 100 -308433
rect -100 -308483 -84 -308449
rect 84 -308483 100 -308449
rect -100 -308530 100 -308483
rect -100 -310977 100 -310930
rect -100 -311011 -84 -310977
rect 84 -311011 100 -310977
rect -100 -311027 100 -311011
rect -100 -311085 100 -311069
rect -100 -311119 -84 -311085
rect 84 -311119 100 -311085
rect -100 -311166 100 -311119
rect -100 -313613 100 -313566
rect -100 -313647 -84 -313613
rect 84 -313647 100 -313613
rect -100 -313663 100 -313647
rect -100 -313721 100 -313705
rect -100 -313755 -84 -313721
rect 84 -313755 100 -313721
rect -100 -313802 100 -313755
rect -100 -316249 100 -316202
rect -100 -316283 -84 -316249
rect 84 -316283 100 -316249
rect -100 -316299 100 -316283
rect -100 -316357 100 -316341
rect -100 -316391 -84 -316357
rect 84 -316391 100 -316357
rect -100 -316438 100 -316391
rect -100 -318885 100 -318838
rect -100 -318919 -84 -318885
rect 84 -318919 100 -318885
rect -100 -318935 100 -318919
rect -100 -318993 100 -318977
rect -100 -319027 -84 -318993
rect 84 -319027 100 -318993
rect -100 -319074 100 -319027
rect -100 -321521 100 -321474
rect -100 -321555 -84 -321521
rect 84 -321555 100 -321521
rect -100 -321571 100 -321555
rect -100 -321629 100 -321613
rect -100 -321663 -84 -321629
rect 84 -321663 100 -321629
rect -100 -321710 100 -321663
rect -100 -324157 100 -324110
rect -100 -324191 -84 -324157
rect 84 -324191 100 -324157
rect -100 -324207 100 -324191
rect -100 -324265 100 -324249
rect -100 -324299 -84 -324265
rect 84 -324299 100 -324265
rect -100 -324346 100 -324299
rect -100 -326793 100 -326746
rect -100 -326827 -84 -326793
rect 84 -326827 100 -326793
rect -100 -326843 100 -326827
rect -100 -326901 100 -326885
rect -100 -326935 -84 -326901
rect 84 -326935 100 -326901
rect -100 -326982 100 -326935
rect -100 -329429 100 -329382
rect -100 -329463 -84 -329429
rect 84 -329463 100 -329429
rect -100 -329479 100 -329463
rect -100 -329537 100 -329521
rect -100 -329571 -84 -329537
rect 84 -329571 100 -329537
rect -100 -329618 100 -329571
rect -100 -332065 100 -332018
rect -100 -332099 -84 -332065
rect 84 -332099 100 -332065
rect -100 -332115 100 -332099
rect -100 -332173 100 -332157
rect -100 -332207 -84 -332173
rect 84 -332207 100 -332173
rect -100 -332254 100 -332207
rect -100 -334701 100 -334654
rect -100 -334735 -84 -334701
rect 84 -334735 100 -334701
rect -100 -334751 100 -334735
rect -100 -334809 100 -334793
rect -100 -334843 -84 -334809
rect 84 -334843 100 -334809
rect -100 -334890 100 -334843
rect -100 -337337 100 -337290
rect -100 -337371 -84 -337337
rect 84 -337371 100 -337337
rect -100 -337387 100 -337371
<< polycont >>
rect -84 337337 84 337371
rect -84 334809 84 334843
rect -84 334701 84 334735
rect -84 332173 84 332207
rect -84 332065 84 332099
rect -84 329537 84 329571
rect -84 329429 84 329463
rect -84 326901 84 326935
rect -84 326793 84 326827
rect -84 324265 84 324299
rect -84 324157 84 324191
rect -84 321629 84 321663
rect -84 321521 84 321555
rect -84 318993 84 319027
rect -84 318885 84 318919
rect -84 316357 84 316391
rect -84 316249 84 316283
rect -84 313721 84 313755
rect -84 313613 84 313647
rect -84 311085 84 311119
rect -84 310977 84 311011
rect -84 308449 84 308483
rect -84 308341 84 308375
rect -84 305813 84 305847
rect -84 305705 84 305739
rect -84 303177 84 303211
rect -84 303069 84 303103
rect -84 300541 84 300575
rect -84 300433 84 300467
rect -84 297905 84 297939
rect -84 297797 84 297831
rect -84 295269 84 295303
rect -84 295161 84 295195
rect -84 292633 84 292667
rect -84 292525 84 292559
rect -84 289997 84 290031
rect -84 289889 84 289923
rect -84 287361 84 287395
rect -84 287253 84 287287
rect -84 284725 84 284759
rect -84 284617 84 284651
rect -84 282089 84 282123
rect -84 281981 84 282015
rect -84 279453 84 279487
rect -84 279345 84 279379
rect -84 276817 84 276851
rect -84 276709 84 276743
rect -84 274181 84 274215
rect -84 274073 84 274107
rect -84 271545 84 271579
rect -84 271437 84 271471
rect -84 268909 84 268943
rect -84 268801 84 268835
rect -84 266273 84 266307
rect -84 266165 84 266199
rect -84 263637 84 263671
rect -84 263529 84 263563
rect -84 261001 84 261035
rect -84 260893 84 260927
rect -84 258365 84 258399
rect -84 258257 84 258291
rect -84 255729 84 255763
rect -84 255621 84 255655
rect -84 253093 84 253127
rect -84 252985 84 253019
rect -84 250457 84 250491
rect -84 250349 84 250383
rect -84 247821 84 247855
rect -84 247713 84 247747
rect -84 245185 84 245219
rect -84 245077 84 245111
rect -84 242549 84 242583
rect -84 242441 84 242475
rect -84 239913 84 239947
rect -84 239805 84 239839
rect -84 237277 84 237311
rect -84 237169 84 237203
rect -84 234641 84 234675
rect -84 234533 84 234567
rect -84 232005 84 232039
rect -84 231897 84 231931
rect -84 229369 84 229403
rect -84 229261 84 229295
rect -84 226733 84 226767
rect -84 226625 84 226659
rect -84 224097 84 224131
rect -84 223989 84 224023
rect -84 221461 84 221495
rect -84 221353 84 221387
rect -84 218825 84 218859
rect -84 218717 84 218751
rect -84 216189 84 216223
rect -84 216081 84 216115
rect -84 213553 84 213587
rect -84 213445 84 213479
rect -84 210917 84 210951
rect -84 210809 84 210843
rect -84 208281 84 208315
rect -84 208173 84 208207
rect -84 205645 84 205679
rect -84 205537 84 205571
rect -84 203009 84 203043
rect -84 202901 84 202935
rect -84 200373 84 200407
rect -84 200265 84 200299
rect -84 197737 84 197771
rect -84 197629 84 197663
rect -84 195101 84 195135
rect -84 194993 84 195027
rect -84 192465 84 192499
rect -84 192357 84 192391
rect -84 189829 84 189863
rect -84 189721 84 189755
rect -84 187193 84 187227
rect -84 187085 84 187119
rect -84 184557 84 184591
rect -84 184449 84 184483
rect -84 181921 84 181955
rect -84 181813 84 181847
rect -84 179285 84 179319
rect -84 179177 84 179211
rect -84 176649 84 176683
rect -84 176541 84 176575
rect -84 174013 84 174047
rect -84 173905 84 173939
rect -84 171377 84 171411
rect -84 171269 84 171303
rect -84 168741 84 168775
rect -84 168633 84 168667
rect -84 166105 84 166139
rect -84 165997 84 166031
rect -84 163469 84 163503
rect -84 163361 84 163395
rect -84 160833 84 160867
rect -84 160725 84 160759
rect -84 158197 84 158231
rect -84 158089 84 158123
rect -84 155561 84 155595
rect -84 155453 84 155487
rect -84 152925 84 152959
rect -84 152817 84 152851
rect -84 150289 84 150323
rect -84 150181 84 150215
rect -84 147653 84 147687
rect -84 147545 84 147579
rect -84 145017 84 145051
rect -84 144909 84 144943
rect -84 142381 84 142415
rect -84 142273 84 142307
rect -84 139745 84 139779
rect -84 139637 84 139671
rect -84 137109 84 137143
rect -84 137001 84 137035
rect -84 134473 84 134507
rect -84 134365 84 134399
rect -84 131837 84 131871
rect -84 131729 84 131763
rect -84 129201 84 129235
rect -84 129093 84 129127
rect -84 126565 84 126599
rect -84 126457 84 126491
rect -84 123929 84 123963
rect -84 123821 84 123855
rect -84 121293 84 121327
rect -84 121185 84 121219
rect -84 118657 84 118691
rect -84 118549 84 118583
rect -84 116021 84 116055
rect -84 115913 84 115947
rect -84 113385 84 113419
rect -84 113277 84 113311
rect -84 110749 84 110783
rect -84 110641 84 110675
rect -84 108113 84 108147
rect -84 108005 84 108039
rect -84 105477 84 105511
rect -84 105369 84 105403
rect -84 102841 84 102875
rect -84 102733 84 102767
rect -84 100205 84 100239
rect -84 100097 84 100131
rect -84 97569 84 97603
rect -84 97461 84 97495
rect -84 94933 84 94967
rect -84 94825 84 94859
rect -84 92297 84 92331
rect -84 92189 84 92223
rect -84 89661 84 89695
rect -84 89553 84 89587
rect -84 87025 84 87059
rect -84 86917 84 86951
rect -84 84389 84 84423
rect -84 84281 84 84315
rect -84 81753 84 81787
rect -84 81645 84 81679
rect -84 79117 84 79151
rect -84 79009 84 79043
rect -84 76481 84 76515
rect -84 76373 84 76407
rect -84 73845 84 73879
rect -84 73737 84 73771
rect -84 71209 84 71243
rect -84 71101 84 71135
rect -84 68573 84 68607
rect -84 68465 84 68499
rect -84 65937 84 65971
rect -84 65829 84 65863
rect -84 63301 84 63335
rect -84 63193 84 63227
rect -84 60665 84 60699
rect -84 60557 84 60591
rect -84 58029 84 58063
rect -84 57921 84 57955
rect -84 55393 84 55427
rect -84 55285 84 55319
rect -84 52757 84 52791
rect -84 52649 84 52683
rect -84 50121 84 50155
rect -84 50013 84 50047
rect -84 47485 84 47519
rect -84 47377 84 47411
rect -84 44849 84 44883
rect -84 44741 84 44775
rect -84 42213 84 42247
rect -84 42105 84 42139
rect -84 39577 84 39611
rect -84 39469 84 39503
rect -84 36941 84 36975
rect -84 36833 84 36867
rect -84 34305 84 34339
rect -84 34197 84 34231
rect -84 31669 84 31703
rect -84 31561 84 31595
rect -84 29033 84 29067
rect -84 28925 84 28959
rect -84 26397 84 26431
rect -84 26289 84 26323
rect -84 23761 84 23795
rect -84 23653 84 23687
rect -84 21125 84 21159
rect -84 21017 84 21051
rect -84 18489 84 18523
rect -84 18381 84 18415
rect -84 15853 84 15887
rect -84 15745 84 15779
rect -84 13217 84 13251
rect -84 13109 84 13143
rect -84 10581 84 10615
rect -84 10473 84 10507
rect -84 7945 84 7979
rect -84 7837 84 7871
rect -84 5309 84 5343
rect -84 5201 84 5235
rect -84 2673 84 2707
rect -84 2565 84 2599
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -2599 84 -2565
rect -84 -2707 84 -2673
rect -84 -5235 84 -5201
rect -84 -5343 84 -5309
rect -84 -7871 84 -7837
rect -84 -7979 84 -7945
rect -84 -10507 84 -10473
rect -84 -10615 84 -10581
rect -84 -13143 84 -13109
rect -84 -13251 84 -13217
rect -84 -15779 84 -15745
rect -84 -15887 84 -15853
rect -84 -18415 84 -18381
rect -84 -18523 84 -18489
rect -84 -21051 84 -21017
rect -84 -21159 84 -21125
rect -84 -23687 84 -23653
rect -84 -23795 84 -23761
rect -84 -26323 84 -26289
rect -84 -26431 84 -26397
rect -84 -28959 84 -28925
rect -84 -29067 84 -29033
rect -84 -31595 84 -31561
rect -84 -31703 84 -31669
rect -84 -34231 84 -34197
rect -84 -34339 84 -34305
rect -84 -36867 84 -36833
rect -84 -36975 84 -36941
rect -84 -39503 84 -39469
rect -84 -39611 84 -39577
rect -84 -42139 84 -42105
rect -84 -42247 84 -42213
rect -84 -44775 84 -44741
rect -84 -44883 84 -44849
rect -84 -47411 84 -47377
rect -84 -47519 84 -47485
rect -84 -50047 84 -50013
rect -84 -50155 84 -50121
rect -84 -52683 84 -52649
rect -84 -52791 84 -52757
rect -84 -55319 84 -55285
rect -84 -55427 84 -55393
rect -84 -57955 84 -57921
rect -84 -58063 84 -58029
rect -84 -60591 84 -60557
rect -84 -60699 84 -60665
rect -84 -63227 84 -63193
rect -84 -63335 84 -63301
rect -84 -65863 84 -65829
rect -84 -65971 84 -65937
rect -84 -68499 84 -68465
rect -84 -68607 84 -68573
rect -84 -71135 84 -71101
rect -84 -71243 84 -71209
rect -84 -73771 84 -73737
rect -84 -73879 84 -73845
rect -84 -76407 84 -76373
rect -84 -76515 84 -76481
rect -84 -79043 84 -79009
rect -84 -79151 84 -79117
rect -84 -81679 84 -81645
rect -84 -81787 84 -81753
rect -84 -84315 84 -84281
rect -84 -84423 84 -84389
rect -84 -86951 84 -86917
rect -84 -87059 84 -87025
rect -84 -89587 84 -89553
rect -84 -89695 84 -89661
rect -84 -92223 84 -92189
rect -84 -92331 84 -92297
rect -84 -94859 84 -94825
rect -84 -94967 84 -94933
rect -84 -97495 84 -97461
rect -84 -97603 84 -97569
rect -84 -100131 84 -100097
rect -84 -100239 84 -100205
rect -84 -102767 84 -102733
rect -84 -102875 84 -102841
rect -84 -105403 84 -105369
rect -84 -105511 84 -105477
rect -84 -108039 84 -108005
rect -84 -108147 84 -108113
rect -84 -110675 84 -110641
rect -84 -110783 84 -110749
rect -84 -113311 84 -113277
rect -84 -113419 84 -113385
rect -84 -115947 84 -115913
rect -84 -116055 84 -116021
rect -84 -118583 84 -118549
rect -84 -118691 84 -118657
rect -84 -121219 84 -121185
rect -84 -121327 84 -121293
rect -84 -123855 84 -123821
rect -84 -123963 84 -123929
rect -84 -126491 84 -126457
rect -84 -126599 84 -126565
rect -84 -129127 84 -129093
rect -84 -129235 84 -129201
rect -84 -131763 84 -131729
rect -84 -131871 84 -131837
rect -84 -134399 84 -134365
rect -84 -134507 84 -134473
rect -84 -137035 84 -137001
rect -84 -137143 84 -137109
rect -84 -139671 84 -139637
rect -84 -139779 84 -139745
rect -84 -142307 84 -142273
rect -84 -142415 84 -142381
rect -84 -144943 84 -144909
rect -84 -145051 84 -145017
rect -84 -147579 84 -147545
rect -84 -147687 84 -147653
rect -84 -150215 84 -150181
rect -84 -150323 84 -150289
rect -84 -152851 84 -152817
rect -84 -152959 84 -152925
rect -84 -155487 84 -155453
rect -84 -155595 84 -155561
rect -84 -158123 84 -158089
rect -84 -158231 84 -158197
rect -84 -160759 84 -160725
rect -84 -160867 84 -160833
rect -84 -163395 84 -163361
rect -84 -163503 84 -163469
rect -84 -166031 84 -165997
rect -84 -166139 84 -166105
rect -84 -168667 84 -168633
rect -84 -168775 84 -168741
rect -84 -171303 84 -171269
rect -84 -171411 84 -171377
rect -84 -173939 84 -173905
rect -84 -174047 84 -174013
rect -84 -176575 84 -176541
rect -84 -176683 84 -176649
rect -84 -179211 84 -179177
rect -84 -179319 84 -179285
rect -84 -181847 84 -181813
rect -84 -181955 84 -181921
rect -84 -184483 84 -184449
rect -84 -184591 84 -184557
rect -84 -187119 84 -187085
rect -84 -187227 84 -187193
rect -84 -189755 84 -189721
rect -84 -189863 84 -189829
rect -84 -192391 84 -192357
rect -84 -192499 84 -192465
rect -84 -195027 84 -194993
rect -84 -195135 84 -195101
rect -84 -197663 84 -197629
rect -84 -197771 84 -197737
rect -84 -200299 84 -200265
rect -84 -200407 84 -200373
rect -84 -202935 84 -202901
rect -84 -203043 84 -203009
rect -84 -205571 84 -205537
rect -84 -205679 84 -205645
rect -84 -208207 84 -208173
rect -84 -208315 84 -208281
rect -84 -210843 84 -210809
rect -84 -210951 84 -210917
rect -84 -213479 84 -213445
rect -84 -213587 84 -213553
rect -84 -216115 84 -216081
rect -84 -216223 84 -216189
rect -84 -218751 84 -218717
rect -84 -218859 84 -218825
rect -84 -221387 84 -221353
rect -84 -221495 84 -221461
rect -84 -224023 84 -223989
rect -84 -224131 84 -224097
rect -84 -226659 84 -226625
rect -84 -226767 84 -226733
rect -84 -229295 84 -229261
rect -84 -229403 84 -229369
rect -84 -231931 84 -231897
rect -84 -232039 84 -232005
rect -84 -234567 84 -234533
rect -84 -234675 84 -234641
rect -84 -237203 84 -237169
rect -84 -237311 84 -237277
rect -84 -239839 84 -239805
rect -84 -239947 84 -239913
rect -84 -242475 84 -242441
rect -84 -242583 84 -242549
rect -84 -245111 84 -245077
rect -84 -245219 84 -245185
rect -84 -247747 84 -247713
rect -84 -247855 84 -247821
rect -84 -250383 84 -250349
rect -84 -250491 84 -250457
rect -84 -253019 84 -252985
rect -84 -253127 84 -253093
rect -84 -255655 84 -255621
rect -84 -255763 84 -255729
rect -84 -258291 84 -258257
rect -84 -258399 84 -258365
rect -84 -260927 84 -260893
rect -84 -261035 84 -261001
rect -84 -263563 84 -263529
rect -84 -263671 84 -263637
rect -84 -266199 84 -266165
rect -84 -266307 84 -266273
rect -84 -268835 84 -268801
rect -84 -268943 84 -268909
rect -84 -271471 84 -271437
rect -84 -271579 84 -271545
rect -84 -274107 84 -274073
rect -84 -274215 84 -274181
rect -84 -276743 84 -276709
rect -84 -276851 84 -276817
rect -84 -279379 84 -279345
rect -84 -279487 84 -279453
rect -84 -282015 84 -281981
rect -84 -282123 84 -282089
rect -84 -284651 84 -284617
rect -84 -284759 84 -284725
rect -84 -287287 84 -287253
rect -84 -287395 84 -287361
rect -84 -289923 84 -289889
rect -84 -290031 84 -289997
rect -84 -292559 84 -292525
rect -84 -292667 84 -292633
rect -84 -295195 84 -295161
rect -84 -295303 84 -295269
rect -84 -297831 84 -297797
rect -84 -297939 84 -297905
rect -84 -300467 84 -300433
rect -84 -300575 84 -300541
rect -84 -303103 84 -303069
rect -84 -303211 84 -303177
rect -84 -305739 84 -305705
rect -84 -305847 84 -305813
rect -84 -308375 84 -308341
rect -84 -308483 84 -308449
rect -84 -311011 84 -310977
rect -84 -311119 84 -311085
rect -84 -313647 84 -313613
rect -84 -313755 84 -313721
rect -84 -316283 84 -316249
rect -84 -316391 84 -316357
rect -84 -318919 84 -318885
rect -84 -319027 84 -318993
rect -84 -321555 84 -321521
rect -84 -321663 84 -321629
rect -84 -324191 84 -324157
rect -84 -324299 84 -324265
rect -84 -326827 84 -326793
rect -84 -326935 84 -326901
rect -84 -329463 84 -329429
rect -84 -329571 84 -329537
rect -84 -332099 84 -332065
rect -84 -332207 84 -332173
rect -84 -334735 84 -334701
rect -84 -334843 84 -334809
rect -84 -337371 84 -337337
<< locali >>
rect -280 337475 -184 337509
rect 184 337475 280 337509
rect -280 337413 -246 337475
rect 246 337413 280 337475
rect -100 337337 -84 337371
rect 84 337337 100 337371
rect -146 337278 -112 337294
rect -146 334886 -112 334902
rect 112 337278 146 337294
rect 112 334886 146 334902
rect -100 334809 -84 334843
rect 84 334809 100 334843
rect -100 334701 -84 334735
rect 84 334701 100 334735
rect -146 334642 -112 334658
rect -146 332250 -112 332266
rect 112 334642 146 334658
rect 112 332250 146 332266
rect -100 332173 -84 332207
rect 84 332173 100 332207
rect -100 332065 -84 332099
rect 84 332065 100 332099
rect -146 332006 -112 332022
rect -146 329614 -112 329630
rect 112 332006 146 332022
rect 112 329614 146 329630
rect -100 329537 -84 329571
rect 84 329537 100 329571
rect -100 329429 -84 329463
rect 84 329429 100 329463
rect -146 329370 -112 329386
rect -146 326978 -112 326994
rect 112 329370 146 329386
rect 112 326978 146 326994
rect -100 326901 -84 326935
rect 84 326901 100 326935
rect -100 326793 -84 326827
rect 84 326793 100 326827
rect -146 326734 -112 326750
rect -146 324342 -112 324358
rect 112 326734 146 326750
rect 112 324342 146 324358
rect -100 324265 -84 324299
rect 84 324265 100 324299
rect -100 324157 -84 324191
rect 84 324157 100 324191
rect -146 324098 -112 324114
rect -146 321706 -112 321722
rect 112 324098 146 324114
rect 112 321706 146 321722
rect -100 321629 -84 321663
rect 84 321629 100 321663
rect -100 321521 -84 321555
rect 84 321521 100 321555
rect -146 321462 -112 321478
rect -146 319070 -112 319086
rect 112 321462 146 321478
rect 112 319070 146 319086
rect -100 318993 -84 319027
rect 84 318993 100 319027
rect -100 318885 -84 318919
rect 84 318885 100 318919
rect -146 318826 -112 318842
rect -146 316434 -112 316450
rect 112 318826 146 318842
rect 112 316434 146 316450
rect -100 316357 -84 316391
rect 84 316357 100 316391
rect -100 316249 -84 316283
rect 84 316249 100 316283
rect -146 316190 -112 316206
rect -146 313798 -112 313814
rect 112 316190 146 316206
rect 112 313798 146 313814
rect -100 313721 -84 313755
rect 84 313721 100 313755
rect -100 313613 -84 313647
rect 84 313613 100 313647
rect -146 313554 -112 313570
rect -146 311162 -112 311178
rect 112 313554 146 313570
rect 112 311162 146 311178
rect -100 311085 -84 311119
rect 84 311085 100 311119
rect -100 310977 -84 311011
rect 84 310977 100 311011
rect -146 310918 -112 310934
rect -146 308526 -112 308542
rect 112 310918 146 310934
rect 112 308526 146 308542
rect -100 308449 -84 308483
rect 84 308449 100 308483
rect -100 308341 -84 308375
rect 84 308341 100 308375
rect -146 308282 -112 308298
rect -146 305890 -112 305906
rect 112 308282 146 308298
rect 112 305890 146 305906
rect -100 305813 -84 305847
rect 84 305813 100 305847
rect -100 305705 -84 305739
rect 84 305705 100 305739
rect -146 305646 -112 305662
rect -146 303254 -112 303270
rect 112 305646 146 305662
rect 112 303254 146 303270
rect -100 303177 -84 303211
rect 84 303177 100 303211
rect -100 303069 -84 303103
rect 84 303069 100 303103
rect -146 303010 -112 303026
rect -146 300618 -112 300634
rect 112 303010 146 303026
rect 112 300618 146 300634
rect -100 300541 -84 300575
rect 84 300541 100 300575
rect -100 300433 -84 300467
rect 84 300433 100 300467
rect -146 300374 -112 300390
rect -146 297982 -112 297998
rect 112 300374 146 300390
rect 112 297982 146 297998
rect -100 297905 -84 297939
rect 84 297905 100 297939
rect -100 297797 -84 297831
rect 84 297797 100 297831
rect -146 297738 -112 297754
rect -146 295346 -112 295362
rect 112 297738 146 297754
rect 112 295346 146 295362
rect -100 295269 -84 295303
rect 84 295269 100 295303
rect -100 295161 -84 295195
rect 84 295161 100 295195
rect -146 295102 -112 295118
rect -146 292710 -112 292726
rect 112 295102 146 295118
rect 112 292710 146 292726
rect -100 292633 -84 292667
rect 84 292633 100 292667
rect -100 292525 -84 292559
rect 84 292525 100 292559
rect -146 292466 -112 292482
rect -146 290074 -112 290090
rect 112 292466 146 292482
rect 112 290074 146 290090
rect -100 289997 -84 290031
rect 84 289997 100 290031
rect -100 289889 -84 289923
rect 84 289889 100 289923
rect -146 289830 -112 289846
rect -146 287438 -112 287454
rect 112 289830 146 289846
rect 112 287438 146 287454
rect -100 287361 -84 287395
rect 84 287361 100 287395
rect -100 287253 -84 287287
rect 84 287253 100 287287
rect -146 287194 -112 287210
rect -146 284802 -112 284818
rect 112 287194 146 287210
rect 112 284802 146 284818
rect -100 284725 -84 284759
rect 84 284725 100 284759
rect -100 284617 -84 284651
rect 84 284617 100 284651
rect -146 284558 -112 284574
rect -146 282166 -112 282182
rect 112 284558 146 284574
rect 112 282166 146 282182
rect -100 282089 -84 282123
rect 84 282089 100 282123
rect -100 281981 -84 282015
rect 84 281981 100 282015
rect -146 281922 -112 281938
rect -146 279530 -112 279546
rect 112 281922 146 281938
rect 112 279530 146 279546
rect -100 279453 -84 279487
rect 84 279453 100 279487
rect -100 279345 -84 279379
rect 84 279345 100 279379
rect -146 279286 -112 279302
rect -146 276894 -112 276910
rect 112 279286 146 279302
rect 112 276894 146 276910
rect -100 276817 -84 276851
rect 84 276817 100 276851
rect -100 276709 -84 276743
rect 84 276709 100 276743
rect -146 276650 -112 276666
rect -146 274258 -112 274274
rect 112 276650 146 276666
rect 112 274258 146 274274
rect -100 274181 -84 274215
rect 84 274181 100 274215
rect -100 274073 -84 274107
rect 84 274073 100 274107
rect -146 274014 -112 274030
rect -146 271622 -112 271638
rect 112 274014 146 274030
rect 112 271622 146 271638
rect -100 271545 -84 271579
rect 84 271545 100 271579
rect -100 271437 -84 271471
rect 84 271437 100 271471
rect -146 271378 -112 271394
rect -146 268986 -112 269002
rect 112 271378 146 271394
rect 112 268986 146 269002
rect -100 268909 -84 268943
rect 84 268909 100 268943
rect -100 268801 -84 268835
rect 84 268801 100 268835
rect -146 268742 -112 268758
rect -146 266350 -112 266366
rect 112 268742 146 268758
rect 112 266350 146 266366
rect -100 266273 -84 266307
rect 84 266273 100 266307
rect -100 266165 -84 266199
rect 84 266165 100 266199
rect -146 266106 -112 266122
rect -146 263714 -112 263730
rect 112 266106 146 266122
rect 112 263714 146 263730
rect -100 263637 -84 263671
rect 84 263637 100 263671
rect -100 263529 -84 263563
rect 84 263529 100 263563
rect -146 263470 -112 263486
rect -146 261078 -112 261094
rect 112 263470 146 263486
rect 112 261078 146 261094
rect -100 261001 -84 261035
rect 84 261001 100 261035
rect -100 260893 -84 260927
rect 84 260893 100 260927
rect -146 260834 -112 260850
rect -146 258442 -112 258458
rect 112 260834 146 260850
rect 112 258442 146 258458
rect -100 258365 -84 258399
rect 84 258365 100 258399
rect -100 258257 -84 258291
rect 84 258257 100 258291
rect -146 258198 -112 258214
rect -146 255806 -112 255822
rect 112 258198 146 258214
rect 112 255806 146 255822
rect -100 255729 -84 255763
rect 84 255729 100 255763
rect -100 255621 -84 255655
rect 84 255621 100 255655
rect -146 255562 -112 255578
rect -146 253170 -112 253186
rect 112 255562 146 255578
rect 112 253170 146 253186
rect -100 253093 -84 253127
rect 84 253093 100 253127
rect -100 252985 -84 253019
rect 84 252985 100 253019
rect -146 252926 -112 252942
rect -146 250534 -112 250550
rect 112 252926 146 252942
rect 112 250534 146 250550
rect -100 250457 -84 250491
rect 84 250457 100 250491
rect -100 250349 -84 250383
rect 84 250349 100 250383
rect -146 250290 -112 250306
rect -146 247898 -112 247914
rect 112 250290 146 250306
rect 112 247898 146 247914
rect -100 247821 -84 247855
rect 84 247821 100 247855
rect -100 247713 -84 247747
rect 84 247713 100 247747
rect -146 247654 -112 247670
rect -146 245262 -112 245278
rect 112 247654 146 247670
rect 112 245262 146 245278
rect -100 245185 -84 245219
rect 84 245185 100 245219
rect -100 245077 -84 245111
rect 84 245077 100 245111
rect -146 245018 -112 245034
rect -146 242626 -112 242642
rect 112 245018 146 245034
rect 112 242626 146 242642
rect -100 242549 -84 242583
rect 84 242549 100 242583
rect -100 242441 -84 242475
rect 84 242441 100 242475
rect -146 242382 -112 242398
rect -146 239990 -112 240006
rect 112 242382 146 242398
rect 112 239990 146 240006
rect -100 239913 -84 239947
rect 84 239913 100 239947
rect -100 239805 -84 239839
rect 84 239805 100 239839
rect -146 239746 -112 239762
rect -146 237354 -112 237370
rect 112 239746 146 239762
rect 112 237354 146 237370
rect -100 237277 -84 237311
rect 84 237277 100 237311
rect -100 237169 -84 237203
rect 84 237169 100 237203
rect -146 237110 -112 237126
rect -146 234718 -112 234734
rect 112 237110 146 237126
rect 112 234718 146 234734
rect -100 234641 -84 234675
rect 84 234641 100 234675
rect -100 234533 -84 234567
rect 84 234533 100 234567
rect -146 234474 -112 234490
rect -146 232082 -112 232098
rect 112 234474 146 234490
rect 112 232082 146 232098
rect -100 232005 -84 232039
rect 84 232005 100 232039
rect -100 231897 -84 231931
rect 84 231897 100 231931
rect -146 231838 -112 231854
rect -146 229446 -112 229462
rect 112 231838 146 231854
rect 112 229446 146 229462
rect -100 229369 -84 229403
rect 84 229369 100 229403
rect -100 229261 -84 229295
rect 84 229261 100 229295
rect -146 229202 -112 229218
rect -146 226810 -112 226826
rect 112 229202 146 229218
rect 112 226810 146 226826
rect -100 226733 -84 226767
rect 84 226733 100 226767
rect -100 226625 -84 226659
rect 84 226625 100 226659
rect -146 226566 -112 226582
rect -146 224174 -112 224190
rect 112 226566 146 226582
rect 112 224174 146 224190
rect -100 224097 -84 224131
rect 84 224097 100 224131
rect -100 223989 -84 224023
rect 84 223989 100 224023
rect -146 223930 -112 223946
rect -146 221538 -112 221554
rect 112 223930 146 223946
rect 112 221538 146 221554
rect -100 221461 -84 221495
rect 84 221461 100 221495
rect -100 221353 -84 221387
rect 84 221353 100 221387
rect -146 221294 -112 221310
rect -146 218902 -112 218918
rect 112 221294 146 221310
rect 112 218902 146 218918
rect -100 218825 -84 218859
rect 84 218825 100 218859
rect -100 218717 -84 218751
rect 84 218717 100 218751
rect -146 218658 -112 218674
rect -146 216266 -112 216282
rect 112 218658 146 218674
rect 112 216266 146 216282
rect -100 216189 -84 216223
rect 84 216189 100 216223
rect -100 216081 -84 216115
rect 84 216081 100 216115
rect -146 216022 -112 216038
rect -146 213630 -112 213646
rect 112 216022 146 216038
rect 112 213630 146 213646
rect -100 213553 -84 213587
rect 84 213553 100 213587
rect -100 213445 -84 213479
rect 84 213445 100 213479
rect -146 213386 -112 213402
rect -146 210994 -112 211010
rect 112 213386 146 213402
rect 112 210994 146 211010
rect -100 210917 -84 210951
rect 84 210917 100 210951
rect -100 210809 -84 210843
rect 84 210809 100 210843
rect -146 210750 -112 210766
rect -146 208358 -112 208374
rect 112 210750 146 210766
rect 112 208358 146 208374
rect -100 208281 -84 208315
rect 84 208281 100 208315
rect -100 208173 -84 208207
rect 84 208173 100 208207
rect -146 208114 -112 208130
rect -146 205722 -112 205738
rect 112 208114 146 208130
rect 112 205722 146 205738
rect -100 205645 -84 205679
rect 84 205645 100 205679
rect -100 205537 -84 205571
rect 84 205537 100 205571
rect -146 205478 -112 205494
rect -146 203086 -112 203102
rect 112 205478 146 205494
rect 112 203086 146 203102
rect -100 203009 -84 203043
rect 84 203009 100 203043
rect -100 202901 -84 202935
rect 84 202901 100 202935
rect -146 202842 -112 202858
rect -146 200450 -112 200466
rect 112 202842 146 202858
rect 112 200450 146 200466
rect -100 200373 -84 200407
rect 84 200373 100 200407
rect -100 200265 -84 200299
rect 84 200265 100 200299
rect -146 200206 -112 200222
rect -146 197814 -112 197830
rect 112 200206 146 200222
rect 112 197814 146 197830
rect -100 197737 -84 197771
rect 84 197737 100 197771
rect -100 197629 -84 197663
rect 84 197629 100 197663
rect -146 197570 -112 197586
rect -146 195178 -112 195194
rect 112 197570 146 197586
rect 112 195178 146 195194
rect -100 195101 -84 195135
rect 84 195101 100 195135
rect -100 194993 -84 195027
rect 84 194993 100 195027
rect -146 194934 -112 194950
rect -146 192542 -112 192558
rect 112 194934 146 194950
rect 112 192542 146 192558
rect -100 192465 -84 192499
rect 84 192465 100 192499
rect -100 192357 -84 192391
rect 84 192357 100 192391
rect -146 192298 -112 192314
rect -146 189906 -112 189922
rect 112 192298 146 192314
rect 112 189906 146 189922
rect -100 189829 -84 189863
rect 84 189829 100 189863
rect -100 189721 -84 189755
rect 84 189721 100 189755
rect -146 189662 -112 189678
rect -146 187270 -112 187286
rect 112 189662 146 189678
rect 112 187270 146 187286
rect -100 187193 -84 187227
rect 84 187193 100 187227
rect -100 187085 -84 187119
rect 84 187085 100 187119
rect -146 187026 -112 187042
rect -146 184634 -112 184650
rect 112 187026 146 187042
rect 112 184634 146 184650
rect -100 184557 -84 184591
rect 84 184557 100 184591
rect -100 184449 -84 184483
rect 84 184449 100 184483
rect -146 184390 -112 184406
rect -146 181998 -112 182014
rect 112 184390 146 184406
rect 112 181998 146 182014
rect -100 181921 -84 181955
rect 84 181921 100 181955
rect -100 181813 -84 181847
rect 84 181813 100 181847
rect -146 181754 -112 181770
rect -146 179362 -112 179378
rect 112 181754 146 181770
rect 112 179362 146 179378
rect -100 179285 -84 179319
rect 84 179285 100 179319
rect -100 179177 -84 179211
rect 84 179177 100 179211
rect -146 179118 -112 179134
rect -146 176726 -112 176742
rect 112 179118 146 179134
rect 112 176726 146 176742
rect -100 176649 -84 176683
rect 84 176649 100 176683
rect -100 176541 -84 176575
rect 84 176541 100 176575
rect -146 176482 -112 176498
rect -146 174090 -112 174106
rect 112 176482 146 176498
rect 112 174090 146 174106
rect -100 174013 -84 174047
rect 84 174013 100 174047
rect -100 173905 -84 173939
rect 84 173905 100 173939
rect -146 173846 -112 173862
rect -146 171454 -112 171470
rect 112 173846 146 173862
rect 112 171454 146 171470
rect -100 171377 -84 171411
rect 84 171377 100 171411
rect -100 171269 -84 171303
rect 84 171269 100 171303
rect -146 171210 -112 171226
rect -146 168818 -112 168834
rect 112 171210 146 171226
rect 112 168818 146 168834
rect -100 168741 -84 168775
rect 84 168741 100 168775
rect -100 168633 -84 168667
rect 84 168633 100 168667
rect -146 168574 -112 168590
rect -146 166182 -112 166198
rect 112 168574 146 168590
rect 112 166182 146 166198
rect -100 166105 -84 166139
rect 84 166105 100 166139
rect -100 165997 -84 166031
rect 84 165997 100 166031
rect -146 165938 -112 165954
rect -146 163546 -112 163562
rect 112 165938 146 165954
rect 112 163546 146 163562
rect -100 163469 -84 163503
rect 84 163469 100 163503
rect -100 163361 -84 163395
rect 84 163361 100 163395
rect -146 163302 -112 163318
rect -146 160910 -112 160926
rect 112 163302 146 163318
rect 112 160910 146 160926
rect -100 160833 -84 160867
rect 84 160833 100 160867
rect -100 160725 -84 160759
rect 84 160725 100 160759
rect -146 160666 -112 160682
rect -146 158274 -112 158290
rect 112 160666 146 160682
rect 112 158274 146 158290
rect -100 158197 -84 158231
rect 84 158197 100 158231
rect -100 158089 -84 158123
rect 84 158089 100 158123
rect -146 158030 -112 158046
rect -146 155638 -112 155654
rect 112 158030 146 158046
rect 112 155638 146 155654
rect -100 155561 -84 155595
rect 84 155561 100 155595
rect -100 155453 -84 155487
rect 84 155453 100 155487
rect -146 155394 -112 155410
rect -146 153002 -112 153018
rect 112 155394 146 155410
rect 112 153002 146 153018
rect -100 152925 -84 152959
rect 84 152925 100 152959
rect -100 152817 -84 152851
rect 84 152817 100 152851
rect -146 152758 -112 152774
rect -146 150366 -112 150382
rect 112 152758 146 152774
rect 112 150366 146 150382
rect -100 150289 -84 150323
rect 84 150289 100 150323
rect -100 150181 -84 150215
rect 84 150181 100 150215
rect -146 150122 -112 150138
rect -146 147730 -112 147746
rect 112 150122 146 150138
rect 112 147730 146 147746
rect -100 147653 -84 147687
rect 84 147653 100 147687
rect -100 147545 -84 147579
rect 84 147545 100 147579
rect -146 147486 -112 147502
rect -146 145094 -112 145110
rect 112 147486 146 147502
rect 112 145094 146 145110
rect -100 145017 -84 145051
rect 84 145017 100 145051
rect -100 144909 -84 144943
rect 84 144909 100 144943
rect -146 144850 -112 144866
rect -146 142458 -112 142474
rect 112 144850 146 144866
rect 112 142458 146 142474
rect -100 142381 -84 142415
rect 84 142381 100 142415
rect -100 142273 -84 142307
rect 84 142273 100 142307
rect -146 142214 -112 142230
rect -146 139822 -112 139838
rect 112 142214 146 142230
rect 112 139822 146 139838
rect -100 139745 -84 139779
rect 84 139745 100 139779
rect -100 139637 -84 139671
rect 84 139637 100 139671
rect -146 139578 -112 139594
rect -146 137186 -112 137202
rect 112 139578 146 139594
rect 112 137186 146 137202
rect -100 137109 -84 137143
rect 84 137109 100 137143
rect -100 137001 -84 137035
rect 84 137001 100 137035
rect -146 136942 -112 136958
rect -146 134550 -112 134566
rect 112 136942 146 136958
rect 112 134550 146 134566
rect -100 134473 -84 134507
rect 84 134473 100 134507
rect -100 134365 -84 134399
rect 84 134365 100 134399
rect -146 134306 -112 134322
rect -146 131914 -112 131930
rect 112 134306 146 134322
rect 112 131914 146 131930
rect -100 131837 -84 131871
rect 84 131837 100 131871
rect -100 131729 -84 131763
rect 84 131729 100 131763
rect -146 131670 -112 131686
rect -146 129278 -112 129294
rect 112 131670 146 131686
rect 112 129278 146 129294
rect -100 129201 -84 129235
rect 84 129201 100 129235
rect -100 129093 -84 129127
rect 84 129093 100 129127
rect -146 129034 -112 129050
rect -146 126642 -112 126658
rect 112 129034 146 129050
rect 112 126642 146 126658
rect -100 126565 -84 126599
rect 84 126565 100 126599
rect -100 126457 -84 126491
rect 84 126457 100 126491
rect -146 126398 -112 126414
rect -146 124006 -112 124022
rect 112 126398 146 126414
rect 112 124006 146 124022
rect -100 123929 -84 123963
rect 84 123929 100 123963
rect -100 123821 -84 123855
rect 84 123821 100 123855
rect -146 123762 -112 123778
rect -146 121370 -112 121386
rect 112 123762 146 123778
rect 112 121370 146 121386
rect -100 121293 -84 121327
rect 84 121293 100 121327
rect -100 121185 -84 121219
rect 84 121185 100 121219
rect -146 121126 -112 121142
rect -146 118734 -112 118750
rect 112 121126 146 121142
rect 112 118734 146 118750
rect -100 118657 -84 118691
rect 84 118657 100 118691
rect -100 118549 -84 118583
rect 84 118549 100 118583
rect -146 118490 -112 118506
rect -146 116098 -112 116114
rect 112 118490 146 118506
rect 112 116098 146 116114
rect -100 116021 -84 116055
rect 84 116021 100 116055
rect -100 115913 -84 115947
rect 84 115913 100 115947
rect -146 115854 -112 115870
rect -146 113462 -112 113478
rect 112 115854 146 115870
rect 112 113462 146 113478
rect -100 113385 -84 113419
rect 84 113385 100 113419
rect -100 113277 -84 113311
rect 84 113277 100 113311
rect -146 113218 -112 113234
rect -146 110826 -112 110842
rect 112 113218 146 113234
rect 112 110826 146 110842
rect -100 110749 -84 110783
rect 84 110749 100 110783
rect -100 110641 -84 110675
rect 84 110641 100 110675
rect -146 110582 -112 110598
rect -146 108190 -112 108206
rect 112 110582 146 110598
rect 112 108190 146 108206
rect -100 108113 -84 108147
rect 84 108113 100 108147
rect -100 108005 -84 108039
rect 84 108005 100 108039
rect -146 107946 -112 107962
rect -146 105554 -112 105570
rect 112 107946 146 107962
rect 112 105554 146 105570
rect -100 105477 -84 105511
rect 84 105477 100 105511
rect -100 105369 -84 105403
rect 84 105369 100 105403
rect -146 105310 -112 105326
rect -146 102918 -112 102934
rect 112 105310 146 105326
rect 112 102918 146 102934
rect -100 102841 -84 102875
rect 84 102841 100 102875
rect -100 102733 -84 102767
rect 84 102733 100 102767
rect -146 102674 -112 102690
rect -146 100282 -112 100298
rect 112 102674 146 102690
rect 112 100282 146 100298
rect -100 100205 -84 100239
rect 84 100205 100 100239
rect -100 100097 -84 100131
rect 84 100097 100 100131
rect -146 100038 -112 100054
rect -146 97646 -112 97662
rect 112 100038 146 100054
rect 112 97646 146 97662
rect -100 97569 -84 97603
rect 84 97569 100 97603
rect -100 97461 -84 97495
rect 84 97461 100 97495
rect -146 97402 -112 97418
rect -146 95010 -112 95026
rect 112 97402 146 97418
rect 112 95010 146 95026
rect -100 94933 -84 94967
rect 84 94933 100 94967
rect -100 94825 -84 94859
rect 84 94825 100 94859
rect -146 94766 -112 94782
rect -146 92374 -112 92390
rect 112 94766 146 94782
rect 112 92374 146 92390
rect -100 92297 -84 92331
rect 84 92297 100 92331
rect -100 92189 -84 92223
rect 84 92189 100 92223
rect -146 92130 -112 92146
rect -146 89738 -112 89754
rect 112 92130 146 92146
rect 112 89738 146 89754
rect -100 89661 -84 89695
rect 84 89661 100 89695
rect -100 89553 -84 89587
rect 84 89553 100 89587
rect -146 89494 -112 89510
rect -146 87102 -112 87118
rect 112 89494 146 89510
rect 112 87102 146 87118
rect -100 87025 -84 87059
rect 84 87025 100 87059
rect -100 86917 -84 86951
rect 84 86917 100 86951
rect -146 86858 -112 86874
rect -146 84466 -112 84482
rect 112 86858 146 86874
rect 112 84466 146 84482
rect -100 84389 -84 84423
rect 84 84389 100 84423
rect -100 84281 -84 84315
rect 84 84281 100 84315
rect -146 84222 -112 84238
rect -146 81830 -112 81846
rect 112 84222 146 84238
rect 112 81830 146 81846
rect -100 81753 -84 81787
rect 84 81753 100 81787
rect -100 81645 -84 81679
rect 84 81645 100 81679
rect -146 81586 -112 81602
rect -146 79194 -112 79210
rect 112 81586 146 81602
rect 112 79194 146 79210
rect -100 79117 -84 79151
rect 84 79117 100 79151
rect -100 79009 -84 79043
rect 84 79009 100 79043
rect -146 78950 -112 78966
rect -146 76558 -112 76574
rect 112 78950 146 78966
rect 112 76558 146 76574
rect -100 76481 -84 76515
rect 84 76481 100 76515
rect -100 76373 -84 76407
rect 84 76373 100 76407
rect -146 76314 -112 76330
rect -146 73922 -112 73938
rect 112 76314 146 76330
rect 112 73922 146 73938
rect -100 73845 -84 73879
rect 84 73845 100 73879
rect -100 73737 -84 73771
rect 84 73737 100 73771
rect -146 73678 -112 73694
rect -146 71286 -112 71302
rect 112 73678 146 73694
rect 112 71286 146 71302
rect -100 71209 -84 71243
rect 84 71209 100 71243
rect -100 71101 -84 71135
rect 84 71101 100 71135
rect -146 71042 -112 71058
rect -146 68650 -112 68666
rect 112 71042 146 71058
rect 112 68650 146 68666
rect -100 68573 -84 68607
rect 84 68573 100 68607
rect -100 68465 -84 68499
rect 84 68465 100 68499
rect -146 68406 -112 68422
rect -146 66014 -112 66030
rect 112 68406 146 68422
rect 112 66014 146 66030
rect -100 65937 -84 65971
rect 84 65937 100 65971
rect -100 65829 -84 65863
rect 84 65829 100 65863
rect -146 65770 -112 65786
rect -146 63378 -112 63394
rect 112 65770 146 65786
rect 112 63378 146 63394
rect -100 63301 -84 63335
rect 84 63301 100 63335
rect -100 63193 -84 63227
rect 84 63193 100 63227
rect -146 63134 -112 63150
rect -146 60742 -112 60758
rect 112 63134 146 63150
rect 112 60742 146 60758
rect -100 60665 -84 60699
rect 84 60665 100 60699
rect -100 60557 -84 60591
rect 84 60557 100 60591
rect -146 60498 -112 60514
rect -146 58106 -112 58122
rect 112 60498 146 60514
rect 112 58106 146 58122
rect -100 58029 -84 58063
rect 84 58029 100 58063
rect -100 57921 -84 57955
rect 84 57921 100 57955
rect -146 57862 -112 57878
rect -146 55470 -112 55486
rect 112 57862 146 57878
rect 112 55470 146 55486
rect -100 55393 -84 55427
rect 84 55393 100 55427
rect -100 55285 -84 55319
rect 84 55285 100 55319
rect -146 55226 -112 55242
rect -146 52834 -112 52850
rect 112 55226 146 55242
rect 112 52834 146 52850
rect -100 52757 -84 52791
rect 84 52757 100 52791
rect -100 52649 -84 52683
rect 84 52649 100 52683
rect -146 52590 -112 52606
rect -146 50198 -112 50214
rect 112 52590 146 52606
rect 112 50198 146 50214
rect -100 50121 -84 50155
rect 84 50121 100 50155
rect -100 50013 -84 50047
rect 84 50013 100 50047
rect -146 49954 -112 49970
rect -146 47562 -112 47578
rect 112 49954 146 49970
rect 112 47562 146 47578
rect -100 47485 -84 47519
rect 84 47485 100 47519
rect -100 47377 -84 47411
rect 84 47377 100 47411
rect -146 47318 -112 47334
rect -146 44926 -112 44942
rect 112 47318 146 47334
rect 112 44926 146 44942
rect -100 44849 -84 44883
rect 84 44849 100 44883
rect -100 44741 -84 44775
rect 84 44741 100 44775
rect -146 44682 -112 44698
rect -146 42290 -112 42306
rect 112 44682 146 44698
rect 112 42290 146 42306
rect -100 42213 -84 42247
rect 84 42213 100 42247
rect -100 42105 -84 42139
rect 84 42105 100 42139
rect -146 42046 -112 42062
rect -146 39654 -112 39670
rect 112 42046 146 42062
rect 112 39654 146 39670
rect -100 39577 -84 39611
rect 84 39577 100 39611
rect -100 39469 -84 39503
rect 84 39469 100 39503
rect -146 39410 -112 39426
rect -146 37018 -112 37034
rect 112 39410 146 39426
rect 112 37018 146 37034
rect -100 36941 -84 36975
rect 84 36941 100 36975
rect -100 36833 -84 36867
rect 84 36833 100 36867
rect -146 36774 -112 36790
rect -146 34382 -112 34398
rect 112 36774 146 36790
rect 112 34382 146 34398
rect -100 34305 -84 34339
rect 84 34305 100 34339
rect -100 34197 -84 34231
rect 84 34197 100 34231
rect -146 34138 -112 34154
rect -146 31746 -112 31762
rect 112 34138 146 34154
rect 112 31746 146 31762
rect -100 31669 -84 31703
rect 84 31669 100 31703
rect -100 31561 -84 31595
rect 84 31561 100 31595
rect -146 31502 -112 31518
rect -146 29110 -112 29126
rect 112 31502 146 31518
rect 112 29110 146 29126
rect -100 29033 -84 29067
rect 84 29033 100 29067
rect -100 28925 -84 28959
rect 84 28925 100 28959
rect -146 28866 -112 28882
rect -146 26474 -112 26490
rect 112 28866 146 28882
rect 112 26474 146 26490
rect -100 26397 -84 26431
rect 84 26397 100 26431
rect -100 26289 -84 26323
rect 84 26289 100 26323
rect -146 26230 -112 26246
rect -146 23838 -112 23854
rect 112 26230 146 26246
rect 112 23838 146 23854
rect -100 23761 -84 23795
rect 84 23761 100 23795
rect -100 23653 -84 23687
rect 84 23653 100 23687
rect -146 23594 -112 23610
rect -146 21202 -112 21218
rect 112 23594 146 23610
rect 112 21202 146 21218
rect -100 21125 -84 21159
rect 84 21125 100 21159
rect -100 21017 -84 21051
rect 84 21017 100 21051
rect -146 20958 -112 20974
rect -146 18566 -112 18582
rect 112 20958 146 20974
rect 112 18566 146 18582
rect -100 18489 -84 18523
rect 84 18489 100 18523
rect -100 18381 -84 18415
rect 84 18381 100 18415
rect -146 18322 -112 18338
rect -146 15930 -112 15946
rect 112 18322 146 18338
rect 112 15930 146 15946
rect -100 15853 -84 15887
rect 84 15853 100 15887
rect -100 15745 -84 15779
rect 84 15745 100 15779
rect -146 15686 -112 15702
rect -146 13294 -112 13310
rect 112 15686 146 15702
rect 112 13294 146 13310
rect -100 13217 -84 13251
rect 84 13217 100 13251
rect -100 13109 -84 13143
rect 84 13109 100 13143
rect -146 13050 -112 13066
rect -146 10658 -112 10674
rect 112 13050 146 13066
rect 112 10658 146 10674
rect -100 10581 -84 10615
rect 84 10581 100 10615
rect -100 10473 -84 10507
rect 84 10473 100 10507
rect -146 10414 -112 10430
rect -146 8022 -112 8038
rect 112 10414 146 10430
rect 112 8022 146 8038
rect -100 7945 -84 7979
rect 84 7945 100 7979
rect -100 7837 -84 7871
rect 84 7837 100 7871
rect -146 7778 -112 7794
rect -146 5386 -112 5402
rect 112 7778 146 7794
rect 112 5386 146 5402
rect -100 5309 -84 5343
rect 84 5309 100 5343
rect -100 5201 -84 5235
rect 84 5201 100 5235
rect -146 5142 -112 5158
rect -146 2750 -112 2766
rect 112 5142 146 5158
rect 112 2750 146 2766
rect -100 2673 -84 2707
rect 84 2673 100 2707
rect -100 2565 -84 2599
rect 84 2565 100 2599
rect -146 2506 -112 2522
rect -146 114 -112 130
rect 112 2506 146 2522
rect 112 114 146 130
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -130 -112 -114
rect -146 -2522 -112 -2506
rect 112 -130 146 -114
rect 112 -2522 146 -2506
rect -100 -2599 -84 -2565
rect 84 -2599 100 -2565
rect -100 -2707 -84 -2673
rect 84 -2707 100 -2673
rect -146 -2766 -112 -2750
rect -146 -5158 -112 -5142
rect 112 -2766 146 -2750
rect 112 -5158 146 -5142
rect -100 -5235 -84 -5201
rect 84 -5235 100 -5201
rect -100 -5343 -84 -5309
rect 84 -5343 100 -5309
rect -146 -5402 -112 -5386
rect -146 -7794 -112 -7778
rect 112 -5402 146 -5386
rect 112 -7794 146 -7778
rect -100 -7871 -84 -7837
rect 84 -7871 100 -7837
rect -100 -7979 -84 -7945
rect 84 -7979 100 -7945
rect -146 -8038 -112 -8022
rect -146 -10430 -112 -10414
rect 112 -8038 146 -8022
rect 112 -10430 146 -10414
rect -100 -10507 -84 -10473
rect 84 -10507 100 -10473
rect -100 -10615 -84 -10581
rect 84 -10615 100 -10581
rect -146 -10674 -112 -10658
rect -146 -13066 -112 -13050
rect 112 -10674 146 -10658
rect 112 -13066 146 -13050
rect -100 -13143 -84 -13109
rect 84 -13143 100 -13109
rect -100 -13251 -84 -13217
rect 84 -13251 100 -13217
rect -146 -13310 -112 -13294
rect -146 -15702 -112 -15686
rect 112 -13310 146 -13294
rect 112 -15702 146 -15686
rect -100 -15779 -84 -15745
rect 84 -15779 100 -15745
rect -100 -15887 -84 -15853
rect 84 -15887 100 -15853
rect -146 -15946 -112 -15930
rect -146 -18338 -112 -18322
rect 112 -15946 146 -15930
rect 112 -18338 146 -18322
rect -100 -18415 -84 -18381
rect 84 -18415 100 -18381
rect -100 -18523 -84 -18489
rect 84 -18523 100 -18489
rect -146 -18582 -112 -18566
rect -146 -20974 -112 -20958
rect 112 -18582 146 -18566
rect 112 -20974 146 -20958
rect -100 -21051 -84 -21017
rect 84 -21051 100 -21017
rect -100 -21159 -84 -21125
rect 84 -21159 100 -21125
rect -146 -21218 -112 -21202
rect -146 -23610 -112 -23594
rect 112 -21218 146 -21202
rect 112 -23610 146 -23594
rect -100 -23687 -84 -23653
rect 84 -23687 100 -23653
rect -100 -23795 -84 -23761
rect 84 -23795 100 -23761
rect -146 -23854 -112 -23838
rect -146 -26246 -112 -26230
rect 112 -23854 146 -23838
rect 112 -26246 146 -26230
rect -100 -26323 -84 -26289
rect 84 -26323 100 -26289
rect -100 -26431 -84 -26397
rect 84 -26431 100 -26397
rect -146 -26490 -112 -26474
rect -146 -28882 -112 -28866
rect 112 -26490 146 -26474
rect 112 -28882 146 -28866
rect -100 -28959 -84 -28925
rect 84 -28959 100 -28925
rect -100 -29067 -84 -29033
rect 84 -29067 100 -29033
rect -146 -29126 -112 -29110
rect -146 -31518 -112 -31502
rect 112 -29126 146 -29110
rect 112 -31518 146 -31502
rect -100 -31595 -84 -31561
rect 84 -31595 100 -31561
rect -100 -31703 -84 -31669
rect 84 -31703 100 -31669
rect -146 -31762 -112 -31746
rect -146 -34154 -112 -34138
rect 112 -31762 146 -31746
rect 112 -34154 146 -34138
rect -100 -34231 -84 -34197
rect 84 -34231 100 -34197
rect -100 -34339 -84 -34305
rect 84 -34339 100 -34305
rect -146 -34398 -112 -34382
rect -146 -36790 -112 -36774
rect 112 -34398 146 -34382
rect 112 -36790 146 -36774
rect -100 -36867 -84 -36833
rect 84 -36867 100 -36833
rect -100 -36975 -84 -36941
rect 84 -36975 100 -36941
rect -146 -37034 -112 -37018
rect -146 -39426 -112 -39410
rect 112 -37034 146 -37018
rect 112 -39426 146 -39410
rect -100 -39503 -84 -39469
rect 84 -39503 100 -39469
rect -100 -39611 -84 -39577
rect 84 -39611 100 -39577
rect -146 -39670 -112 -39654
rect -146 -42062 -112 -42046
rect 112 -39670 146 -39654
rect 112 -42062 146 -42046
rect -100 -42139 -84 -42105
rect 84 -42139 100 -42105
rect -100 -42247 -84 -42213
rect 84 -42247 100 -42213
rect -146 -42306 -112 -42290
rect -146 -44698 -112 -44682
rect 112 -42306 146 -42290
rect 112 -44698 146 -44682
rect -100 -44775 -84 -44741
rect 84 -44775 100 -44741
rect -100 -44883 -84 -44849
rect 84 -44883 100 -44849
rect -146 -44942 -112 -44926
rect -146 -47334 -112 -47318
rect 112 -44942 146 -44926
rect 112 -47334 146 -47318
rect -100 -47411 -84 -47377
rect 84 -47411 100 -47377
rect -100 -47519 -84 -47485
rect 84 -47519 100 -47485
rect -146 -47578 -112 -47562
rect -146 -49970 -112 -49954
rect 112 -47578 146 -47562
rect 112 -49970 146 -49954
rect -100 -50047 -84 -50013
rect 84 -50047 100 -50013
rect -100 -50155 -84 -50121
rect 84 -50155 100 -50121
rect -146 -50214 -112 -50198
rect -146 -52606 -112 -52590
rect 112 -50214 146 -50198
rect 112 -52606 146 -52590
rect -100 -52683 -84 -52649
rect 84 -52683 100 -52649
rect -100 -52791 -84 -52757
rect 84 -52791 100 -52757
rect -146 -52850 -112 -52834
rect -146 -55242 -112 -55226
rect 112 -52850 146 -52834
rect 112 -55242 146 -55226
rect -100 -55319 -84 -55285
rect 84 -55319 100 -55285
rect -100 -55427 -84 -55393
rect 84 -55427 100 -55393
rect -146 -55486 -112 -55470
rect -146 -57878 -112 -57862
rect 112 -55486 146 -55470
rect 112 -57878 146 -57862
rect -100 -57955 -84 -57921
rect 84 -57955 100 -57921
rect -100 -58063 -84 -58029
rect 84 -58063 100 -58029
rect -146 -58122 -112 -58106
rect -146 -60514 -112 -60498
rect 112 -58122 146 -58106
rect 112 -60514 146 -60498
rect -100 -60591 -84 -60557
rect 84 -60591 100 -60557
rect -100 -60699 -84 -60665
rect 84 -60699 100 -60665
rect -146 -60758 -112 -60742
rect -146 -63150 -112 -63134
rect 112 -60758 146 -60742
rect 112 -63150 146 -63134
rect -100 -63227 -84 -63193
rect 84 -63227 100 -63193
rect -100 -63335 -84 -63301
rect 84 -63335 100 -63301
rect -146 -63394 -112 -63378
rect -146 -65786 -112 -65770
rect 112 -63394 146 -63378
rect 112 -65786 146 -65770
rect -100 -65863 -84 -65829
rect 84 -65863 100 -65829
rect -100 -65971 -84 -65937
rect 84 -65971 100 -65937
rect -146 -66030 -112 -66014
rect -146 -68422 -112 -68406
rect 112 -66030 146 -66014
rect 112 -68422 146 -68406
rect -100 -68499 -84 -68465
rect 84 -68499 100 -68465
rect -100 -68607 -84 -68573
rect 84 -68607 100 -68573
rect -146 -68666 -112 -68650
rect -146 -71058 -112 -71042
rect 112 -68666 146 -68650
rect 112 -71058 146 -71042
rect -100 -71135 -84 -71101
rect 84 -71135 100 -71101
rect -100 -71243 -84 -71209
rect 84 -71243 100 -71209
rect -146 -71302 -112 -71286
rect -146 -73694 -112 -73678
rect 112 -71302 146 -71286
rect 112 -73694 146 -73678
rect -100 -73771 -84 -73737
rect 84 -73771 100 -73737
rect -100 -73879 -84 -73845
rect 84 -73879 100 -73845
rect -146 -73938 -112 -73922
rect -146 -76330 -112 -76314
rect 112 -73938 146 -73922
rect 112 -76330 146 -76314
rect -100 -76407 -84 -76373
rect 84 -76407 100 -76373
rect -100 -76515 -84 -76481
rect 84 -76515 100 -76481
rect -146 -76574 -112 -76558
rect -146 -78966 -112 -78950
rect 112 -76574 146 -76558
rect 112 -78966 146 -78950
rect -100 -79043 -84 -79009
rect 84 -79043 100 -79009
rect -100 -79151 -84 -79117
rect 84 -79151 100 -79117
rect -146 -79210 -112 -79194
rect -146 -81602 -112 -81586
rect 112 -79210 146 -79194
rect 112 -81602 146 -81586
rect -100 -81679 -84 -81645
rect 84 -81679 100 -81645
rect -100 -81787 -84 -81753
rect 84 -81787 100 -81753
rect -146 -81846 -112 -81830
rect -146 -84238 -112 -84222
rect 112 -81846 146 -81830
rect 112 -84238 146 -84222
rect -100 -84315 -84 -84281
rect 84 -84315 100 -84281
rect -100 -84423 -84 -84389
rect 84 -84423 100 -84389
rect -146 -84482 -112 -84466
rect -146 -86874 -112 -86858
rect 112 -84482 146 -84466
rect 112 -86874 146 -86858
rect -100 -86951 -84 -86917
rect 84 -86951 100 -86917
rect -100 -87059 -84 -87025
rect 84 -87059 100 -87025
rect -146 -87118 -112 -87102
rect -146 -89510 -112 -89494
rect 112 -87118 146 -87102
rect 112 -89510 146 -89494
rect -100 -89587 -84 -89553
rect 84 -89587 100 -89553
rect -100 -89695 -84 -89661
rect 84 -89695 100 -89661
rect -146 -89754 -112 -89738
rect -146 -92146 -112 -92130
rect 112 -89754 146 -89738
rect 112 -92146 146 -92130
rect -100 -92223 -84 -92189
rect 84 -92223 100 -92189
rect -100 -92331 -84 -92297
rect 84 -92331 100 -92297
rect -146 -92390 -112 -92374
rect -146 -94782 -112 -94766
rect 112 -92390 146 -92374
rect 112 -94782 146 -94766
rect -100 -94859 -84 -94825
rect 84 -94859 100 -94825
rect -100 -94967 -84 -94933
rect 84 -94967 100 -94933
rect -146 -95026 -112 -95010
rect -146 -97418 -112 -97402
rect 112 -95026 146 -95010
rect 112 -97418 146 -97402
rect -100 -97495 -84 -97461
rect 84 -97495 100 -97461
rect -100 -97603 -84 -97569
rect 84 -97603 100 -97569
rect -146 -97662 -112 -97646
rect -146 -100054 -112 -100038
rect 112 -97662 146 -97646
rect 112 -100054 146 -100038
rect -100 -100131 -84 -100097
rect 84 -100131 100 -100097
rect -100 -100239 -84 -100205
rect 84 -100239 100 -100205
rect -146 -100298 -112 -100282
rect -146 -102690 -112 -102674
rect 112 -100298 146 -100282
rect 112 -102690 146 -102674
rect -100 -102767 -84 -102733
rect 84 -102767 100 -102733
rect -100 -102875 -84 -102841
rect 84 -102875 100 -102841
rect -146 -102934 -112 -102918
rect -146 -105326 -112 -105310
rect 112 -102934 146 -102918
rect 112 -105326 146 -105310
rect -100 -105403 -84 -105369
rect 84 -105403 100 -105369
rect -100 -105511 -84 -105477
rect 84 -105511 100 -105477
rect -146 -105570 -112 -105554
rect -146 -107962 -112 -107946
rect 112 -105570 146 -105554
rect 112 -107962 146 -107946
rect -100 -108039 -84 -108005
rect 84 -108039 100 -108005
rect -100 -108147 -84 -108113
rect 84 -108147 100 -108113
rect -146 -108206 -112 -108190
rect -146 -110598 -112 -110582
rect 112 -108206 146 -108190
rect 112 -110598 146 -110582
rect -100 -110675 -84 -110641
rect 84 -110675 100 -110641
rect -100 -110783 -84 -110749
rect 84 -110783 100 -110749
rect -146 -110842 -112 -110826
rect -146 -113234 -112 -113218
rect 112 -110842 146 -110826
rect 112 -113234 146 -113218
rect -100 -113311 -84 -113277
rect 84 -113311 100 -113277
rect -100 -113419 -84 -113385
rect 84 -113419 100 -113385
rect -146 -113478 -112 -113462
rect -146 -115870 -112 -115854
rect 112 -113478 146 -113462
rect 112 -115870 146 -115854
rect -100 -115947 -84 -115913
rect 84 -115947 100 -115913
rect -100 -116055 -84 -116021
rect 84 -116055 100 -116021
rect -146 -116114 -112 -116098
rect -146 -118506 -112 -118490
rect 112 -116114 146 -116098
rect 112 -118506 146 -118490
rect -100 -118583 -84 -118549
rect 84 -118583 100 -118549
rect -100 -118691 -84 -118657
rect 84 -118691 100 -118657
rect -146 -118750 -112 -118734
rect -146 -121142 -112 -121126
rect 112 -118750 146 -118734
rect 112 -121142 146 -121126
rect -100 -121219 -84 -121185
rect 84 -121219 100 -121185
rect -100 -121327 -84 -121293
rect 84 -121327 100 -121293
rect -146 -121386 -112 -121370
rect -146 -123778 -112 -123762
rect 112 -121386 146 -121370
rect 112 -123778 146 -123762
rect -100 -123855 -84 -123821
rect 84 -123855 100 -123821
rect -100 -123963 -84 -123929
rect 84 -123963 100 -123929
rect -146 -124022 -112 -124006
rect -146 -126414 -112 -126398
rect 112 -124022 146 -124006
rect 112 -126414 146 -126398
rect -100 -126491 -84 -126457
rect 84 -126491 100 -126457
rect -100 -126599 -84 -126565
rect 84 -126599 100 -126565
rect -146 -126658 -112 -126642
rect -146 -129050 -112 -129034
rect 112 -126658 146 -126642
rect 112 -129050 146 -129034
rect -100 -129127 -84 -129093
rect 84 -129127 100 -129093
rect -100 -129235 -84 -129201
rect 84 -129235 100 -129201
rect -146 -129294 -112 -129278
rect -146 -131686 -112 -131670
rect 112 -129294 146 -129278
rect 112 -131686 146 -131670
rect -100 -131763 -84 -131729
rect 84 -131763 100 -131729
rect -100 -131871 -84 -131837
rect 84 -131871 100 -131837
rect -146 -131930 -112 -131914
rect -146 -134322 -112 -134306
rect 112 -131930 146 -131914
rect 112 -134322 146 -134306
rect -100 -134399 -84 -134365
rect 84 -134399 100 -134365
rect -100 -134507 -84 -134473
rect 84 -134507 100 -134473
rect -146 -134566 -112 -134550
rect -146 -136958 -112 -136942
rect 112 -134566 146 -134550
rect 112 -136958 146 -136942
rect -100 -137035 -84 -137001
rect 84 -137035 100 -137001
rect -100 -137143 -84 -137109
rect 84 -137143 100 -137109
rect -146 -137202 -112 -137186
rect -146 -139594 -112 -139578
rect 112 -137202 146 -137186
rect 112 -139594 146 -139578
rect -100 -139671 -84 -139637
rect 84 -139671 100 -139637
rect -100 -139779 -84 -139745
rect 84 -139779 100 -139745
rect -146 -139838 -112 -139822
rect -146 -142230 -112 -142214
rect 112 -139838 146 -139822
rect 112 -142230 146 -142214
rect -100 -142307 -84 -142273
rect 84 -142307 100 -142273
rect -100 -142415 -84 -142381
rect 84 -142415 100 -142381
rect -146 -142474 -112 -142458
rect -146 -144866 -112 -144850
rect 112 -142474 146 -142458
rect 112 -144866 146 -144850
rect -100 -144943 -84 -144909
rect 84 -144943 100 -144909
rect -100 -145051 -84 -145017
rect 84 -145051 100 -145017
rect -146 -145110 -112 -145094
rect -146 -147502 -112 -147486
rect 112 -145110 146 -145094
rect 112 -147502 146 -147486
rect -100 -147579 -84 -147545
rect 84 -147579 100 -147545
rect -100 -147687 -84 -147653
rect 84 -147687 100 -147653
rect -146 -147746 -112 -147730
rect -146 -150138 -112 -150122
rect 112 -147746 146 -147730
rect 112 -150138 146 -150122
rect -100 -150215 -84 -150181
rect 84 -150215 100 -150181
rect -100 -150323 -84 -150289
rect 84 -150323 100 -150289
rect -146 -150382 -112 -150366
rect -146 -152774 -112 -152758
rect 112 -150382 146 -150366
rect 112 -152774 146 -152758
rect -100 -152851 -84 -152817
rect 84 -152851 100 -152817
rect -100 -152959 -84 -152925
rect 84 -152959 100 -152925
rect -146 -153018 -112 -153002
rect -146 -155410 -112 -155394
rect 112 -153018 146 -153002
rect 112 -155410 146 -155394
rect -100 -155487 -84 -155453
rect 84 -155487 100 -155453
rect -100 -155595 -84 -155561
rect 84 -155595 100 -155561
rect -146 -155654 -112 -155638
rect -146 -158046 -112 -158030
rect 112 -155654 146 -155638
rect 112 -158046 146 -158030
rect -100 -158123 -84 -158089
rect 84 -158123 100 -158089
rect -100 -158231 -84 -158197
rect 84 -158231 100 -158197
rect -146 -158290 -112 -158274
rect -146 -160682 -112 -160666
rect 112 -158290 146 -158274
rect 112 -160682 146 -160666
rect -100 -160759 -84 -160725
rect 84 -160759 100 -160725
rect -100 -160867 -84 -160833
rect 84 -160867 100 -160833
rect -146 -160926 -112 -160910
rect -146 -163318 -112 -163302
rect 112 -160926 146 -160910
rect 112 -163318 146 -163302
rect -100 -163395 -84 -163361
rect 84 -163395 100 -163361
rect -100 -163503 -84 -163469
rect 84 -163503 100 -163469
rect -146 -163562 -112 -163546
rect -146 -165954 -112 -165938
rect 112 -163562 146 -163546
rect 112 -165954 146 -165938
rect -100 -166031 -84 -165997
rect 84 -166031 100 -165997
rect -100 -166139 -84 -166105
rect 84 -166139 100 -166105
rect -146 -166198 -112 -166182
rect -146 -168590 -112 -168574
rect 112 -166198 146 -166182
rect 112 -168590 146 -168574
rect -100 -168667 -84 -168633
rect 84 -168667 100 -168633
rect -100 -168775 -84 -168741
rect 84 -168775 100 -168741
rect -146 -168834 -112 -168818
rect -146 -171226 -112 -171210
rect 112 -168834 146 -168818
rect 112 -171226 146 -171210
rect -100 -171303 -84 -171269
rect 84 -171303 100 -171269
rect -100 -171411 -84 -171377
rect 84 -171411 100 -171377
rect -146 -171470 -112 -171454
rect -146 -173862 -112 -173846
rect 112 -171470 146 -171454
rect 112 -173862 146 -173846
rect -100 -173939 -84 -173905
rect 84 -173939 100 -173905
rect -100 -174047 -84 -174013
rect 84 -174047 100 -174013
rect -146 -174106 -112 -174090
rect -146 -176498 -112 -176482
rect 112 -174106 146 -174090
rect 112 -176498 146 -176482
rect -100 -176575 -84 -176541
rect 84 -176575 100 -176541
rect -100 -176683 -84 -176649
rect 84 -176683 100 -176649
rect -146 -176742 -112 -176726
rect -146 -179134 -112 -179118
rect 112 -176742 146 -176726
rect 112 -179134 146 -179118
rect -100 -179211 -84 -179177
rect 84 -179211 100 -179177
rect -100 -179319 -84 -179285
rect 84 -179319 100 -179285
rect -146 -179378 -112 -179362
rect -146 -181770 -112 -181754
rect 112 -179378 146 -179362
rect 112 -181770 146 -181754
rect -100 -181847 -84 -181813
rect 84 -181847 100 -181813
rect -100 -181955 -84 -181921
rect 84 -181955 100 -181921
rect -146 -182014 -112 -181998
rect -146 -184406 -112 -184390
rect 112 -182014 146 -181998
rect 112 -184406 146 -184390
rect -100 -184483 -84 -184449
rect 84 -184483 100 -184449
rect -100 -184591 -84 -184557
rect 84 -184591 100 -184557
rect -146 -184650 -112 -184634
rect -146 -187042 -112 -187026
rect 112 -184650 146 -184634
rect 112 -187042 146 -187026
rect -100 -187119 -84 -187085
rect 84 -187119 100 -187085
rect -100 -187227 -84 -187193
rect 84 -187227 100 -187193
rect -146 -187286 -112 -187270
rect -146 -189678 -112 -189662
rect 112 -187286 146 -187270
rect 112 -189678 146 -189662
rect -100 -189755 -84 -189721
rect 84 -189755 100 -189721
rect -100 -189863 -84 -189829
rect 84 -189863 100 -189829
rect -146 -189922 -112 -189906
rect -146 -192314 -112 -192298
rect 112 -189922 146 -189906
rect 112 -192314 146 -192298
rect -100 -192391 -84 -192357
rect 84 -192391 100 -192357
rect -100 -192499 -84 -192465
rect 84 -192499 100 -192465
rect -146 -192558 -112 -192542
rect -146 -194950 -112 -194934
rect 112 -192558 146 -192542
rect 112 -194950 146 -194934
rect -100 -195027 -84 -194993
rect 84 -195027 100 -194993
rect -100 -195135 -84 -195101
rect 84 -195135 100 -195101
rect -146 -195194 -112 -195178
rect -146 -197586 -112 -197570
rect 112 -195194 146 -195178
rect 112 -197586 146 -197570
rect -100 -197663 -84 -197629
rect 84 -197663 100 -197629
rect -100 -197771 -84 -197737
rect 84 -197771 100 -197737
rect -146 -197830 -112 -197814
rect -146 -200222 -112 -200206
rect 112 -197830 146 -197814
rect 112 -200222 146 -200206
rect -100 -200299 -84 -200265
rect 84 -200299 100 -200265
rect -100 -200407 -84 -200373
rect 84 -200407 100 -200373
rect -146 -200466 -112 -200450
rect -146 -202858 -112 -202842
rect 112 -200466 146 -200450
rect 112 -202858 146 -202842
rect -100 -202935 -84 -202901
rect 84 -202935 100 -202901
rect -100 -203043 -84 -203009
rect 84 -203043 100 -203009
rect -146 -203102 -112 -203086
rect -146 -205494 -112 -205478
rect 112 -203102 146 -203086
rect 112 -205494 146 -205478
rect -100 -205571 -84 -205537
rect 84 -205571 100 -205537
rect -100 -205679 -84 -205645
rect 84 -205679 100 -205645
rect -146 -205738 -112 -205722
rect -146 -208130 -112 -208114
rect 112 -205738 146 -205722
rect 112 -208130 146 -208114
rect -100 -208207 -84 -208173
rect 84 -208207 100 -208173
rect -100 -208315 -84 -208281
rect 84 -208315 100 -208281
rect -146 -208374 -112 -208358
rect -146 -210766 -112 -210750
rect 112 -208374 146 -208358
rect 112 -210766 146 -210750
rect -100 -210843 -84 -210809
rect 84 -210843 100 -210809
rect -100 -210951 -84 -210917
rect 84 -210951 100 -210917
rect -146 -211010 -112 -210994
rect -146 -213402 -112 -213386
rect 112 -211010 146 -210994
rect 112 -213402 146 -213386
rect -100 -213479 -84 -213445
rect 84 -213479 100 -213445
rect -100 -213587 -84 -213553
rect 84 -213587 100 -213553
rect -146 -213646 -112 -213630
rect -146 -216038 -112 -216022
rect 112 -213646 146 -213630
rect 112 -216038 146 -216022
rect -100 -216115 -84 -216081
rect 84 -216115 100 -216081
rect -100 -216223 -84 -216189
rect 84 -216223 100 -216189
rect -146 -216282 -112 -216266
rect -146 -218674 -112 -218658
rect 112 -216282 146 -216266
rect 112 -218674 146 -218658
rect -100 -218751 -84 -218717
rect 84 -218751 100 -218717
rect -100 -218859 -84 -218825
rect 84 -218859 100 -218825
rect -146 -218918 -112 -218902
rect -146 -221310 -112 -221294
rect 112 -218918 146 -218902
rect 112 -221310 146 -221294
rect -100 -221387 -84 -221353
rect 84 -221387 100 -221353
rect -100 -221495 -84 -221461
rect 84 -221495 100 -221461
rect -146 -221554 -112 -221538
rect -146 -223946 -112 -223930
rect 112 -221554 146 -221538
rect 112 -223946 146 -223930
rect -100 -224023 -84 -223989
rect 84 -224023 100 -223989
rect -100 -224131 -84 -224097
rect 84 -224131 100 -224097
rect -146 -224190 -112 -224174
rect -146 -226582 -112 -226566
rect 112 -224190 146 -224174
rect 112 -226582 146 -226566
rect -100 -226659 -84 -226625
rect 84 -226659 100 -226625
rect -100 -226767 -84 -226733
rect 84 -226767 100 -226733
rect -146 -226826 -112 -226810
rect -146 -229218 -112 -229202
rect 112 -226826 146 -226810
rect 112 -229218 146 -229202
rect -100 -229295 -84 -229261
rect 84 -229295 100 -229261
rect -100 -229403 -84 -229369
rect 84 -229403 100 -229369
rect -146 -229462 -112 -229446
rect -146 -231854 -112 -231838
rect 112 -229462 146 -229446
rect 112 -231854 146 -231838
rect -100 -231931 -84 -231897
rect 84 -231931 100 -231897
rect -100 -232039 -84 -232005
rect 84 -232039 100 -232005
rect -146 -232098 -112 -232082
rect -146 -234490 -112 -234474
rect 112 -232098 146 -232082
rect 112 -234490 146 -234474
rect -100 -234567 -84 -234533
rect 84 -234567 100 -234533
rect -100 -234675 -84 -234641
rect 84 -234675 100 -234641
rect -146 -234734 -112 -234718
rect -146 -237126 -112 -237110
rect 112 -234734 146 -234718
rect 112 -237126 146 -237110
rect -100 -237203 -84 -237169
rect 84 -237203 100 -237169
rect -100 -237311 -84 -237277
rect 84 -237311 100 -237277
rect -146 -237370 -112 -237354
rect -146 -239762 -112 -239746
rect 112 -237370 146 -237354
rect 112 -239762 146 -239746
rect -100 -239839 -84 -239805
rect 84 -239839 100 -239805
rect -100 -239947 -84 -239913
rect 84 -239947 100 -239913
rect -146 -240006 -112 -239990
rect -146 -242398 -112 -242382
rect 112 -240006 146 -239990
rect 112 -242398 146 -242382
rect -100 -242475 -84 -242441
rect 84 -242475 100 -242441
rect -100 -242583 -84 -242549
rect 84 -242583 100 -242549
rect -146 -242642 -112 -242626
rect -146 -245034 -112 -245018
rect 112 -242642 146 -242626
rect 112 -245034 146 -245018
rect -100 -245111 -84 -245077
rect 84 -245111 100 -245077
rect -100 -245219 -84 -245185
rect 84 -245219 100 -245185
rect -146 -245278 -112 -245262
rect -146 -247670 -112 -247654
rect 112 -245278 146 -245262
rect 112 -247670 146 -247654
rect -100 -247747 -84 -247713
rect 84 -247747 100 -247713
rect -100 -247855 -84 -247821
rect 84 -247855 100 -247821
rect -146 -247914 -112 -247898
rect -146 -250306 -112 -250290
rect 112 -247914 146 -247898
rect 112 -250306 146 -250290
rect -100 -250383 -84 -250349
rect 84 -250383 100 -250349
rect -100 -250491 -84 -250457
rect 84 -250491 100 -250457
rect -146 -250550 -112 -250534
rect -146 -252942 -112 -252926
rect 112 -250550 146 -250534
rect 112 -252942 146 -252926
rect -100 -253019 -84 -252985
rect 84 -253019 100 -252985
rect -100 -253127 -84 -253093
rect 84 -253127 100 -253093
rect -146 -253186 -112 -253170
rect -146 -255578 -112 -255562
rect 112 -253186 146 -253170
rect 112 -255578 146 -255562
rect -100 -255655 -84 -255621
rect 84 -255655 100 -255621
rect -100 -255763 -84 -255729
rect 84 -255763 100 -255729
rect -146 -255822 -112 -255806
rect -146 -258214 -112 -258198
rect 112 -255822 146 -255806
rect 112 -258214 146 -258198
rect -100 -258291 -84 -258257
rect 84 -258291 100 -258257
rect -100 -258399 -84 -258365
rect 84 -258399 100 -258365
rect -146 -258458 -112 -258442
rect -146 -260850 -112 -260834
rect 112 -258458 146 -258442
rect 112 -260850 146 -260834
rect -100 -260927 -84 -260893
rect 84 -260927 100 -260893
rect -100 -261035 -84 -261001
rect 84 -261035 100 -261001
rect -146 -261094 -112 -261078
rect -146 -263486 -112 -263470
rect 112 -261094 146 -261078
rect 112 -263486 146 -263470
rect -100 -263563 -84 -263529
rect 84 -263563 100 -263529
rect -100 -263671 -84 -263637
rect 84 -263671 100 -263637
rect -146 -263730 -112 -263714
rect -146 -266122 -112 -266106
rect 112 -263730 146 -263714
rect 112 -266122 146 -266106
rect -100 -266199 -84 -266165
rect 84 -266199 100 -266165
rect -100 -266307 -84 -266273
rect 84 -266307 100 -266273
rect -146 -266366 -112 -266350
rect -146 -268758 -112 -268742
rect 112 -266366 146 -266350
rect 112 -268758 146 -268742
rect -100 -268835 -84 -268801
rect 84 -268835 100 -268801
rect -100 -268943 -84 -268909
rect 84 -268943 100 -268909
rect -146 -269002 -112 -268986
rect -146 -271394 -112 -271378
rect 112 -269002 146 -268986
rect 112 -271394 146 -271378
rect -100 -271471 -84 -271437
rect 84 -271471 100 -271437
rect -100 -271579 -84 -271545
rect 84 -271579 100 -271545
rect -146 -271638 -112 -271622
rect -146 -274030 -112 -274014
rect 112 -271638 146 -271622
rect 112 -274030 146 -274014
rect -100 -274107 -84 -274073
rect 84 -274107 100 -274073
rect -100 -274215 -84 -274181
rect 84 -274215 100 -274181
rect -146 -274274 -112 -274258
rect -146 -276666 -112 -276650
rect 112 -274274 146 -274258
rect 112 -276666 146 -276650
rect -100 -276743 -84 -276709
rect 84 -276743 100 -276709
rect -100 -276851 -84 -276817
rect 84 -276851 100 -276817
rect -146 -276910 -112 -276894
rect -146 -279302 -112 -279286
rect 112 -276910 146 -276894
rect 112 -279302 146 -279286
rect -100 -279379 -84 -279345
rect 84 -279379 100 -279345
rect -100 -279487 -84 -279453
rect 84 -279487 100 -279453
rect -146 -279546 -112 -279530
rect -146 -281938 -112 -281922
rect 112 -279546 146 -279530
rect 112 -281938 146 -281922
rect -100 -282015 -84 -281981
rect 84 -282015 100 -281981
rect -100 -282123 -84 -282089
rect 84 -282123 100 -282089
rect -146 -282182 -112 -282166
rect -146 -284574 -112 -284558
rect 112 -282182 146 -282166
rect 112 -284574 146 -284558
rect -100 -284651 -84 -284617
rect 84 -284651 100 -284617
rect -100 -284759 -84 -284725
rect 84 -284759 100 -284725
rect -146 -284818 -112 -284802
rect -146 -287210 -112 -287194
rect 112 -284818 146 -284802
rect 112 -287210 146 -287194
rect -100 -287287 -84 -287253
rect 84 -287287 100 -287253
rect -100 -287395 -84 -287361
rect 84 -287395 100 -287361
rect -146 -287454 -112 -287438
rect -146 -289846 -112 -289830
rect 112 -287454 146 -287438
rect 112 -289846 146 -289830
rect -100 -289923 -84 -289889
rect 84 -289923 100 -289889
rect -100 -290031 -84 -289997
rect 84 -290031 100 -289997
rect -146 -290090 -112 -290074
rect -146 -292482 -112 -292466
rect 112 -290090 146 -290074
rect 112 -292482 146 -292466
rect -100 -292559 -84 -292525
rect 84 -292559 100 -292525
rect -100 -292667 -84 -292633
rect 84 -292667 100 -292633
rect -146 -292726 -112 -292710
rect -146 -295118 -112 -295102
rect 112 -292726 146 -292710
rect 112 -295118 146 -295102
rect -100 -295195 -84 -295161
rect 84 -295195 100 -295161
rect -100 -295303 -84 -295269
rect 84 -295303 100 -295269
rect -146 -295362 -112 -295346
rect -146 -297754 -112 -297738
rect 112 -295362 146 -295346
rect 112 -297754 146 -297738
rect -100 -297831 -84 -297797
rect 84 -297831 100 -297797
rect -100 -297939 -84 -297905
rect 84 -297939 100 -297905
rect -146 -297998 -112 -297982
rect -146 -300390 -112 -300374
rect 112 -297998 146 -297982
rect 112 -300390 146 -300374
rect -100 -300467 -84 -300433
rect 84 -300467 100 -300433
rect -100 -300575 -84 -300541
rect 84 -300575 100 -300541
rect -146 -300634 -112 -300618
rect -146 -303026 -112 -303010
rect 112 -300634 146 -300618
rect 112 -303026 146 -303010
rect -100 -303103 -84 -303069
rect 84 -303103 100 -303069
rect -100 -303211 -84 -303177
rect 84 -303211 100 -303177
rect -146 -303270 -112 -303254
rect -146 -305662 -112 -305646
rect 112 -303270 146 -303254
rect 112 -305662 146 -305646
rect -100 -305739 -84 -305705
rect 84 -305739 100 -305705
rect -100 -305847 -84 -305813
rect 84 -305847 100 -305813
rect -146 -305906 -112 -305890
rect -146 -308298 -112 -308282
rect 112 -305906 146 -305890
rect 112 -308298 146 -308282
rect -100 -308375 -84 -308341
rect 84 -308375 100 -308341
rect -100 -308483 -84 -308449
rect 84 -308483 100 -308449
rect -146 -308542 -112 -308526
rect -146 -310934 -112 -310918
rect 112 -308542 146 -308526
rect 112 -310934 146 -310918
rect -100 -311011 -84 -310977
rect 84 -311011 100 -310977
rect -100 -311119 -84 -311085
rect 84 -311119 100 -311085
rect -146 -311178 -112 -311162
rect -146 -313570 -112 -313554
rect 112 -311178 146 -311162
rect 112 -313570 146 -313554
rect -100 -313647 -84 -313613
rect 84 -313647 100 -313613
rect -100 -313755 -84 -313721
rect 84 -313755 100 -313721
rect -146 -313814 -112 -313798
rect -146 -316206 -112 -316190
rect 112 -313814 146 -313798
rect 112 -316206 146 -316190
rect -100 -316283 -84 -316249
rect 84 -316283 100 -316249
rect -100 -316391 -84 -316357
rect 84 -316391 100 -316357
rect -146 -316450 -112 -316434
rect -146 -318842 -112 -318826
rect 112 -316450 146 -316434
rect 112 -318842 146 -318826
rect -100 -318919 -84 -318885
rect 84 -318919 100 -318885
rect -100 -319027 -84 -318993
rect 84 -319027 100 -318993
rect -146 -319086 -112 -319070
rect -146 -321478 -112 -321462
rect 112 -319086 146 -319070
rect 112 -321478 146 -321462
rect -100 -321555 -84 -321521
rect 84 -321555 100 -321521
rect -100 -321663 -84 -321629
rect 84 -321663 100 -321629
rect -146 -321722 -112 -321706
rect -146 -324114 -112 -324098
rect 112 -321722 146 -321706
rect 112 -324114 146 -324098
rect -100 -324191 -84 -324157
rect 84 -324191 100 -324157
rect -100 -324299 -84 -324265
rect 84 -324299 100 -324265
rect -146 -324358 -112 -324342
rect -146 -326750 -112 -326734
rect 112 -324358 146 -324342
rect 112 -326750 146 -326734
rect -100 -326827 -84 -326793
rect 84 -326827 100 -326793
rect -100 -326935 -84 -326901
rect 84 -326935 100 -326901
rect -146 -326994 -112 -326978
rect -146 -329386 -112 -329370
rect 112 -326994 146 -326978
rect 112 -329386 146 -329370
rect -100 -329463 -84 -329429
rect 84 -329463 100 -329429
rect -100 -329571 -84 -329537
rect 84 -329571 100 -329537
rect -146 -329630 -112 -329614
rect -146 -332022 -112 -332006
rect 112 -329630 146 -329614
rect 112 -332022 146 -332006
rect -100 -332099 -84 -332065
rect 84 -332099 100 -332065
rect -100 -332207 -84 -332173
rect 84 -332207 100 -332173
rect -146 -332266 -112 -332250
rect -146 -334658 -112 -334642
rect 112 -332266 146 -332250
rect 112 -334658 146 -334642
rect -100 -334735 -84 -334701
rect 84 -334735 100 -334701
rect -100 -334843 -84 -334809
rect 84 -334843 100 -334809
rect -146 -334902 -112 -334886
rect -146 -337294 -112 -337278
rect 112 -334902 146 -334886
rect 112 -337294 146 -337278
rect -100 -337371 -84 -337337
rect 84 -337371 100 -337337
rect -280 -337475 -246 -337413
rect 246 -337475 280 -337413
rect -280 -337509 -184 -337475
rect 184 -337509 280 -337475
<< viali >>
rect -84 337337 84 337371
rect -146 334902 -112 337278
rect 112 334902 146 337278
rect -84 334809 84 334843
rect -84 334701 84 334735
rect -146 332266 -112 334642
rect 112 332266 146 334642
rect -84 332173 84 332207
rect -84 332065 84 332099
rect -146 329630 -112 332006
rect 112 329630 146 332006
rect -84 329537 84 329571
rect -84 329429 84 329463
rect -146 326994 -112 329370
rect 112 326994 146 329370
rect -84 326901 84 326935
rect -84 326793 84 326827
rect -146 324358 -112 326734
rect 112 324358 146 326734
rect -84 324265 84 324299
rect -84 324157 84 324191
rect -146 321722 -112 324098
rect 112 321722 146 324098
rect -84 321629 84 321663
rect -84 321521 84 321555
rect -146 319086 -112 321462
rect 112 319086 146 321462
rect -84 318993 84 319027
rect -84 318885 84 318919
rect -146 316450 -112 318826
rect 112 316450 146 318826
rect -84 316357 84 316391
rect -84 316249 84 316283
rect -146 313814 -112 316190
rect 112 313814 146 316190
rect -84 313721 84 313755
rect -84 313613 84 313647
rect -146 311178 -112 313554
rect 112 311178 146 313554
rect -84 311085 84 311119
rect -84 310977 84 311011
rect -146 308542 -112 310918
rect 112 308542 146 310918
rect -84 308449 84 308483
rect -84 308341 84 308375
rect -146 305906 -112 308282
rect 112 305906 146 308282
rect -84 305813 84 305847
rect -84 305705 84 305739
rect -146 303270 -112 305646
rect 112 303270 146 305646
rect -84 303177 84 303211
rect -84 303069 84 303103
rect -146 300634 -112 303010
rect 112 300634 146 303010
rect -84 300541 84 300575
rect -84 300433 84 300467
rect -146 297998 -112 300374
rect 112 297998 146 300374
rect -84 297905 84 297939
rect -84 297797 84 297831
rect -146 295362 -112 297738
rect 112 295362 146 297738
rect -84 295269 84 295303
rect -84 295161 84 295195
rect -146 292726 -112 295102
rect 112 292726 146 295102
rect -84 292633 84 292667
rect -84 292525 84 292559
rect -146 290090 -112 292466
rect 112 290090 146 292466
rect -84 289997 84 290031
rect -84 289889 84 289923
rect -146 287454 -112 289830
rect 112 287454 146 289830
rect -84 287361 84 287395
rect -84 287253 84 287287
rect -146 284818 -112 287194
rect 112 284818 146 287194
rect -84 284725 84 284759
rect -84 284617 84 284651
rect -146 282182 -112 284558
rect 112 282182 146 284558
rect -84 282089 84 282123
rect -84 281981 84 282015
rect -146 279546 -112 281922
rect 112 279546 146 281922
rect -84 279453 84 279487
rect -84 279345 84 279379
rect -146 276910 -112 279286
rect 112 276910 146 279286
rect -84 276817 84 276851
rect -84 276709 84 276743
rect -146 274274 -112 276650
rect 112 274274 146 276650
rect -84 274181 84 274215
rect -84 274073 84 274107
rect -146 271638 -112 274014
rect 112 271638 146 274014
rect -84 271545 84 271579
rect -84 271437 84 271471
rect -146 269002 -112 271378
rect 112 269002 146 271378
rect -84 268909 84 268943
rect -84 268801 84 268835
rect -146 266366 -112 268742
rect 112 266366 146 268742
rect -84 266273 84 266307
rect -84 266165 84 266199
rect -146 263730 -112 266106
rect 112 263730 146 266106
rect -84 263637 84 263671
rect -84 263529 84 263563
rect -146 261094 -112 263470
rect 112 261094 146 263470
rect -84 261001 84 261035
rect -84 260893 84 260927
rect -146 258458 -112 260834
rect 112 258458 146 260834
rect -84 258365 84 258399
rect -84 258257 84 258291
rect -146 255822 -112 258198
rect 112 255822 146 258198
rect -84 255729 84 255763
rect -84 255621 84 255655
rect -146 253186 -112 255562
rect 112 253186 146 255562
rect -84 253093 84 253127
rect -84 252985 84 253019
rect -146 250550 -112 252926
rect 112 250550 146 252926
rect -84 250457 84 250491
rect -84 250349 84 250383
rect -146 247914 -112 250290
rect 112 247914 146 250290
rect -84 247821 84 247855
rect -84 247713 84 247747
rect -146 245278 -112 247654
rect 112 245278 146 247654
rect -84 245185 84 245219
rect -84 245077 84 245111
rect -146 242642 -112 245018
rect 112 242642 146 245018
rect -84 242549 84 242583
rect -84 242441 84 242475
rect -146 240006 -112 242382
rect 112 240006 146 242382
rect -84 239913 84 239947
rect -84 239805 84 239839
rect -146 237370 -112 239746
rect 112 237370 146 239746
rect -84 237277 84 237311
rect -84 237169 84 237203
rect -146 234734 -112 237110
rect 112 234734 146 237110
rect -84 234641 84 234675
rect -84 234533 84 234567
rect -146 232098 -112 234474
rect 112 232098 146 234474
rect -84 232005 84 232039
rect -84 231897 84 231931
rect -146 229462 -112 231838
rect 112 229462 146 231838
rect -84 229369 84 229403
rect -84 229261 84 229295
rect -146 226826 -112 229202
rect 112 226826 146 229202
rect -84 226733 84 226767
rect -84 226625 84 226659
rect -146 224190 -112 226566
rect 112 224190 146 226566
rect -84 224097 84 224131
rect -84 223989 84 224023
rect -146 221554 -112 223930
rect 112 221554 146 223930
rect -84 221461 84 221495
rect -84 221353 84 221387
rect -146 218918 -112 221294
rect 112 218918 146 221294
rect -84 218825 84 218859
rect -84 218717 84 218751
rect -146 216282 -112 218658
rect 112 216282 146 218658
rect -84 216189 84 216223
rect -84 216081 84 216115
rect -146 213646 -112 216022
rect 112 213646 146 216022
rect -84 213553 84 213587
rect -84 213445 84 213479
rect -146 211010 -112 213386
rect 112 211010 146 213386
rect -84 210917 84 210951
rect -84 210809 84 210843
rect -146 208374 -112 210750
rect 112 208374 146 210750
rect -84 208281 84 208315
rect -84 208173 84 208207
rect -146 205738 -112 208114
rect 112 205738 146 208114
rect -84 205645 84 205679
rect -84 205537 84 205571
rect -146 203102 -112 205478
rect 112 203102 146 205478
rect -84 203009 84 203043
rect -84 202901 84 202935
rect -146 200466 -112 202842
rect 112 200466 146 202842
rect -84 200373 84 200407
rect -84 200265 84 200299
rect -146 197830 -112 200206
rect 112 197830 146 200206
rect -84 197737 84 197771
rect -84 197629 84 197663
rect -146 195194 -112 197570
rect 112 195194 146 197570
rect -84 195101 84 195135
rect -84 194993 84 195027
rect -146 192558 -112 194934
rect 112 192558 146 194934
rect -84 192465 84 192499
rect -84 192357 84 192391
rect -146 189922 -112 192298
rect 112 189922 146 192298
rect -84 189829 84 189863
rect -84 189721 84 189755
rect -146 187286 -112 189662
rect 112 187286 146 189662
rect -84 187193 84 187227
rect -84 187085 84 187119
rect -146 184650 -112 187026
rect 112 184650 146 187026
rect -84 184557 84 184591
rect -84 184449 84 184483
rect -146 182014 -112 184390
rect 112 182014 146 184390
rect -84 181921 84 181955
rect -84 181813 84 181847
rect -146 179378 -112 181754
rect 112 179378 146 181754
rect -84 179285 84 179319
rect -84 179177 84 179211
rect -146 176742 -112 179118
rect 112 176742 146 179118
rect -84 176649 84 176683
rect -84 176541 84 176575
rect -146 174106 -112 176482
rect 112 174106 146 176482
rect -84 174013 84 174047
rect -84 173905 84 173939
rect -146 171470 -112 173846
rect 112 171470 146 173846
rect -84 171377 84 171411
rect -84 171269 84 171303
rect -146 168834 -112 171210
rect 112 168834 146 171210
rect -84 168741 84 168775
rect -84 168633 84 168667
rect -146 166198 -112 168574
rect 112 166198 146 168574
rect -84 166105 84 166139
rect -84 165997 84 166031
rect -146 163562 -112 165938
rect 112 163562 146 165938
rect -84 163469 84 163503
rect -84 163361 84 163395
rect -146 160926 -112 163302
rect 112 160926 146 163302
rect -84 160833 84 160867
rect -84 160725 84 160759
rect -146 158290 -112 160666
rect 112 158290 146 160666
rect -84 158197 84 158231
rect -84 158089 84 158123
rect -146 155654 -112 158030
rect 112 155654 146 158030
rect -84 155561 84 155595
rect -84 155453 84 155487
rect -146 153018 -112 155394
rect 112 153018 146 155394
rect -84 152925 84 152959
rect -84 152817 84 152851
rect -146 150382 -112 152758
rect 112 150382 146 152758
rect -84 150289 84 150323
rect -84 150181 84 150215
rect -146 147746 -112 150122
rect 112 147746 146 150122
rect -84 147653 84 147687
rect -84 147545 84 147579
rect -146 145110 -112 147486
rect 112 145110 146 147486
rect -84 145017 84 145051
rect -84 144909 84 144943
rect -146 142474 -112 144850
rect 112 142474 146 144850
rect -84 142381 84 142415
rect -84 142273 84 142307
rect -146 139838 -112 142214
rect 112 139838 146 142214
rect -84 139745 84 139779
rect -84 139637 84 139671
rect -146 137202 -112 139578
rect 112 137202 146 139578
rect -84 137109 84 137143
rect -84 137001 84 137035
rect -146 134566 -112 136942
rect 112 134566 146 136942
rect -84 134473 84 134507
rect -84 134365 84 134399
rect -146 131930 -112 134306
rect 112 131930 146 134306
rect -84 131837 84 131871
rect -84 131729 84 131763
rect -146 129294 -112 131670
rect 112 129294 146 131670
rect -84 129201 84 129235
rect -84 129093 84 129127
rect -146 126658 -112 129034
rect 112 126658 146 129034
rect -84 126565 84 126599
rect -84 126457 84 126491
rect -146 124022 -112 126398
rect 112 124022 146 126398
rect -84 123929 84 123963
rect -84 123821 84 123855
rect -146 121386 -112 123762
rect 112 121386 146 123762
rect -84 121293 84 121327
rect -84 121185 84 121219
rect -146 118750 -112 121126
rect 112 118750 146 121126
rect -84 118657 84 118691
rect -84 118549 84 118583
rect -146 116114 -112 118490
rect 112 116114 146 118490
rect -84 116021 84 116055
rect -84 115913 84 115947
rect -146 113478 -112 115854
rect 112 113478 146 115854
rect -84 113385 84 113419
rect -84 113277 84 113311
rect -146 110842 -112 113218
rect 112 110842 146 113218
rect -84 110749 84 110783
rect -84 110641 84 110675
rect -146 108206 -112 110582
rect 112 108206 146 110582
rect -84 108113 84 108147
rect -84 108005 84 108039
rect -146 105570 -112 107946
rect 112 105570 146 107946
rect -84 105477 84 105511
rect -84 105369 84 105403
rect -146 102934 -112 105310
rect 112 102934 146 105310
rect -84 102841 84 102875
rect -84 102733 84 102767
rect -146 100298 -112 102674
rect 112 100298 146 102674
rect -84 100205 84 100239
rect -84 100097 84 100131
rect -146 97662 -112 100038
rect 112 97662 146 100038
rect -84 97569 84 97603
rect -84 97461 84 97495
rect -146 95026 -112 97402
rect 112 95026 146 97402
rect -84 94933 84 94967
rect -84 94825 84 94859
rect -146 92390 -112 94766
rect 112 92390 146 94766
rect -84 92297 84 92331
rect -84 92189 84 92223
rect -146 89754 -112 92130
rect 112 89754 146 92130
rect -84 89661 84 89695
rect -84 89553 84 89587
rect -146 87118 -112 89494
rect 112 87118 146 89494
rect -84 87025 84 87059
rect -84 86917 84 86951
rect -146 84482 -112 86858
rect 112 84482 146 86858
rect -84 84389 84 84423
rect -84 84281 84 84315
rect -146 81846 -112 84222
rect 112 81846 146 84222
rect -84 81753 84 81787
rect -84 81645 84 81679
rect -146 79210 -112 81586
rect 112 79210 146 81586
rect -84 79117 84 79151
rect -84 79009 84 79043
rect -146 76574 -112 78950
rect 112 76574 146 78950
rect -84 76481 84 76515
rect -84 76373 84 76407
rect -146 73938 -112 76314
rect 112 73938 146 76314
rect -84 73845 84 73879
rect -84 73737 84 73771
rect -146 71302 -112 73678
rect 112 71302 146 73678
rect -84 71209 84 71243
rect -84 71101 84 71135
rect -146 68666 -112 71042
rect 112 68666 146 71042
rect -84 68573 84 68607
rect -84 68465 84 68499
rect -146 66030 -112 68406
rect 112 66030 146 68406
rect -84 65937 84 65971
rect -84 65829 84 65863
rect -146 63394 -112 65770
rect 112 63394 146 65770
rect -84 63301 84 63335
rect -84 63193 84 63227
rect -146 60758 -112 63134
rect 112 60758 146 63134
rect -84 60665 84 60699
rect -84 60557 84 60591
rect -146 58122 -112 60498
rect 112 58122 146 60498
rect -84 58029 84 58063
rect -84 57921 84 57955
rect -146 55486 -112 57862
rect 112 55486 146 57862
rect -84 55393 84 55427
rect -84 55285 84 55319
rect -146 52850 -112 55226
rect 112 52850 146 55226
rect -84 52757 84 52791
rect -84 52649 84 52683
rect -146 50214 -112 52590
rect 112 50214 146 52590
rect -84 50121 84 50155
rect -84 50013 84 50047
rect -146 47578 -112 49954
rect 112 47578 146 49954
rect -84 47485 84 47519
rect -84 47377 84 47411
rect -146 44942 -112 47318
rect 112 44942 146 47318
rect -84 44849 84 44883
rect -84 44741 84 44775
rect -146 42306 -112 44682
rect 112 42306 146 44682
rect -84 42213 84 42247
rect -84 42105 84 42139
rect -146 39670 -112 42046
rect 112 39670 146 42046
rect -84 39577 84 39611
rect -84 39469 84 39503
rect -146 37034 -112 39410
rect 112 37034 146 39410
rect -84 36941 84 36975
rect -84 36833 84 36867
rect -146 34398 -112 36774
rect 112 34398 146 36774
rect -84 34305 84 34339
rect -84 34197 84 34231
rect -146 31762 -112 34138
rect 112 31762 146 34138
rect -84 31669 84 31703
rect -84 31561 84 31595
rect -146 29126 -112 31502
rect 112 29126 146 31502
rect -84 29033 84 29067
rect -84 28925 84 28959
rect -146 26490 -112 28866
rect 112 26490 146 28866
rect -84 26397 84 26431
rect -84 26289 84 26323
rect -146 23854 -112 26230
rect 112 23854 146 26230
rect -84 23761 84 23795
rect -84 23653 84 23687
rect -146 21218 -112 23594
rect 112 21218 146 23594
rect -84 21125 84 21159
rect -84 21017 84 21051
rect -146 18582 -112 20958
rect 112 18582 146 20958
rect -84 18489 84 18523
rect -84 18381 84 18415
rect -146 15946 -112 18322
rect 112 15946 146 18322
rect -84 15853 84 15887
rect -84 15745 84 15779
rect -146 13310 -112 15686
rect 112 13310 146 15686
rect -84 13217 84 13251
rect -84 13109 84 13143
rect -146 10674 -112 13050
rect 112 10674 146 13050
rect -84 10581 84 10615
rect -84 10473 84 10507
rect -146 8038 -112 10414
rect 112 8038 146 10414
rect -84 7945 84 7979
rect -84 7837 84 7871
rect -146 5402 -112 7778
rect 112 5402 146 7778
rect -84 5309 84 5343
rect -84 5201 84 5235
rect -146 2766 -112 5142
rect 112 2766 146 5142
rect -84 2673 84 2707
rect -84 2565 84 2599
rect -146 130 -112 2506
rect 112 130 146 2506
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -2506 -112 -130
rect 112 -2506 146 -130
rect -84 -2599 84 -2565
rect -84 -2707 84 -2673
rect -146 -5142 -112 -2766
rect 112 -5142 146 -2766
rect -84 -5235 84 -5201
rect -84 -5343 84 -5309
rect -146 -7778 -112 -5402
rect 112 -7778 146 -5402
rect -84 -7871 84 -7837
rect -84 -7979 84 -7945
rect -146 -10414 -112 -8038
rect 112 -10414 146 -8038
rect -84 -10507 84 -10473
rect -84 -10615 84 -10581
rect -146 -13050 -112 -10674
rect 112 -13050 146 -10674
rect -84 -13143 84 -13109
rect -84 -13251 84 -13217
rect -146 -15686 -112 -13310
rect 112 -15686 146 -13310
rect -84 -15779 84 -15745
rect -84 -15887 84 -15853
rect -146 -18322 -112 -15946
rect 112 -18322 146 -15946
rect -84 -18415 84 -18381
rect -84 -18523 84 -18489
rect -146 -20958 -112 -18582
rect 112 -20958 146 -18582
rect -84 -21051 84 -21017
rect -84 -21159 84 -21125
rect -146 -23594 -112 -21218
rect 112 -23594 146 -21218
rect -84 -23687 84 -23653
rect -84 -23795 84 -23761
rect -146 -26230 -112 -23854
rect 112 -26230 146 -23854
rect -84 -26323 84 -26289
rect -84 -26431 84 -26397
rect -146 -28866 -112 -26490
rect 112 -28866 146 -26490
rect -84 -28959 84 -28925
rect -84 -29067 84 -29033
rect -146 -31502 -112 -29126
rect 112 -31502 146 -29126
rect -84 -31595 84 -31561
rect -84 -31703 84 -31669
rect -146 -34138 -112 -31762
rect 112 -34138 146 -31762
rect -84 -34231 84 -34197
rect -84 -34339 84 -34305
rect -146 -36774 -112 -34398
rect 112 -36774 146 -34398
rect -84 -36867 84 -36833
rect -84 -36975 84 -36941
rect -146 -39410 -112 -37034
rect 112 -39410 146 -37034
rect -84 -39503 84 -39469
rect -84 -39611 84 -39577
rect -146 -42046 -112 -39670
rect 112 -42046 146 -39670
rect -84 -42139 84 -42105
rect -84 -42247 84 -42213
rect -146 -44682 -112 -42306
rect 112 -44682 146 -42306
rect -84 -44775 84 -44741
rect -84 -44883 84 -44849
rect -146 -47318 -112 -44942
rect 112 -47318 146 -44942
rect -84 -47411 84 -47377
rect -84 -47519 84 -47485
rect -146 -49954 -112 -47578
rect 112 -49954 146 -47578
rect -84 -50047 84 -50013
rect -84 -50155 84 -50121
rect -146 -52590 -112 -50214
rect 112 -52590 146 -50214
rect -84 -52683 84 -52649
rect -84 -52791 84 -52757
rect -146 -55226 -112 -52850
rect 112 -55226 146 -52850
rect -84 -55319 84 -55285
rect -84 -55427 84 -55393
rect -146 -57862 -112 -55486
rect 112 -57862 146 -55486
rect -84 -57955 84 -57921
rect -84 -58063 84 -58029
rect -146 -60498 -112 -58122
rect 112 -60498 146 -58122
rect -84 -60591 84 -60557
rect -84 -60699 84 -60665
rect -146 -63134 -112 -60758
rect 112 -63134 146 -60758
rect -84 -63227 84 -63193
rect -84 -63335 84 -63301
rect -146 -65770 -112 -63394
rect 112 -65770 146 -63394
rect -84 -65863 84 -65829
rect -84 -65971 84 -65937
rect -146 -68406 -112 -66030
rect 112 -68406 146 -66030
rect -84 -68499 84 -68465
rect -84 -68607 84 -68573
rect -146 -71042 -112 -68666
rect 112 -71042 146 -68666
rect -84 -71135 84 -71101
rect -84 -71243 84 -71209
rect -146 -73678 -112 -71302
rect 112 -73678 146 -71302
rect -84 -73771 84 -73737
rect -84 -73879 84 -73845
rect -146 -76314 -112 -73938
rect 112 -76314 146 -73938
rect -84 -76407 84 -76373
rect -84 -76515 84 -76481
rect -146 -78950 -112 -76574
rect 112 -78950 146 -76574
rect -84 -79043 84 -79009
rect -84 -79151 84 -79117
rect -146 -81586 -112 -79210
rect 112 -81586 146 -79210
rect -84 -81679 84 -81645
rect -84 -81787 84 -81753
rect -146 -84222 -112 -81846
rect 112 -84222 146 -81846
rect -84 -84315 84 -84281
rect -84 -84423 84 -84389
rect -146 -86858 -112 -84482
rect 112 -86858 146 -84482
rect -84 -86951 84 -86917
rect -84 -87059 84 -87025
rect -146 -89494 -112 -87118
rect 112 -89494 146 -87118
rect -84 -89587 84 -89553
rect -84 -89695 84 -89661
rect -146 -92130 -112 -89754
rect 112 -92130 146 -89754
rect -84 -92223 84 -92189
rect -84 -92331 84 -92297
rect -146 -94766 -112 -92390
rect 112 -94766 146 -92390
rect -84 -94859 84 -94825
rect -84 -94967 84 -94933
rect -146 -97402 -112 -95026
rect 112 -97402 146 -95026
rect -84 -97495 84 -97461
rect -84 -97603 84 -97569
rect -146 -100038 -112 -97662
rect 112 -100038 146 -97662
rect -84 -100131 84 -100097
rect -84 -100239 84 -100205
rect -146 -102674 -112 -100298
rect 112 -102674 146 -100298
rect -84 -102767 84 -102733
rect -84 -102875 84 -102841
rect -146 -105310 -112 -102934
rect 112 -105310 146 -102934
rect -84 -105403 84 -105369
rect -84 -105511 84 -105477
rect -146 -107946 -112 -105570
rect 112 -107946 146 -105570
rect -84 -108039 84 -108005
rect -84 -108147 84 -108113
rect -146 -110582 -112 -108206
rect 112 -110582 146 -108206
rect -84 -110675 84 -110641
rect -84 -110783 84 -110749
rect -146 -113218 -112 -110842
rect 112 -113218 146 -110842
rect -84 -113311 84 -113277
rect -84 -113419 84 -113385
rect -146 -115854 -112 -113478
rect 112 -115854 146 -113478
rect -84 -115947 84 -115913
rect -84 -116055 84 -116021
rect -146 -118490 -112 -116114
rect 112 -118490 146 -116114
rect -84 -118583 84 -118549
rect -84 -118691 84 -118657
rect -146 -121126 -112 -118750
rect 112 -121126 146 -118750
rect -84 -121219 84 -121185
rect -84 -121327 84 -121293
rect -146 -123762 -112 -121386
rect 112 -123762 146 -121386
rect -84 -123855 84 -123821
rect -84 -123963 84 -123929
rect -146 -126398 -112 -124022
rect 112 -126398 146 -124022
rect -84 -126491 84 -126457
rect -84 -126599 84 -126565
rect -146 -129034 -112 -126658
rect 112 -129034 146 -126658
rect -84 -129127 84 -129093
rect -84 -129235 84 -129201
rect -146 -131670 -112 -129294
rect 112 -131670 146 -129294
rect -84 -131763 84 -131729
rect -84 -131871 84 -131837
rect -146 -134306 -112 -131930
rect 112 -134306 146 -131930
rect -84 -134399 84 -134365
rect -84 -134507 84 -134473
rect -146 -136942 -112 -134566
rect 112 -136942 146 -134566
rect -84 -137035 84 -137001
rect -84 -137143 84 -137109
rect -146 -139578 -112 -137202
rect 112 -139578 146 -137202
rect -84 -139671 84 -139637
rect -84 -139779 84 -139745
rect -146 -142214 -112 -139838
rect 112 -142214 146 -139838
rect -84 -142307 84 -142273
rect -84 -142415 84 -142381
rect -146 -144850 -112 -142474
rect 112 -144850 146 -142474
rect -84 -144943 84 -144909
rect -84 -145051 84 -145017
rect -146 -147486 -112 -145110
rect 112 -147486 146 -145110
rect -84 -147579 84 -147545
rect -84 -147687 84 -147653
rect -146 -150122 -112 -147746
rect 112 -150122 146 -147746
rect -84 -150215 84 -150181
rect -84 -150323 84 -150289
rect -146 -152758 -112 -150382
rect 112 -152758 146 -150382
rect -84 -152851 84 -152817
rect -84 -152959 84 -152925
rect -146 -155394 -112 -153018
rect 112 -155394 146 -153018
rect -84 -155487 84 -155453
rect -84 -155595 84 -155561
rect -146 -158030 -112 -155654
rect 112 -158030 146 -155654
rect -84 -158123 84 -158089
rect -84 -158231 84 -158197
rect -146 -160666 -112 -158290
rect 112 -160666 146 -158290
rect -84 -160759 84 -160725
rect -84 -160867 84 -160833
rect -146 -163302 -112 -160926
rect 112 -163302 146 -160926
rect -84 -163395 84 -163361
rect -84 -163503 84 -163469
rect -146 -165938 -112 -163562
rect 112 -165938 146 -163562
rect -84 -166031 84 -165997
rect -84 -166139 84 -166105
rect -146 -168574 -112 -166198
rect 112 -168574 146 -166198
rect -84 -168667 84 -168633
rect -84 -168775 84 -168741
rect -146 -171210 -112 -168834
rect 112 -171210 146 -168834
rect -84 -171303 84 -171269
rect -84 -171411 84 -171377
rect -146 -173846 -112 -171470
rect 112 -173846 146 -171470
rect -84 -173939 84 -173905
rect -84 -174047 84 -174013
rect -146 -176482 -112 -174106
rect 112 -176482 146 -174106
rect -84 -176575 84 -176541
rect -84 -176683 84 -176649
rect -146 -179118 -112 -176742
rect 112 -179118 146 -176742
rect -84 -179211 84 -179177
rect -84 -179319 84 -179285
rect -146 -181754 -112 -179378
rect 112 -181754 146 -179378
rect -84 -181847 84 -181813
rect -84 -181955 84 -181921
rect -146 -184390 -112 -182014
rect 112 -184390 146 -182014
rect -84 -184483 84 -184449
rect -84 -184591 84 -184557
rect -146 -187026 -112 -184650
rect 112 -187026 146 -184650
rect -84 -187119 84 -187085
rect -84 -187227 84 -187193
rect -146 -189662 -112 -187286
rect 112 -189662 146 -187286
rect -84 -189755 84 -189721
rect -84 -189863 84 -189829
rect -146 -192298 -112 -189922
rect 112 -192298 146 -189922
rect -84 -192391 84 -192357
rect -84 -192499 84 -192465
rect -146 -194934 -112 -192558
rect 112 -194934 146 -192558
rect -84 -195027 84 -194993
rect -84 -195135 84 -195101
rect -146 -197570 -112 -195194
rect 112 -197570 146 -195194
rect -84 -197663 84 -197629
rect -84 -197771 84 -197737
rect -146 -200206 -112 -197830
rect 112 -200206 146 -197830
rect -84 -200299 84 -200265
rect -84 -200407 84 -200373
rect -146 -202842 -112 -200466
rect 112 -202842 146 -200466
rect -84 -202935 84 -202901
rect -84 -203043 84 -203009
rect -146 -205478 -112 -203102
rect 112 -205478 146 -203102
rect -84 -205571 84 -205537
rect -84 -205679 84 -205645
rect -146 -208114 -112 -205738
rect 112 -208114 146 -205738
rect -84 -208207 84 -208173
rect -84 -208315 84 -208281
rect -146 -210750 -112 -208374
rect 112 -210750 146 -208374
rect -84 -210843 84 -210809
rect -84 -210951 84 -210917
rect -146 -213386 -112 -211010
rect 112 -213386 146 -211010
rect -84 -213479 84 -213445
rect -84 -213587 84 -213553
rect -146 -216022 -112 -213646
rect 112 -216022 146 -213646
rect -84 -216115 84 -216081
rect -84 -216223 84 -216189
rect -146 -218658 -112 -216282
rect 112 -218658 146 -216282
rect -84 -218751 84 -218717
rect -84 -218859 84 -218825
rect -146 -221294 -112 -218918
rect 112 -221294 146 -218918
rect -84 -221387 84 -221353
rect -84 -221495 84 -221461
rect -146 -223930 -112 -221554
rect 112 -223930 146 -221554
rect -84 -224023 84 -223989
rect -84 -224131 84 -224097
rect -146 -226566 -112 -224190
rect 112 -226566 146 -224190
rect -84 -226659 84 -226625
rect -84 -226767 84 -226733
rect -146 -229202 -112 -226826
rect 112 -229202 146 -226826
rect -84 -229295 84 -229261
rect -84 -229403 84 -229369
rect -146 -231838 -112 -229462
rect 112 -231838 146 -229462
rect -84 -231931 84 -231897
rect -84 -232039 84 -232005
rect -146 -234474 -112 -232098
rect 112 -234474 146 -232098
rect -84 -234567 84 -234533
rect -84 -234675 84 -234641
rect -146 -237110 -112 -234734
rect 112 -237110 146 -234734
rect -84 -237203 84 -237169
rect -84 -237311 84 -237277
rect -146 -239746 -112 -237370
rect 112 -239746 146 -237370
rect -84 -239839 84 -239805
rect -84 -239947 84 -239913
rect -146 -242382 -112 -240006
rect 112 -242382 146 -240006
rect -84 -242475 84 -242441
rect -84 -242583 84 -242549
rect -146 -245018 -112 -242642
rect 112 -245018 146 -242642
rect -84 -245111 84 -245077
rect -84 -245219 84 -245185
rect -146 -247654 -112 -245278
rect 112 -247654 146 -245278
rect -84 -247747 84 -247713
rect -84 -247855 84 -247821
rect -146 -250290 -112 -247914
rect 112 -250290 146 -247914
rect -84 -250383 84 -250349
rect -84 -250491 84 -250457
rect -146 -252926 -112 -250550
rect 112 -252926 146 -250550
rect -84 -253019 84 -252985
rect -84 -253127 84 -253093
rect -146 -255562 -112 -253186
rect 112 -255562 146 -253186
rect -84 -255655 84 -255621
rect -84 -255763 84 -255729
rect -146 -258198 -112 -255822
rect 112 -258198 146 -255822
rect -84 -258291 84 -258257
rect -84 -258399 84 -258365
rect -146 -260834 -112 -258458
rect 112 -260834 146 -258458
rect -84 -260927 84 -260893
rect -84 -261035 84 -261001
rect -146 -263470 -112 -261094
rect 112 -263470 146 -261094
rect -84 -263563 84 -263529
rect -84 -263671 84 -263637
rect -146 -266106 -112 -263730
rect 112 -266106 146 -263730
rect -84 -266199 84 -266165
rect -84 -266307 84 -266273
rect -146 -268742 -112 -266366
rect 112 -268742 146 -266366
rect -84 -268835 84 -268801
rect -84 -268943 84 -268909
rect -146 -271378 -112 -269002
rect 112 -271378 146 -269002
rect -84 -271471 84 -271437
rect -84 -271579 84 -271545
rect -146 -274014 -112 -271638
rect 112 -274014 146 -271638
rect -84 -274107 84 -274073
rect -84 -274215 84 -274181
rect -146 -276650 -112 -274274
rect 112 -276650 146 -274274
rect -84 -276743 84 -276709
rect -84 -276851 84 -276817
rect -146 -279286 -112 -276910
rect 112 -279286 146 -276910
rect -84 -279379 84 -279345
rect -84 -279487 84 -279453
rect -146 -281922 -112 -279546
rect 112 -281922 146 -279546
rect -84 -282015 84 -281981
rect -84 -282123 84 -282089
rect -146 -284558 -112 -282182
rect 112 -284558 146 -282182
rect -84 -284651 84 -284617
rect -84 -284759 84 -284725
rect -146 -287194 -112 -284818
rect 112 -287194 146 -284818
rect -84 -287287 84 -287253
rect -84 -287395 84 -287361
rect -146 -289830 -112 -287454
rect 112 -289830 146 -287454
rect -84 -289923 84 -289889
rect -84 -290031 84 -289997
rect -146 -292466 -112 -290090
rect 112 -292466 146 -290090
rect -84 -292559 84 -292525
rect -84 -292667 84 -292633
rect -146 -295102 -112 -292726
rect 112 -295102 146 -292726
rect -84 -295195 84 -295161
rect -84 -295303 84 -295269
rect -146 -297738 -112 -295362
rect 112 -297738 146 -295362
rect -84 -297831 84 -297797
rect -84 -297939 84 -297905
rect -146 -300374 -112 -297998
rect 112 -300374 146 -297998
rect -84 -300467 84 -300433
rect -84 -300575 84 -300541
rect -146 -303010 -112 -300634
rect 112 -303010 146 -300634
rect -84 -303103 84 -303069
rect -84 -303211 84 -303177
rect -146 -305646 -112 -303270
rect 112 -305646 146 -303270
rect -84 -305739 84 -305705
rect -84 -305847 84 -305813
rect -146 -308282 -112 -305906
rect 112 -308282 146 -305906
rect -84 -308375 84 -308341
rect -84 -308483 84 -308449
rect -146 -310918 -112 -308542
rect 112 -310918 146 -308542
rect -84 -311011 84 -310977
rect -84 -311119 84 -311085
rect -146 -313554 -112 -311178
rect 112 -313554 146 -311178
rect -84 -313647 84 -313613
rect -84 -313755 84 -313721
rect -146 -316190 -112 -313814
rect 112 -316190 146 -313814
rect -84 -316283 84 -316249
rect -84 -316391 84 -316357
rect -146 -318826 -112 -316450
rect 112 -318826 146 -316450
rect -84 -318919 84 -318885
rect -84 -319027 84 -318993
rect -146 -321462 -112 -319086
rect 112 -321462 146 -319086
rect -84 -321555 84 -321521
rect -84 -321663 84 -321629
rect -146 -324098 -112 -321722
rect 112 -324098 146 -321722
rect -84 -324191 84 -324157
rect -84 -324299 84 -324265
rect -146 -326734 -112 -324358
rect 112 -326734 146 -324358
rect -84 -326827 84 -326793
rect -84 -326935 84 -326901
rect -146 -329370 -112 -326994
rect 112 -329370 146 -326994
rect -84 -329463 84 -329429
rect -84 -329571 84 -329537
rect -146 -332006 -112 -329630
rect 112 -332006 146 -329630
rect -84 -332099 84 -332065
rect -84 -332207 84 -332173
rect -146 -334642 -112 -332266
rect 112 -334642 146 -332266
rect -84 -334735 84 -334701
rect -84 -334843 84 -334809
rect -146 -337278 -112 -334902
rect 112 -337278 146 -334902
rect -84 -337371 84 -337337
<< metal1 >>
rect -96 337371 96 337377
rect -96 337337 -84 337371
rect 84 337337 96 337371
rect -96 337331 96 337337
rect -152 337278 -106 337290
rect -152 334902 -146 337278
rect -112 334902 -106 337278
rect -152 334890 -106 334902
rect 106 337278 152 337290
rect 106 334902 112 337278
rect 146 334902 152 337278
rect 106 334890 152 334902
rect -96 334843 96 334849
rect -96 334809 -84 334843
rect 84 334809 96 334843
rect -96 334803 96 334809
rect -96 334735 96 334741
rect -96 334701 -84 334735
rect 84 334701 96 334735
rect -96 334695 96 334701
rect -152 334642 -106 334654
rect -152 332266 -146 334642
rect -112 332266 -106 334642
rect -152 332254 -106 332266
rect 106 334642 152 334654
rect 106 332266 112 334642
rect 146 332266 152 334642
rect 106 332254 152 332266
rect -96 332207 96 332213
rect -96 332173 -84 332207
rect 84 332173 96 332207
rect -96 332167 96 332173
rect -96 332099 96 332105
rect -96 332065 -84 332099
rect 84 332065 96 332099
rect -96 332059 96 332065
rect -152 332006 -106 332018
rect -152 329630 -146 332006
rect -112 329630 -106 332006
rect -152 329618 -106 329630
rect 106 332006 152 332018
rect 106 329630 112 332006
rect 146 329630 152 332006
rect 106 329618 152 329630
rect -96 329571 96 329577
rect -96 329537 -84 329571
rect 84 329537 96 329571
rect -96 329531 96 329537
rect -96 329463 96 329469
rect -96 329429 -84 329463
rect 84 329429 96 329463
rect -96 329423 96 329429
rect -152 329370 -106 329382
rect -152 326994 -146 329370
rect -112 326994 -106 329370
rect -152 326982 -106 326994
rect 106 329370 152 329382
rect 106 326994 112 329370
rect 146 326994 152 329370
rect 106 326982 152 326994
rect -96 326935 96 326941
rect -96 326901 -84 326935
rect 84 326901 96 326935
rect -96 326895 96 326901
rect -96 326827 96 326833
rect -96 326793 -84 326827
rect 84 326793 96 326827
rect -96 326787 96 326793
rect -152 326734 -106 326746
rect -152 324358 -146 326734
rect -112 324358 -106 326734
rect -152 324346 -106 324358
rect 106 326734 152 326746
rect 106 324358 112 326734
rect 146 324358 152 326734
rect 106 324346 152 324358
rect -96 324299 96 324305
rect -96 324265 -84 324299
rect 84 324265 96 324299
rect -96 324259 96 324265
rect -96 324191 96 324197
rect -96 324157 -84 324191
rect 84 324157 96 324191
rect -96 324151 96 324157
rect -152 324098 -106 324110
rect -152 321722 -146 324098
rect -112 321722 -106 324098
rect -152 321710 -106 321722
rect 106 324098 152 324110
rect 106 321722 112 324098
rect 146 321722 152 324098
rect 106 321710 152 321722
rect -96 321663 96 321669
rect -96 321629 -84 321663
rect 84 321629 96 321663
rect -96 321623 96 321629
rect -96 321555 96 321561
rect -96 321521 -84 321555
rect 84 321521 96 321555
rect -96 321515 96 321521
rect -152 321462 -106 321474
rect -152 319086 -146 321462
rect -112 319086 -106 321462
rect -152 319074 -106 319086
rect 106 321462 152 321474
rect 106 319086 112 321462
rect 146 319086 152 321462
rect 106 319074 152 319086
rect -96 319027 96 319033
rect -96 318993 -84 319027
rect 84 318993 96 319027
rect -96 318987 96 318993
rect -96 318919 96 318925
rect -96 318885 -84 318919
rect 84 318885 96 318919
rect -96 318879 96 318885
rect -152 318826 -106 318838
rect -152 316450 -146 318826
rect -112 316450 -106 318826
rect -152 316438 -106 316450
rect 106 318826 152 318838
rect 106 316450 112 318826
rect 146 316450 152 318826
rect 106 316438 152 316450
rect -96 316391 96 316397
rect -96 316357 -84 316391
rect 84 316357 96 316391
rect -96 316351 96 316357
rect -96 316283 96 316289
rect -96 316249 -84 316283
rect 84 316249 96 316283
rect -96 316243 96 316249
rect -152 316190 -106 316202
rect -152 313814 -146 316190
rect -112 313814 -106 316190
rect -152 313802 -106 313814
rect 106 316190 152 316202
rect 106 313814 112 316190
rect 146 313814 152 316190
rect 106 313802 152 313814
rect -96 313755 96 313761
rect -96 313721 -84 313755
rect 84 313721 96 313755
rect -96 313715 96 313721
rect -96 313647 96 313653
rect -96 313613 -84 313647
rect 84 313613 96 313647
rect -96 313607 96 313613
rect -152 313554 -106 313566
rect -152 311178 -146 313554
rect -112 311178 -106 313554
rect -152 311166 -106 311178
rect 106 313554 152 313566
rect 106 311178 112 313554
rect 146 311178 152 313554
rect 106 311166 152 311178
rect -96 311119 96 311125
rect -96 311085 -84 311119
rect 84 311085 96 311119
rect -96 311079 96 311085
rect -96 311011 96 311017
rect -96 310977 -84 311011
rect 84 310977 96 311011
rect -96 310971 96 310977
rect -152 310918 -106 310930
rect -152 308542 -146 310918
rect -112 308542 -106 310918
rect -152 308530 -106 308542
rect 106 310918 152 310930
rect 106 308542 112 310918
rect 146 308542 152 310918
rect 106 308530 152 308542
rect -96 308483 96 308489
rect -96 308449 -84 308483
rect 84 308449 96 308483
rect -96 308443 96 308449
rect -96 308375 96 308381
rect -96 308341 -84 308375
rect 84 308341 96 308375
rect -96 308335 96 308341
rect -152 308282 -106 308294
rect -152 305906 -146 308282
rect -112 305906 -106 308282
rect -152 305894 -106 305906
rect 106 308282 152 308294
rect 106 305906 112 308282
rect 146 305906 152 308282
rect 106 305894 152 305906
rect -96 305847 96 305853
rect -96 305813 -84 305847
rect 84 305813 96 305847
rect -96 305807 96 305813
rect -96 305739 96 305745
rect -96 305705 -84 305739
rect 84 305705 96 305739
rect -96 305699 96 305705
rect -152 305646 -106 305658
rect -152 303270 -146 305646
rect -112 303270 -106 305646
rect -152 303258 -106 303270
rect 106 305646 152 305658
rect 106 303270 112 305646
rect 146 303270 152 305646
rect 106 303258 152 303270
rect -96 303211 96 303217
rect -96 303177 -84 303211
rect 84 303177 96 303211
rect -96 303171 96 303177
rect -96 303103 96 303109
rect -96 303069 -84 303103
rect 84 303069 96 303103
rect -96 303063 96 303069
rect -152 303010 -106 303022
rect -152 300634 -146 303010
rect -112 300634 -106 303010
rect -152 300622 -106 300634
rect 106 303010 152 303022
rect 106 300634 112 303010
rect 146 300634 152 303010
rect 106 300622 152 300634
rect -96 300575 96 300581
rect -96 300541 -84 300575
rect 84 300541 96 300575
rect -96 300535 96 300541
rect -96 300467 96 300473
rect -96 300433 -84 300467
rect 84 300433 96 300467
rect -96 300427 96 300433
rect -152 300374 -106 300386
rect -152 297998 -146 300374
rect -112 297998 -106 300374
rect -152 297986 -106 297998
rect 106 300374 152 300386
rect 106 297998 112 300374
rect 146 297998 152 300374
rect 106 297986 152 297998
rect -96 297939 96 297945
rect -96 297905 -84 297939
rect 84 297905 96 297939
rect -96 297899 96 297905
rect -96 297831 96 297837
rect -96 297797 -84 297831
rect 84 297797 96 297831
rect -96 297791 96 297797
rect -152 297738 -106 297750
rect -152 295362 -146 297738
rect -112 295362 -106 297738
rect -152 295350 -106 295362
rect 106 297738 152 297750
rect 106 295362 112 297738
rect 146 295362 152 297738
rect 106 295350 152 295362
rect -96 295303 96 295309
rect -96 295269 -84 295303
rect 84 295269 96 295303
rect -96 295263 96 295269
rect -96 295195 96 295201
rect -96 295161 -84 295195
rect 84 295161 96 295195
rect -96 295155 96 295161
rect -152 295102 -106 295114
rect -152 292726 -146 295102
rect -112 292726 -106 295102
rect -152 292714 -106 292726
rect 106 295102 152 295114
rect 106 292726 112 295102
rect 146 292726 152 295102
rect 106 292714 152 292726
rect -96 292667 96 292673
rect -96 292633 -84 292667
rect 84 292633 96 292667
rect -96 292627 96 292633
rect -96 292559 96 292565
rect -96 292525 -84 292559
rect 84 292525 96 292559
rect -96 292519 96 292525
rect -152 292466 -106 292478
rect -152 290090 -146 292466
rect -112 290090 -106 292466
rect -152 290078 -106 290090
rect 106 292466 152 292478
rect 106 290090 112 292466
rect 146 290090 152 292466
rect 106 290078 152 290090
rect -96 290031 96 290037
rect -96 289997 -84 290031
rect 84 289997 96 290031
rect -96 289991 96 289997
rect -96 289923 96 289929
rect -96 289889 -84 289923
rect 84 289889 96 289923
rect -96 289883 96 289889
rect -152 289830 -106 289842
rect -152 287454 -146 289830
rect -112 287454 -106 289830
rect -152 287442 -106 287454
rect 106 289830 152 289842
rect 106 287454 112 289830
rect 146 287454 152 289830
rect 106 287442 152 287454
rect -96 287395 96 287401
rect -96 287361 -84 287395
rect 84 287361 96 287395
rect -96 287355 96 287361
rect -96 287287 96 287293
rect -96 287253 -84 287287
rect 84 287253 96 287287
rect -96 287247 96 287253
rect -152 287194 -106 287206
rect -152 284818 -146 287194
rect -112 284818 -106 287194
rect -152 284806 -106 284818
rect 106 287194 152 287206
rect 106 284818 112 287194
rect 146 284818 152 287194
rect 106 284806 152 284818
rect -96 284759 96 284765
rect -96 284725 -84 284759
rect 84 284725 96 284759
rect -96 284719 96 284725
rect -96 284651 96 284657
rect -96 284617 -84 284651
rect 84 284617 96 284651
rect -96 284611 96 284617
rect -152 284558 -106 284570
rect -152 282182 -146 284558
rect -112 282182 -106 284558
rect -152 282170 -106 282182
rect 106 284558 152 284570
rect 106 282182 112 284558
rect 146 282182 152 284558
rect 106 282170 152 282182
rect -96 282123 96 282129
rect -96 282089 -84 282123
rect 84 282089 96 282123
rect -96 282083 96 282089
rect -96 282015 96 282021
rect -96 281981 -84 282015
rect 84 281981 96 282015
rect -96 281975 96 281981
rect -152 281922 -106 281934
rect -152 279546 -146 281922
rect -112 279546 -106 281922
rect -152 279534 -106 279546
rect 106 281922 152 281934
rect 106 279546 112 281922
rect 146 279546 152 281922
rect 106 279534 152 279546
rect -96 279487 96 279493
rect -96 279453 -84 279487
rect 84 279453 96 279487
rect -96 279447 96 279453
rect -96 279379 96 279385
rect -96 279345 -84 279379
rect 84 279345 96 279379
rect -96 279339 96 279345
rect -152 279286 -106 279298
rect -152 276910 -146 279286
rect -112 276910 -106 279286
rect -152 276898 -106 276910
rect 106 279286 152 279298
rect 106 276910 112 279286
rect 146 276910 152 279286
rect 106 276898 152 276910
rect -96 276851 96 276857
rect -96 276817 -84 276851
rect 84 276817 96 276851
rect -96 276811 96 276817
rect -96 276743 96 276749
rect -96 276709 -84 276743
rect 84 276709 96 276743
rect -96 276703 96 276709
rect -152 276650 -106 276662
rect -152 274274 -146 276650
rect -112 274274 -106 276650
rect -152 274262 -106 274274
rect 106 276650 152 276662
rect 106 274274 112 276650
rect 146 274274 152 276650
rect 106 274262 152 274274
rect -96 274215 96 274221
rect -96 274181 -84 274215
rect 84 274181 96 274215
rect -96 274175 96 274181
rect -96 274107 96 274113
rect -96 274073 -84 274107
rect 84 274073 96 274107
rect -96 274067 96 274073
rect -152 274014 -106 274026
rect -152 271638 -146 274014
rect -112 271638 -106 274014
rect -152 271626 -106 271638
rect 106 274014 152 274026
rect 106 271638 112 274014
rect 146 271638 152 274014
rect 106 271626 152 271638
rect -96 271579 96 271585
rect -96 271545 -84 271579
rect 84 271545 96 271579
rect -96 271539 96 271545
rect -96 271471 96 271477
rect -96 271437 -84 271471
rect 84 271437 96 271471
rect -96 271431 96 271437
rect -152 271378 -106 271390
rect -152 269002 -146 271378
rect -112 269002 -106 271378
rect -152 268990 -106 269002
rect 106 271378 152 271390
rect 106 269002 112 271378
rect 146 269002 152 271378
rect 106 268990 152 269002
rect -96 268943 96 268949
rect -96 268909 -84 268943
rect 84 268909 96 268943
rect -96 268903 96 268909
rect -96 268835 96 268841
rect -96 268801 -84 268835
rect 84 268801 96 268835
rect -96 268795 96 268801
rect -152 268742 -106 268754
rect -152 266366 -146 268742
rect -112 266366 -106 268742
rect -152 266354 -106 266366
rect 106 268742 152 268754
rect 106 266366 112 268742
rect 146 266366 152 268742
rect 106 266354 152 266366
rect -96 266307 96 266313
rect -96 266273 -84 266307
rect 84 266273 96 266307
rect -96 266267 96 266273
rect -96 266199 96 266205
rect -96 266165 -84 266199
rect 84 266165 96 266199
rect -96 266159 96 266165
rect -152 266106 -106 266118
rect -152 263730 -146 266106
rect -112 263730 -106 266106
rect -152 263718 -106 263730
rect 106 266106 152 266118
rect 106 263730 112 266106
rect 146 263730 152 266106
rect 106 263718 152 263730
rect -96 263671 96 263677
rect -96 263637 -84 263671
rect 84 263637 96 263671
rect -96 263631 96 263637
rect -96 263563 96 263569
rect -96 263529 -84 263563
rect 84 263529 96 263563
rect -96 263523 96 263529
rect -152 263470 -106 263482
rect -152 261094 -146 263470
rect -112 261094 -106 263470
rect -152 261082 -106 261094
rect 106 263470 152 263482
rect 106 261094 112 263470
rect 146 261094 152 263470
rect 106 261082 152 261094
rect -96 261035 96 261041
rect -96 261001 -84 261035
rect 84 261001 96 261035
rect -96 260995 96 261001
rect -96 260927 96 260933
rect -96 260893 -84 260927
rect 84 260893 96 260927
rect -96 260887 96 260893
rect -152 260834 -106 260846
rect -152 258458 -146 260834
rect -112 258458 -106 260834
rect -152 258446 -106 258458
rect 106 260834 152 260846
rect 106 258458 112 260834
rect 146 258458 152 260834
rect 106 258446 152 258458
rect -96 258399 96 258405
rect -96 258365 -84 258399
rect 84 258365 96 258399
rect -96 258359 96 258365
rect -96 258291 96 258297
rect -96 258257 -84 258291
rect 84 258257 96 258291
rect -96 258251 96 258257
rect -152 258198 -106 258210
rect -152 255822 -146 258198
rect -112 255822 -106 258198
rect -152 255810 -106 255822
rect 106 258198 152 258210
rect 106 255822 112 258198
rect 146 255822 152 258198
rect 106 255810 152 255822
rect -96 255763 96 255769
rect -96 255729 -84 255763
rect 84 255729 96 255763
rect -96 255723 96 255729
rect -96 255655 96 255661
rect -96 255621 -84 255655
rect 84 255621 96 255655
rect -96 255615 96 255621
rect -152 255562 -106 255574
rect -152 253186 -146 255562
rect -112 253186 -106 255562
rect -152 253174 -106 253186
rect 106 255562 152 255574
rect 106 253186 112 255562
rect 146 253186 152 255562
rect 106 253174 152 253186
rect -96 253127 96 253133
rect -96 253093 -84 253127
rect 84 253093 96 253127
rect -96 253087 96 253093
rect -96 253019 96 253025
rect -96 252985 -84 253019
rect 84 252985 96 253019
rect -96 252979 96 252985
rect -152 252926 -106 252938
rect -152 250550 -146 252926
rect -112 250550 -106 252926
rect -152 250538 -106 250550
rect 106 252926 152 252938
rect 106 250550 112 252926
rect 146 250550 152 252926
rect 106 250538 152 250550
rect -96 250491 96 250497
rect -96 250457 -84 250491
rect 84 250457 96 250491
rect -96 250451 96 250457
rect -96 250383 96 250389
rect -96 250349 -84 250383
rect 84 250349 96 250383
rect -96 250343 96 250349
rect -152 250290 -106 250302
rect -152 247914 -146 250290
rect -112 247914 -106 250290
rect -152 247902 -106 247914
rect 106 250290 152 250302
rect 106 247914 112 250290
rect 146 247914 152 250290
rect 106 247902 152 247914
rect -96 247855 96 247861
rect -96 247821 -84 247855
rect 84 247821 96 247855
rect -96 247815 96 247821
rect -96 247747 96 247753
rect -96 247713 -84 247747
rect 84 247713 96 247747
rect -96 247707 96 247713
rect -152 247654 -106 247666
rect -152 245278 -146 247654
rect -112 245278 -106 247654
rect -152 245266 -106 245278
rect 106 247654 152 247666
rect 106 245278 112 247654
rect 146 245278 152 247654
rect 106 245266 152 245278
rect -96 245219 96 245225
rect -96 245185 -84 245219
rect 84 245185 96 245219
rect -96 245179 96 245185
rect -96 245111 96 245117
rect -96 245077 -84 245111
rect 84 245077 96 245111
rect -96 245071 96 245077
rect -152 245018 -106 245030
rect -152 242642 -146 245018
rect -112 242642 -106 245018
rect -152 242630 -106 242642
rect 106 245018 152 245030
rect 106 242642 112 245018
rect 146 242642 152 245018
rect 106 242630 152 242642
rect -96 242583 96 242589
rect -96 242549 -84 242583
rect 84 242549 96 242583
rect -96 242543 96 242549
rect -96 242475 96 242481
rect -96 242441 -84 242475
rect 84 242441 96 242475
rect -96 242435 96 242441
rect -152 242382 -106 242394
rect -152 240006 -146 242382
rect -112 240006 -106 242382
rect -152 239994 -106 240006
rect 106 242382 152 242394
rect 106 240006 112 242382
rect 146 240006 152 242382
rect 106 239994 152 240006
rect -96 239947 96 239953
rect -96 239913 -84 239947
rect 84 239913 96 239947
rect -96 239907 96 239913
rect -96 239839 96 239845
rect -96 239805 -84 239839
rect 84 239805 96 239839
rect -96 239799 96 239805
rect -152 239746 -106 239758
rect -152 237370 -146 239746
rect -112 237370 -106 239746
rect -152 237358 -106 237370
rect 106 239746 152 239758
rect 106 237370 112 239746
rect 146 237370 152 239746
rect 106 237358 152 237370
rect -96 237311 96 237317
rect -96 237277 -84 237311
rect 84 237277 96 237311
rect -96 237271 96 237277
rect -96 237203 96 237209
rect -96 237169 -84 237203
rect 84 237169 96 237203
rect -96 237163 96 237169
rect -152 237110 -106 237122
rect -152 234734 -146 237110
rect -112 234734 -106 237110
rect -152 234722 -106 234734
rect 106 237110 152 237122
rect 106 234734 112 237110
rect 146 234734 152 237110
rect 106 234722 152 234734
rect -96 234675 96 234681
rect -96 234641 -84 234675
rect 84 234641 96 234675
rect -96 234635 96 234641
rect -96 234567 96 234573
rect -96 234533 -84 234567
rect 84 234533 96 234567
rect -96 234527 96 234533
rect -152 234474 -106 234486
rect -152 232098 -146 234474
rect -112 232098 -106 234474
rect -152 232086 -106 232098
rect 106 234474 152 234486
rect 106 232098 112 234474
rect 146 232098 152 234474
rect 106 232086 152 232098
rect -96 232039 96 232045
rect -96 232005 -84 232039
rect 84 232005 96 232039
rect -96 231999 96 232005
rect -96 231931 96 231937
rect -96 231897 -84 231931
rect 84 231897 96 231931
rect -96 231891 96 231897
rect -152 231838 -106 231850
rect -152 229462 -146 231838
rect -112 229462 -106 231838
rect -152 229450 -106 229462
rect 106 231838 152 231850
rect 106 229462 112 231838
rect 146 229462 152 231838
rect 106 229450 152 229462
rect -96 229403 96 229409
rect -96 229369 -84 229403
rect 84 229369 96 229403
rect -96 229363 96 229369
rect -96 229295 96 229301
rect -96 229261 -84 229295
rect 84 229261 96 229295
rect -96 229255 96 229261
rect -152 229202 -106 229214
rect -152 226826 -146 229202
rect -112 226826 -106 229202
rect -152 226814 -106 226826
rect 106 229202 152 229214
rect 106 226826 112 229202
rect 146 226826 152 229202
rect 106 226814 152 226826
rect -96 226767 96 226773
rect -96 226733 -84 226767
rect 84 226733 96 226767
rect -96 226727 96 226733
rect -96 226659 96 226665
rect -96 226625 -84 226659
rect 84 226625 96 226659
rect -96 226619 96 226625
rect -152 226566 -106 226578
rect -152 224190 -146 226566
rect -112 224190 -106 226566
rect -152 224178 -106 224190
rect 106 226566 152 226578
rect 106 224190 112 226566
rect 146 224190 152 226566
rect 106 224178 152 224190
rect -96 224131 96 224137
rect -96 224097 -84 224131
rect 84 224097 96 224131
rect -96 224091 96 224097
rect -96 224023 96 224029
rect -96 223989 -84 224023
rect 84 223989 96 224023
rect -96 223983 96 223989
rect -152 223930 -106 223942
rect -152 221554 -146 223930
rect -112 221554 -106 223930
rect -152 221542 -106 221554
rect 106 223930 152 223942
rect 106 221554 112 223930
rect 146 221554 152 223930
rect 106 221542 152 221554
rect -96 221495 96 221501
rect -96 221461 -84 221495
rect 84 221461 96 221495
rect -96 221455 96 221461
rect -96 221387 96 221393
rect -96 221353 -84 221387
rect 84 221353 96 221387
rect -96 221347 96 221353
rect -152 221294 -106 221306
rect -152 218918 -146 221294
rect -112 218918 -106 221294
rect -152 218906 -106 218918
rect 106 221294 152 221306
rect 106 218918 112 221294
rect 146 218918 152 221294
rect 106 218906 152 218918
rect -96 218859 96 218865
rect -96 218825 -84 218859
rect 84 218825 96 218859
rect -96 218819 96 218825
rect -96 218751 96 218757
rect -96 218717 -84 218751
rect 84 218717 96 218751
rect -96 218711 96 218717
rect -152 218658 -106 218670
rect -152 216282 -146 218658
rect -112 216282 -106 218658
rect -152 216270 -106 216282
rect 106 218658 152 218670
rect 106 216282 112 218658
rect 146 216282 152 218658
rect 106 216270 152 216282
rect -96 216223 96 216229
rect -96 216189 -84 216223
rect 84 216189 96 216223
rect -96 216183 96 216189
rect -96 216115 96 216121
rect -96 216081 -84 216115
rect 84 216081 96 216115
rect -96 216075 96 216081
rect -152 216022 -106 216034
rect -152 213646 -146 216022
rect -112 213646 -106 216022
rect -152 213634 -106 213646
rect 106 216022 152 216034
rect 106 213646 112 216022
rect 146 213646 152 216022
rect 106 213634 152 213646
rect -96 213587 96 213593
rect -96 213553 -84 213587
rect 84 213553 96 213587
rect -96 213547 96 213553
rect -96 213479 96 213485
rect -96 213445 -84 213479
rect 84 213445 96 213479
rect -96 213439 96 213445
rect -152 213386 -106 213398
rect -152 211010 -146 213386
rect -112 211010 -106 213386
rect -152 210998 -106 211010
rect 106 213386 152 213398
rect 106 211010 112 213386
rect 146 211010 152 213386
rect 106 210998 152 211010
rect -96 210951 96 210957
rect -96 210917 -84 210951
rect 84 210917 96 210951
rect -96 210911 96 210917
rect -96 210843 96 210849
rect -96 210809 -84 210843
rect 84 210809 96 210843
rect -96 210803 96 210809
rect -152 210750 -106 210762
rect -152 208374 -146 210750
rect -112 208374 -106 210750
rect -152 208362 -106 208374
rect 106 210750 152 210762
rect 106 208374 112 210750
rect 146 208374 152 210750
rect 106 208362 152 208374
rect -96 208315 96 208321
rect -96 208281 -84 208315
rect 84 208281 96 208315
rect -96 208275 96 208281
rect -96 208207 96 208213
rect -96 208173 -84 208207
rect 84 208173 96 208207
rect -96 208167 96 208173
rect -152 208114 -106 208126
rect -152 205738 -146 208114
rect -112 205738 -106 208114
rect -152 205726 -106 205738
rect 106 208114 152 208126
rect 106 205738 112 208114
rect 146 205738 152 208114
rect 106 205726 152 205738
rect -96 205679 96 205685
rect -96 205645 -84 205679
rect 84 205645 96 205679
rect -96 205639 96 205645
rect -96 205571 96 205577
rect -96 205537 -84 205571
rect 84 205537 96 205571
rect -96 205531 96 205537
rect -152 205478 -106 205490
rect -152 203102 -146 205478
rect -112 203102 -106 205478
rect -152 203090 -106 203102
rect 106 205478 152 205490
rect 106 203102 112 205478
rect 146 203102 152 205478
rect 106 203090 152 203102
rect -96 203043 96 203049
rect -96 203009 -84 203043
rect 84 203009 96 203043
rect -96 203003 96 203009
rect -96 202935 96 202941
rect -96 202901 -84 202935
rect 84 202901 96 202935
rect -96 202895 96 202901
rect -152 202842 -106 202854
rect -152 200466 -146 202842
rect -112 200466 -106 202842
rect -152 200454 -106 200466
rect 106 202842 152 202854
rect 106 200466 112 202842
rect 146 200466 152 202842
rect 106 200454 152 200466
rect -96 200407 96 200413
rect -96 200373 -84 200407
rect 84 200373 96 200407
rect -96 200367 96 200373
rect -96 200299 96 200305
rect -96 200265 -84 200299
rect 84 200265 96 200299
rect -96 200259 96 200265
rect -152 200206 -106 200218
rect -152 197830 -146 200206
rect -112 197830 -106 200206
rect -152 197818 -106 197830
rect 106 200206 152 200218
rect 106 197830 112 200206
rect 146 197830 152 200206
rect 106 197818 152 197830
rect -96 197771 96 197777
rect -96 197737 -84 197771
rect 84 197737 96 197771
rect -96 197731 96 197737
rect -96 197663 96 197669
rect -96 197629 -84 197663
rect 84 197629 96 197663
rect -96 197623 96 197629
rect -152 197570 -106 197582
rect -152 195194 -146 197570
rect -112 195194 -106 197570
rect -152 195182 -106 195194
rect 106 197570 152 197582
rect 106 195194 112 197570
rect 146 195194 152 197570
rect 106 195182 152 195194
rect -96 195135 96 195141
rect -96 195101 -84 195135
rect 84 195101 96 195135
rect -96 195095 96 195101
rect -96 195027 96 195033
rect -96 194993 -84 195027
rect 84 194993 96 195027
rect -96 194987 96 194993
rect -152 194934 -106 194946
rect -152 192558 -146 194934
rect -112 192558 -106 194934
rect -152 192546 -106 192558
rect 106 194934 152 194946
rect 106 192558 112 194934
rect 146 192558 152 194934
rect 106 192546 152 192558
rect -96 192499 96 192505
rect -96 192465 -84 192499
rect 84 192465 96 192499
rect -96 192459 96 192465
rect -96 192391 96 192397
rect -96 192357 -84 192391
rect 84 192357 96 192391
rect -96 192351 96 192357
rect -152 192298 -106 192310
rect -152 189922 -146 192298
rect -112 189922 -106 192298
rect -152 189910 -106 189922
rect 106 192298 152 192310
rect 106 189922 112 192298
rect 146 189922 152 192298
rect 106 189910 152 189922
rect -96 189863 96 189869
rect -96 189829 -84 189863
rect 84 189829 96 189863
rect -96 189823 96 189829
rect -96 189755 96 189761
rect -96 189721 -84 189755
rect 84 189721 96 189755
rect -96 189715 96 189721
rect -152 189662 -106 189674
rect -152 187286 -146 189662
rect -112 187286 -106 189662
rect -152 187274 -106 187286
rect 106 189662 152 189674
rect 106 187286 112 189662
rect 146 187286 152 189662
rect 106 187274 152 187286
rect -96 187227 96 187233
rect -96 187193 -84 187227
rect 84 187193 96 187227
rect -96 187187 96 187193
rect -96 187119 96 187125
rect -96 187085 -84 187119
rect 84 187085 96 187119
rect -96 187079 96 187085
rect -152 187026 -106 187038
rect -152 184650 -146 187026
rect -112 184650 -106 187026
rect -152 184638 -106 184650
rect 106 187026 152 187038
rect 106 184650 112 187026
rect 146 184650 152 187026
rect 106 184638 152 184650
rect -96 184591 96 184597
rect -96 184557 -84 184591
rect 84 184557 96 184591
rect -96 184551 96 184557
rect -96 184483 96 184489
rect -96 184449 -84 184483
rect 84 184449 96 184483
rect -96 184443 96 184449
rect -152 184390 -106 184402
rect -152 182014 -146 184390
rect -112 182014 -106 184390
rect -152 182002 -106 182014
rect 106 184390 152 184402
rect 106 182014 112 184390
rect 146 182014 152 184390
rect 106 182002 152 182014
rect -96 181955 96 181961
rect -96 181921 -84 181955
rect 84 181921 96 181955
rect -96 181915 96 181921
rect -96 181847 96 181853
rect -96 181813 -84 181847
rect 84 181813 96 181847
rect -96 181807 96 181813
rect -152 181754 -106 181766
rect -152 179378 -146 181754
rect -112 179378 -106 181754
rect -152 179366 -106 179378
rect 106 181754 152 181766
rect 106 179378 112 181754
rect 146 179378 152 181754
rect 106 179366 152 179378
rect -96 179319 96 179325
rect -96 179285 -84 179319
rect 84 179285 96 179319
rect -96 179279 96 179285
rect -96 179211 96 179217
rect -96 179177 -84 179211
rect 84 179177 96 179211
rect -96 179171 96 179177
rect -152 179118 -106 179130
rect -152 176742 -146 179118
rect -112 176742 -106 179118
rect -152 176730 -106 176742
rect 106 179118 152 179130
rect 106 176742 112 179118
rect 146 176742 152 179118
rect 106 176730 152 176742
rect -96 176683 96 176689
rect -96 176649 -84 176683
rect 84 176649 96 176683
rect -96 176643 96 176649
rect -96 176575 96 176581
rect -96 176541 -84 176575
rect 84 176541 96 176575
rect -96 176535 96 176541
rect -152 176482 -106 176494
rect -152 174106 -146 176482
rect -112 174106 -106 176482
rect -152 174094 -106 174106
rect 106 176482 152 176494
rect 106 174106 112 176482
rect 146 174106 152 176482
rect 106 174094 152 174106
rect -96 174047 96 174053
rect -96 174013 -84 174047
rect 84 174013 96 174047
rect -96 174007 96 174013
rect -96 173939 96 173945
rect -96 173905 -84 173939
rect 84 173905 96 173939
rect -96 173899 96 173905
rect -152 173846 -106 173858
rect -152 171470 -146 173846
rect -112 171470 -106 173846
rect -152 171458 -106 171470
rect 106 173846 152 173858
rect 106 171470 112 173846
rect 146 171470 152 173846
rect 106 171458 152 171470
rect -96 171411 96 171417
rect -96 171377 -84 171411
rect 84 171377 96 171411
rect -96 171371 96 171377
rect -96 171303 96 171309
rect -96 171269 -84 171303
rect 84 171269 96 171303
rect -96 171263 96 171269
rect -152 171210 -106 171222
rect -152 168834 -146 171210
rect -112 168834 -106 171210
rect -152 168822 -106 168834
rect 106 171210 152 171222
rect 106 168834 112 171210
rect 146 168834 152 171210
rect 106 168822 152 168834
rect -96 168775 96 168781
rect -96 168741 -84 168775
rect 84 168741 96 168775
rect -96 168735 96 168741
rect -96 168667 96 168673
rect -96 168633 -84 168667
rect 84 168633 96 168667
rect -96 168627 96 168633
rect -152 168574 -106 168586
rect -152 166198 -146 168574
rect -112 166198 -106 168574
rect -152 166186 -106 166198
rect 106 168574 152 168586
rect 106 166198 112 168574
rect 146 166198 152 168574
rect 106 166186 152 166198
rect -96 166139 96 166145
rect -96 166105 -84 166139
rect 84 166105 96 166139
rect -96 166099 96 166105
rect -96 166031 96 166037
rect -96 165997 -84 166031
rect 84 165997 96 166031
rect -96 165991 96 165997
rect -152 165938 -106 165950
rect -152 163562 -146 165938
rect -112 163562 -106 165938
rect -152 163550 -106 163562
rect 106 165938 152 165950
rect 106 163562 112 165938
rect 146 163562 152 165938
rect 106 163550 152 163562
rect -96 163503 96 163509
rect -96 163469 -84 163503
rect 84 163469 96 163503
rect -96 163463 96 163469
rect -96 163395 96 163401
rect -96 163361 -84 163395
rect 84 163361 96 163395
rect -96 163355 96 163361
rect -152 163302 -106 163314
rect -152 160926 -146 163302
rect -112 160926 -106 163302
rect -152 160914 -106 160926
rect 106 163302 152 163314
rect 106 160926 112 163302
rect 146 160926 152 163302
rect 106 160914 152 160926
rect -96 160867 96 160873
rect -96 160833 -84 160867
rect 84 160833 96 160867
rect -96 160827 96 160833
rect -96 160759 96 160765
rect -96 160725 -84 160759
rect 84 160725 96 160759
rect -96 160719 96 160725
rect -152 160666 -106 160678
rect -152 158290 -146 160666
rect -112 158290 -106 160666
rect -152 158278 -106 158290
rect 106 160666 152 160678
rect 106 158290 112 160666
rect 146 158290 152 160666
rect 106 158278 152 158290
rect -96 158231 96 158237
rect -96 158197 -84 158231
rect 84 158197 96 158231
rect -96 158191 96 158197
rect -96 158123 96 158129
rect -96 158089 -84 158123
rect 84 158089 96 158123
rect -96 158083 96 158089
rect -152 158030 -106 158042
rect -152 155654 -146 158030
rect -112 155654 -106 158030
rect -152 155642 -106 155654
rect 106 158030 152 158042
rect 106 155654 112 158030
rect 146 155654 152 158030
rect 106 155642 152 155654
rect -96 155595 96 155601
rect -96 155561 -84 155595
rect 84 155561 96 155595
rect -96 155555 96 155561
rect -96 155487 96 155493
rect -96 155453 -84 155487
rect 84 155453 96 155487
rect -96 155447 96 155453
rect -152 155394 -106 155406
rect -152 153018 -146 155394
rect -112 153018 -106 155394
rect -152 153006 -106 153018
rect 106 155394 152 155406
rect 106 153018 112 155394
rect 146 153018 152 155394
rect 106 153006 152 153018
rect -96 152959 96 152965
rect -96 152925 -84 152959
rect 84 152925 96 152959
rect -96 152919 96 152925
rect -96 152851 96 152857
rect -96 152817 -84 152851
rect 84 152817 96 152851
rect -96 152811 96 152817
rect -152 152758 -106 152770
rect -152 150382 -146 152758
rect -112 150382 -106 152758
rect -152 150370 -106 150382
rect 106 152758 152 152770
rect 106 150382 112 152758
rect 146 150382 152 152758
rect 106 150370 152 150382
rect -96 150323 96 150329
rect -96 150289 -84 150323
rect 84 150289 96 150323
rect -96 150283 96 150289
rect -96 150215 96 150221
rect -96 150181 -84 150215
rect 84 150181 96 150215
rect -96 150175 96 150181
rect -152 150122 -106 150134
rect -152 147746 -146 150122
rect -112 147746 -106 150122
rect -152 147734 -106 147746
rect 106 150122 152 150134
rect 106 147746 112 150122
rect 146 147746 152 150122
rect 106 147734 152 147746
rect -96 147687 96 147693
rect -96 147653 -84 147687
rect 84 147653 96 147687
rect -96 147647 96 147653
rect -96 147579 96 147585
rect -96 147545 -84 147579
rect 84 147545 96 147579
rect -96 147539 96 147545
rect -152 147486 -106 147498
rect -152 145110 -146 147486
rect -112 145110 -106 147486
rect -152 145098 -106 145110
rect 106 147486 152 147498
rect 106 145110 112 147486
rect 146 145110 152 147486
rect 106 145098 152 145110
rect -96 145051 96 145057
rect -96 145017 -84 145051
rect 84 145017 96 145051
rect -96 145011 96 145017
rect -96 144943 96 144949
rect -96 144909 -84 144943
rect 84 144909 96 144943
rect -96 144903 96 144909
rect -152 144850 -106 144862
rect -152 142474 -146 144850
rect -112 142474 -106 144850
rect -152 142462 -106 142474
rect 106 144850 152 144862
rect 106 142474 112 144850
rect 146 142474 152 144850
rect 106 142462 152 142474
rect -96 142415 96 142421
rect -96 142381 -84 142415
rect 84 142381 96 142415
rect -96 142375 96 142381
rect -96 142307 96 142313
rect -96 142273 -84 142307
rect 84 142273 96 142307
rect -96 142267 96 142273
rect -152 142214 -106 142226
rect -152 139838 -146 142214
rect -112 139838 -106 142214
rect -152 139826 -106 139838
rect 106 142214 152 142226
rect 106 139838 112 142214
rect 146 139838 152 142214
rect 106 139826 152 139838
rect -96 139779 96 139785
rect -96 139745 -84 139779
rect 84 139745 96 139779
rect -96 139739 96 139745
rect -96 139671 96 139677
rect -96 139637 -84 139671
rect 84 139637 96 139671
rect -96 139631 96 139637
rect -152 139578 -106 139590
rect -152 137202 -146 139578
rect -112 137202 -106 139578
rect -152 137190 -106 137202
rect 106 139578 152 139590
rect 106 137202 112 139578
rect 146 137202 152 139578
rect 106 137190 152 137202
rect -96 137143 96 137149
rect -96 137109 -84 137143
rect 84 137109 96 137143
rect -96 137103 96 137109
rect -96 137035 96 137041
rect -96 137001 -84 137035
rect 84 137001 96 137035
rect -96 136995 96 137001
rect -152 136942 -106 136954
rect -152 134566 -146 136942
rect -112 134566 -106 136942
rect -152 134554 -106 134566
rect 106 136942 152 136954
rect 106 134566 112 136942
rect 146 134566 152 136942
rect 106 134554 152 134566
rect -96 134507 96 134513
rect -96 134473 -84 134507
rect 84 134473 96 134507
rect -96 134467 96 134473
rect -96 134399 96 134405
rect -96 134365 -84 134399
rect 84 134365 96 134399
rect -96 134359 96 134365
rect -152 134306 -106 134318
rect -152 131930 -146 134306
rect -112 131930 -106 134306
rect -152 131918 -106 131930
rect 106 134306 152 134318
rect 106 131930 112 134306
rect 146 131930 152 134306
rect 106 131918 152 131930
rect -96 131871 96 131877
rect -96 131837 -84 131871
rect 84 131837 96 131871
rect -96 131831 96 131837
rect -96 131763 96 131769
rect -96 131729 -84 131763
rect 84 131729 96 131763
rect -96 131723 96 131729
rect -152 131670 -106 131682
rect -152 129294 -146 131670
rect -112 129294 -106 131670
rect -152 129282 -106 129294
rect 106 131670 152 131682
rect 106 129294 112 131670
rect 146 129294 152 131670
rect 106 129282 152 129294
rect -96 129235 96 129241
rect -96 129201 -84 129235
rect 84 129201 96 129235
rect -96 129195 96 129201
rect -96 129127 96 129133
rect -96 129093 -84 129127
rect 84 129093 96 129127
rect -96 129087 96 129093
rect -152 129034 -106 129046
rect -152 126658 -146 129034
rect -112 126658 -106 129034
rect -152 126646 -106 126658
rect 106 129034 152 129046
rect 106 126658 112 129034
rect 146 126658 152 129034
rect 106 126646 152 126658
rect -96 126599 96 126605
rect -96 126565 -84 126599
rect 84 126565 96 126599
rect -96 126559 96 126565
rect -96 126491 96 126497
rect -96 126457 -84 126491
rect 84 126457 96 126491
rect -96 126451 96 126457
rect -152 126398 -106 126410
rect -152 124022 -146 126398
rect -112 124022 -106 126398
rect -152 124010 -106 124022
rect 106 126398 152 126410
rect 106 124022 112 126398
rect 146 124022 152 126398
rect 106 124010 152 124022
rect -96 123963 96 123969
rect -96 123929 -84 123963
rect 84 123929 96 123963
rect -96 123923 96 123929
rect -96 123855 96 123861
rect -96 123821 -84 123855
rect 84 123821 96 123855
rect -96 123815 96 123821
rect -152 123762 -106 123774
rect -152 121386 -146 123762
rect -112 121386 -106 123762
rect -152 121374 -106 121386
rect 106 123762 152 123774
rect 106 121386 112 123762
rect 146 121386 152 123762
rect 106 121374 152 121386
rect -96 121327 96 121333
rect -96 121293 -84 121327
rect 84 121293 96 121327
rect -96 121287 96 121293
rect -96 121219 96 121225
rect -96 121185 -84 121219
rect 84 121185 96 121219
rect -96 121179 96 121185
rect -152 121126 -106 121138
rect -152 118750 -146 121126
rect -112 118750 -106 121126
rect -152 118738 -106 118750
rect 106 121126 152 121138
rect 106 118750 112 121126
rect 146 118750 152 121126
rect 106 118738 152 118750
rect -96 118691 96 118697
rect -96 118657 -84 118691
rect 84 118657 96 118691
rect -96 118651 96 118657
rect -96 118583 96 118589
rect -96 118549 -84 118583
rect 84 118549 96 118583
rect -96 118543 96 118549
rect -152 118490 -106 118502
rect -152 116114 -146 118490
rect -112 116114 -106 118490
rect -152 116102 -106 116114
rect 106 118490 152 118502
rect 106 116114 112 118490
rect 146 116114 152 118490
rect 106 116102 152 116114
rect -96 116055 96 116061
rect -96 116021 -84 116055
rect 84 116021 96 116055
rect -96 116015 96 116021
rect -96 115947 96 115953
rect -96 115913 -84 115947
rect 84 115913 96 115947
rect -96 115907 96 115913
rect -152 115854 -106 115866
rect -152 113478 -146 115854
rect -112 113478 -106 115854
rect -152 113466 -106 113478
rect 106 115854 152 115866
rect 106 113478 112 115854
rect 146 113478 152 115854
rect 106 113466 152 113478
rect -96 113419 96 113425
rect -96 113385 -84 113419
rect 84 113385 96 113419
rect -96 113379 96 113385
rect -96 113311 96 113317
rect -96 113277 -84 113311
rect 84 113277 96 113311
rect -96 113271 96 113277
rect -152 113218 -106 113230
rect -152 110842 -146 113218
rect -112 110842 -106 113218
rect -152 110830 -106 110842
rect 106 113218 152 113230
rect 106 110842 112 113218
rect 146 110842 152 113218
rect 106 110830 152 110842
rect -96 110783 96 110789
rect -96 110749 -84 110783
rect 84 110749 96 110783
rect -96 110743 96 110749
rect -96 110675 96 110681
rect -96 110641 -84 110675
rect 84 110641 96 110675
rect -96 110635 96 110641
rect -152 110582 -106 110594
rect -152 108206 -146 110582
rect -112 108206 -106 110582
rect -152 108194 -106 108206
rect 106 110582 152 110594
rect 106 108206 112 110582
rect 146 108206 152 110582
rect 106 108194 152 108206
rect -96 108147 96 108153
rect -96 108113 -84 108147
rect 84 108113 96 108147
rect -96 108107 96 108113
rect -96 108039 96 108045
rect -96 108005 -84 108039
rect 84 108005 96 108039
rect -96 107999 96 108005
rect -152 107946 -106 107958
rect -152 105570 -146 107946
rect -112 105570 -106 107946
rect -152 105558 -106 105570
rect 106 107946 152 107958
rect 106 105570 112 107946
rect 146 105570 152 107946
rect 106 105558 152 105570
rect -96 105511 96 105517
rect -96 105477 -84 105511
rect 84 105477 96 105511
rect -96 105471 96 105477
rect -96 105403 96 105409
rect -96 105369 -84 105403
rect 84 105369 96 105403
rect -96 105363 96 105369
rect -152 105310 -106 105322
rect -152 102934 -146 105310
rect -112 102934 -106 105310
rect -152 102922 -106 102934
rect 106 105310 152 105322
rect 106 102934 112 105310
rect 146 102934 152 105310
rect 106 102922 152 102934
rect -96 102875 96 102881
rect -96 102841 -84 102875
rect 84 102841 96 102875
rect -96 102835 96 102841
rect -96 102767 96 102773
rect -96 102733 -84 102767
rect 84 102733 96 102767
rect -96 102727 96 102733
rect -152 102674 -106 102686
rect -152 100298 -146 102674
rect -112 100298 -106 102674
rect -152 100286 -106 100298
rect 106 102674 152 102686
rect 106 100298 112 102674
rect 146 100298 152 102674
rect 106 100286 152 100298
rect -96 100239 96 100245
rect -96 100205 -84 100239
rect 84 100205 96 100239
rect -96 100199 96 100205
rect -96 100131 96 100137
rect -96 100097 -84 100131
rect 84 100097 96 100131
rect -96 100091 96 100097
rect -152 100038 -106 100050
rect -152 97662 -146 100038
rect -112 97662 -106 100038
rect -152 97650 -106 97662
rect 106 100038 152 100050
rect 106 97662 112 100038
rect 146 97662 152 100038
rect 106 97650 152 97662
rect -96 97603 96 97609
rect -96 97569 -84 97603
rect 84 97569 96 97603
rect -96 97563 96 97569
rect -96 97495 96 97501
rect -96 97461 -84 97495
rect 84 97461 96 97495
rect -96 97455 96 97461
rect -152 97402 -106 97414
rect -152 95026 -146 97402
rect -112 95026 -106 97402
rect -152 95014 -106 95026
rect 106 97402 152 97414
rect 106 95026 112 97402
rect 146 95026 152 97402
rect 106 95014 152 95026
rect -96 94967 96 94973
rect -96 94933 -84 94967
rect 84 94933 96 94967
rect -96 94927 96 94933
rect -96 94859 96 94865
rect -96 94825 -84 94859
rect 84 94825 96 94859
rect -96 94819 96 94825
rect -152 94766 -106 94778
rect -152 92390 -146 94766
rect -112 92390 -106 94766
rect -152 92378 -106 92390
rect 106 94766 152 94778
rect 106 92390 112 94766
rect 146 92390 152 94766
rect 106 92378 152 92390
rect -96 92331 96 92337
rect -96 92297 -84 92331
rect 84 92297 96 92331
rect -96 92291 96 92297
rect -96 92223 96 92229
rect -96 92189 -84 92223
rect 84 92189 96 92223
rect -96 92183 96 92189
rect -152 92130 -106 92142
rect -152 89754 -146 92130
rect -112 89754 -106 92130
rect -152 89742 -106 89754
rect 106 92130 152 92142
rect 106 89754 112 92130
rect 146 89754 152 92130
rect 106 89742 152 89754
rect -96 89695 96 89701
rect -96 89661 -84 89695
rect 84 89661 96 89695
rect -96 89655 96 89661
rect -96 89587 96 89593
rect -96 89553 -84 89587
rect 84 89553 96 89587
rect -96 89547 96 89553
rect -152 89494 -106 89506
rect -152 87118 -146 89494
rect -112 87118 -106 89494
rect -152 87106 -106 87118
rect 106 89494 152 89506
rect 106 87118 112 89494
rect 146 87118 152 89494
rect 106 87106 152 87118
rect -96 87059 96 87065
rect -96 87025 -84 87059
rect 84 87025 96 87059
rect -96 87019 96 87025
rect -96 86951 96 86957
rect -96 86917 -84 86951
rect 84 86917 96 86951
rect -96 86911 96 86917
rect -152 86858 -106 86870
rect -152 84482 -146 86858
rect -112 84482 -106 86858
rect -152 84470 -106 84482
rect 106 86858 152 86870
rect 106 84482 112 86858
rect 146 84482 152 86858
rect 106 84470 152 84482
rect -96 84423 96 84429
rect -96 84389 -84 84423
rect 84 84389 96 84423
rect -96 84383 96 84389
rect -96 84315 96 84321
rect -96 84281 -84 84315
rect 84 84281 96 84315
rect -96 84275 96 84281
rect -152 84222 -106 84234
rect -152 81846 -146 84222
rect -112 81846 -106 84222
rect -152 81834 -106 81846
rect 106 84222 152 84234
rect 106 81846 112 84222
rect 146 81846 152 84222
rect 106 81834 152 81846
rect -96 81787 96 81793
rect -96 81753 -84 81787
rect 84 81753 96 81787
rect -96 81747 96 81753
rect -96 81679 96 81685
rect -96 81645 -84 81679
rect 84 81645 96 81679
rect -96 81639 96 81645
rect -152 81586 -106 81598
rect -152 79210 -146 81586
rect -112 79210 -106 81586
rect -152 79198 -106 79210
rect 106 81586 152 81598
rect 106 79210 112 81586
rect 146 79210 152 81586
rect 106 79198 152 79210
rect -96 79151 96 79157
rect -96 79117 -84 79151
rect 84 79117 96 79151
rect -96 79111 96 79117
rect -96 79043 96 79049
rect -96 79009 -84 79043
rect 84 79009 96 79043
rect -96 79003 96 79009
rect -152 78950 -106 78962
rect -152 76574 -146 78950
rect -112 76574 -106 78950
rect -152 76562 -106 76574
rect 106 78950 152 78962
rect 106 76574 112 78950
rect 146 76574 152 78950
rect 106 76562 152 76574
rect -96 76515 96 76521
rect -96 76481 -84 76515
rect 84 76481 96 76515
rect -96 76475 96 76481
rect -96 76407 96 76413
rect -96 76373 -84 76407
rect 84 76373 96 76407
rect -96 76367 96 76373
rect -152 76314 -106 76326
rect -152 73938 -146 76314
rect -112 73938 -106 76314
rect -152 73926 -106 73938
rect 106 76314 152 76326
rect 106 73938 112 76314
rect 146 73938 152 76314
rect 106 73926 152 73938
rect -96 73879 96 73885
rect -96 73845 -84 73879
rect 84 73845 96 73879
rect -96 73839 96 73845
rect -96 73771 96 73777
rect -96 73737 -84 73771
rect 84 73737 96 73771
rect -96 73731 96 73737
rect -152 73678 -106 73690
rect -152 71302 -146 73678
rect -112 71302 -106 73678
rect -152 71290 -106 71302
rect 106 73678 152 73690
rect 106 71302 112 73678
rect 146 71302 152 73678
rect 106 71290 152 71302
rect -96 71243 96 71249
rect -96 71209 -84 71243
rect 84 71209 96 71243
rect -96 71203 96 71209
rect -96 71135 96 71141
rect -96 71101 -84 71135
rect 84 71101 96 71135
rect -96 71095 96 71101
rect -152 71042 -106 71054
rect -152 68666 -146 71042
rect -112 68666 -106 71042
rect -152 68654 -106 68666
rect 106 71042 152 71054
rect 106 68666 112 71042
rect 146 68666 152 71042
rect 106 68654 152 68666
rect -96 68607 96 68613
rect -96 68573 -84 68607
rect 84 68573 96 68607
rect -96 68567 96 68573
rect -96 68499 96 68505
rect -96 68465 -84 68499
rect 84 68465 96 68499
rect -96 68459 96 68465
rect -152 68406 -106 68418
rect -152 66030 -146 68406
rect -112 66030 -106 68406
rect -152 66018 -106 66030
rect 106 68406 152 68418
rect 106 66030 112 68406
rect 146 66030 152 68406
rect 106 66018 152 66030
rect -96 65971 96 65977
rect -96 65937 -84 65971
rect 84 65937 96 65971
rect -96 65931 96 65937
rect -96 65863 96 65869
rect -96 65829 -84 65863
rect 84 65829 96 65863
rect -96 65823 96 65829
rect -152 65770 -106 65782
rect -152 63394 -146 65770
rect -112 63394 -106 65770
rect -152 63382 -106 63394
rect 106 65770 152 65782
rect 106 63394 112 65770
rect 146 63394 152 65770
rect 106 63382 152 63394
rect -96 63335 96 63341
rect -96 63301 -84 63335
rect 84 63301 96 63335
rect -96 63295 96 63301
rect -96 63227 96 63233
rect -96 63193 -84 63227
rect 84 63193 96 63227
rect -96 63187 96 63193
rect -152 63134 -106 63146
rect -152 60758 -146 63134
rect -112 60758 -106 63134
rect -152 60746 -106 60758
rect 106 63134 152 63146
rect 106 60758 112 63134
rect 146 60758 152 63134
rect 106 60746 152 60758
rect -96 60699 96 60705
rect -96 60665 -84 60699
rect 84 60665 96 60699
rect -96 60659 96 60665
rect -96 60591 96 60597
rect -96 60557 -84 60591
rect 84 60557 96 60591
rect -96 60551 96 60557
rect -152 60498 -106 60510
rect -152 58122 -146 60498
rect -112 58122 -106 60498
rect -152 58110 -106 58122
rect 106 60498 152 60510
rect 106 58122 112 60498
rect 146 58122 152 60498
rect 106 58110 152 58122
rect -96 58063 96 58069
rect -96 58029 -84 58063
rect 84 58029 96 58063
rect -96 58023 96 58029
rect -96 57955 96 57961
rect -96 57921 -84 57955
rect 84 57921 96 57955
rect -96 57915 96 57921
rect -152 57862 -106 57874
rect -152 55486 -146 57862
rect -112 55486 -106 57862
rect -152 55474 -106 55486
rect 106 57862 152 57874
rect 106 55486 112 57862
rect 146 55486 152 57862
rect 106 55474 152 55486
rect -96 55427 96 55433
rect -96 55393 -84 55427
rect 84 55393 96 55427
rect -96 55387 96 55393
rect -96 55319 96 55325
rect -96 55285 -84 55319
rect 84 55285 96 55319
rect -96 55279 96 55285
rect -152 55226 -106 55238
rect -152 52850 -146 55226
rect -112 52850 -106 55226
rect -152 52838 -106 52850
rect 106 55226 152 55238
rect 106 52850 112 55226
rect 146 52850 152 55226
rect 106 52838 152 52850
rect -96 52791 96 52797
rect -96 52757 -84 52791
rect 84 52757 96 52791
rect -96 52751 96 52757
rect -96 52683 96 52689
rect -96 52649 -84 52683
rect 84 52649 96 52683
rect -96 52643 96 52649
rect -152 52590 -106 52602
rect -152 50214 -146 52590
rect -112 50214 -106 52590
rect -152 50202 -106 50214
rect 106 52590 152 52602
rect 106 50214 112 52590
rect 146 50214 152 52590
rect 106 50202 152 50214
rect -96 50155 96 50161
rect -96 50121 -84 50155
rect 84 50121 96 50155
rect -96 50115 96 50121
rect -96 50047 96 50053
rect -96 50013 -84 50047
rect 84 50013 96 50047
rect -96 50007 96 50013
rect -152 49954 -106 49966
rect -152 47578 -146 49954
rect -112 47578 -106 49954
rect -152 47566 -106 47578
rect 106 49954 152 49966
rect 106 47578 112 49954
rect 146 47578 152 49954
rect 106 47566 152 47578
rect -96 47519 96 47525
rect -96 47485 -84 47519
rect 84 47485 96 47519
rect -96 47479 96 47485
rect -96 47411 96 47417
rect -96 47377 -84 47411
rect 84 47377 96 47411
rect -96 47371 96 47377
rect -152 47318 -106 47330
rect -152 44942 -146 47318
rect -112 44942 -106 47318
rect -152 44930 -106 44942
rect 106 47318 152 47330
rect 106 44942 112 47318
rect 146 44942 152 47318
rect 106 44930 152 44942
rect -96 44883 96 44889
rect -96 44849 -84 44883
rect 84 44849 96 44883
rect -96 44843 96 44849
rect -96 44775 96 44781
rect -96 44741 -84 44775
rect 84 44741 96 44775
rect -96 44735 96 44741
rect -152 44682 -106 44694
rect -152 42306 -146 44682
rect -112 42306 -106 44682
rect -152 42294 -106 42306
rect 106 44682 152 44694
rect 106 42306 112 44682
rect 146 42306 152 44682
rect 106 42294 152 42306
rect -96 42247 96 42253
rect -96 42213 -84 42247
rect 84 42213 96 42247
rect -96 42207 96 42213
rect -96 42139 96 42145
rect -96 42105 -84 42139
rect 84 42105 96 42139
rect -96 42099 96 42105
rect -152 42046 -106 42058
rect -152 39670 -146 42046
rect -112 39670 -106 42046
rect -152 39658 -106 39670
rect 106 42046 152 42058
rect 106 39670 112 42046
rect 146 39670 152 42046
rect 106 39658 152 39670
rect -96 39611 96 39617
rect -96 39577 -84 39611
rect 84 39577 96 39611
rect -96 39571 96 39577
rect -96 39503 96 39509
rect -96 39469 -84 39503
rect 84 39469 96 39503
rect -96 39463 96 39469
rect -152 39410 -106 39422
rect -152 37034 -146 39410
rect -112 37034 -106 39410
rect -152 37022 -106 37034
rect 106 39410 152 39422
rect 106 37034 112 39410
rect 146 37034 152 39410
rect 106 37022 152 37034
rect -96 36975 96 36981
rect -96 36941 -84 36975
rect 84 36941 96 36975
rect -96 36935 96 36941
rect -96 36867 96 36873
rect -96 36833 -84 36867
rect 84 36833 96 36867
rect -96 36827 96 36833
rect -152 36774 -106 36786
rect -152 34398 -146 36774
rect -112 34398 -106 36774
rect -152 34386 -106 34398
rect 106 36774 152 36786
rect 106 34398 112 36774
rect 146 34398 152 36774
rect 106 34386 152 34398
rect -96 34339 96 34345
rect -96 34305 -84 34339
rect 84 34305 96 34339
rect -96 34299 96 34305
rect -96 34231 96 34237
rect -96 34197 -84 34231
rect 84 34197 96 34231
rect -96 34191 96 34197
rect -152 34138 -106 34150
rect -152 31762 -146 34138
rect -112 31762 -106 34138
rect -152 31750 -106 31762
rect 106 34138 152 34150
rect 106 31762 112 34138
rect 146 31762 152 34138
rect 106 31750 152 31762
rect -96 31703 96 31709
rect -96 31669 -84 31703
rect 84 31669 96 31703
rect -96 31663 96 31669
rect -96 31595 96 31601
rect -96 31561 -84 31595
rect 84 31561 96 31595
rect -96 31555 96 31561
rect -152 31502 -106 31514
rect -152 29126 -146 31502
rect -112 29126 -106 31502
rect -152 29114 -106 29126
rect 106 31502 152 31514
rect 106 29126 112 31502
rect 146 29126 152 31502
rect 106 29114 152 29126
rect -96 29067 96 29073
rect -96 29033 -84 29067
rect 84 29033 96 29067
rect -96 29027 96 29033
rect -96 28959 96 28965
rect -96 28925 -84 28959
rect 84 28925 96 28959
rect -96 28919 96 28925
rect -152 28866 -106 28878
rect -152 26490 -146 28866
rect -112 26490 -106 28866
rect -152 26478 -106 26490
rect 106 28866 152 28878
rect 106 26490 112 28866
rect 146 26490 152 28866
rect 106 26478 152 26490
rect -96 26431 96 26437
rect -96 26397 -84 26431
rect 84 26397 96 26431
rect -96 26391 96 26397
rect -96 26323 96 26329
rect -96 26289 -84 26323
rect 84 26289 96 26323
rect -96 26283 96 26289
rect -152 26230 -106 26242
rect -152 23854 -146 26230
rect -112 23854 -106 26230
rect -152 23842 -106 23854
rect 106 26230 152 26242
rect 106 23854 112 26230
rect 146 23854 152 26230
rect 106 23842 152 23854
rect -96 23795 96 23801
rect -96 23761 -84 23795
rect 84 23761 96 23795
rect -96 23755 96 23761
rect -96 23687 96 23693
rect -96 23653 -84 23687
rect 84 23653 96 23687
rect -96 23647 96 23653
rect -152 23594 -106 23606
rect -152 21218 -146 23594
rect -112 21218 -106 23594
rect -152 21206 -106 21218
rect 106 23594 152 23606
rect 106 21218 112 23594
rect 146 21218 152 23594
rect 106 21206 152 21218
rect -96 21159 96 21165
rect -96 21125 -84 21159
rect 84 21125 96 21159
rect -96 21119 96 21125
rect -96 21051 96 21057
rect -96 21017 -84 21051
rect 84 21017 96 21051
rect -96 21011 96 21017
rect -152 20958 -106 20970
rect -152 18582 -146 20958
rect -112 18582 -106 20958
rect -152 18570 -106 18582
rect 106 20958 152 20970
rect 106 18582 112 20958
rect 146 18582 152 20958
rect 106 18570 152 18582
rect -96 18523 96 18529
rect -96 18489 -84 18523
rect 84 18489 96 18523
rect -96 18483 96 18489
rect -96 18415 96 18421
rect -96 18381 -84 18415
rect 84 18381 96 18415
rect -96 18375 96 18381
rect -152 18322 -106 18334
rect -152 15946 -146 18322
rect -112 15946 -106 18322
rect -152 15934 -106 15946
rect 106 18322 152 18334
rect 106 15946 112 18322
rect 146 15946 152 18322
rect 106 15934 152 15946
rect -96 15887 96 15893
rect -96 15853 -84 15887
rect 84 15853 96 15887
rect -96 15847 96 15853
rect -96 15779 96 15785
rect -96 15745 -84 15779
rect 84 15745 96 15779
rect -96 15739 96 15745
rect -152 15686 -106 15698
rect -152 13310 -146 15686
rect -112 13310 -106 15686
rect -152 13298 -106 13310
rect 106 15686 152 15698
rect 106 13310 112 15686
rect 146 13310 152 15686
rect 106 13298 152 13310
rect -96 13251 96 13257
rect -96 13217 -84 13251
rect 84 13217 96 13251
rect -96 13211 96 13217
rect -96 13143 96 13149
rect -96 13109 -84 13143
rect 84 13109 96 13143
rect -96 13103 96 13109
rect -152 13050 -106 13062
rect -152 10674 -146 13050
rect -112 10674 -106 13050
rect -152 10662 -106 10674
rect 106 13050 152 13062
rect 106 10674 112 13050
rect 146 10674 152 13050
rect 106 10662 152 10674
rect -96 10615 96 10621
rect -96 10581 -84 10615
rect 84 10581 96 10615
rect -96 10575 96 10581
rect -96 10507 96 10513
rect -96 10473 -84 10507
rect 84 10473 96 10507
rect -96 10467 96 10473
rect -152 10414 -106 10426
rect -152 8038 -146 10414
rect -112 8038 -106 10414
rect -152 8026 -106 8038
rect 106 10414 152 10426
rect 106 8038 112 10414
rect 146 8038 152 10414
rect 106 8026 152 8038
rect -96 7979 96 7985
rect -96 7945 -84 7979
rect 84 7945 96 7979
rect -96 7939 96 7945
rect -96 7871 96 7877
rect -96 7837 -84 7871
rect 84 7837 96 7871
rect -96 7831 96 7837
rect -152 7778 -106 7790
rect -152 5402 -146 7778
rect -112 5402 -106 7778
rect -152 5390 -106 5402
rect 106 7778 152 7790
rect 106 5402 112 7778
rect 146 5402 152 7778
rect 106 5390 152 5402
rect -96 5343 96 5349
rect -96 5309 -84 5343
rect 84 5309 96 5343
rect -96 5303 96 5309
rect -96 5235 96 5241
rect -96 5201 -84 5235
rect 84 5201 96 5235
rect -96 5195 96 5201
rect -152 5142 -106 5154
rect -152 2766 -146 5142
rect -112 2766 -106 5142
rect -152 2754 -106 2766
rect 106 5142 152 5154
rect 106 2766 112 5142
rect 146 2766 152 5142
rect 106 2754 152 2766
rect -96 2707 96 2713
rect -96 2673 -84 2707
rect 84 2673 96 2707
rect -96 2667 96 2673
rect -96 2599 96 2605
rect -96 2565 -84 2599
rect 84 2565 96 2599
rect -96 2559 96 2565
rect -152 2506 -106 2518
rect -152 130 -146 2506
rect -112 130 -106 2506
rect -152 118 -106 130
rect 106 2506 152 2518
rect 106 130 112 2506
rect 146 130 152 2506
rect 106 118 152 130
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -130 -106 -118
rect -152 -2506 -146 -130
rect -112 -2506 -106 -130
rect -152 -2518 -106 -2506
rect 106 -130 152 -118
rect 106 -2506 112 -130
rect 146 -2506 152 -130
rect 106 -2518 152 -2506
rect -96 -2565 96 -2559
rect -96 -2599 -84 -2565
rect 84 -2599 96 -2565
rect -96 -2605 96 -2599
rect -96 -2673 96 -2667
rect -96 -2707 -84 -2673
rect 84 -2707 96 -2673
rect -96 -2713 96 -2707
rect -152 -2766 -106 -2754
rect -152 -5142 -146 -2766
rect -112 -5142 -106 -2766
rect -152 -5154 -106 -5142
rect 106 -2766 152 -2754
rect 106 -5142 112 -2766
rect 146 -5142 152 -2766
rect 106 -5154 152 -5142
rect -96 -5201 96 -5195
rect -96 -5235 -84 -5201
rect 84 -5235 96 -5201
rect -96 -5241 96 -5235
rect -96 -5309 96 -5303
rect -96 -5343 -84 -5309
rect 84 -5343 96 -5309
rect -96 -5349 96 -5343
rect -152 -5402 -106 -5390
rect -152 -7778 -146 -5402
rect -112 -7778 -106 -5402
rect -152 -7790 -106 -7778
rect 106 -5402 152 -5390
rect 106 -7778 112 -5402
rect 146 -7778 152 -5402
rect 106 -7790 152 -7778
rect -96 -7837 96 -7831
rect -96 -7871 -84 -7837
rect 84 -7871 96 -7837
rect -96 -7877 96 -7871
rect -96 -7945 96 -7939
rect -96 -7979 -84 -7945
rect 84 -7979 96 -7945
rect -96 -7985 96 -7979
rect -152 -8038 -106 -8026
rect -152 -10414 -146 -8038
rect -112 -10414 -106 -8038
rect -152 -10426 -106 -10414
rect 106 -8038 152 -8026
rect 106 -10414 112 -8038
rect 146 -10414 152 -8038
rect 106 -10426 152 -10414
rect -96 -10473 96 -10467
rect -96 -10507 -84 -10473
rect 84 -10507 96 -10473
rect -96 -10513 96 -10507
rect -96 -10581 96 -10575
rect -96 -10615 -84 -10581
rect 84 -10615 96 -10581
rect -96 -10621 96 -10615
rect -152 -10674 -106 -10662
rect -152 -13050 -146 -10674
rect -112 -13050 -106 -10674
rect -152 -13062 -106 -13050
rect 106 -10674 152 -10662
rect 106 -13050 112 -10674
rect 146 -13050 152 -10674
rect 106 -13062 152 -13050
rect -96 -13109 96 -13103
rect -96 -13143 -84 -13109
rect 84 -13143 96 -13109
rect -96 -13149 96 -13143
rect -96 -13217 96 -13211
rect -96 -13251 -84 -13217
rect 84 -13251 96 -13217
rect -96 -13257 96 -13251
rect -152 -13310 -106 -13298
rect -152 -15686 -146 -13310
rect -112 -15686 -106 -13310
rect -152 -15698 -106 -15686
rect 106 -13310 152 -13298
rect 106 -15686 112 -13310
rect 146 -15686 152 -13310
rect 106 -15698 152 -15686
rect -96 -15745 96 -15739
rect -96 -15779 -84 -15745
rect 84 -15779 96 -15745
rect -96 -15785 96 -15779
rect -96 -15853 96 -15847
rect -96 -15887 -84 -15853
rect 84 -15887 96 -15853
rect -96 -15893 96 -15887
rect -152 -15946 -106 -15934
rect -152 -18322 -146 -15946
rect -112 -18322 -106 -15946
rect -152 -18334 -106 -18322
rect 106 -15946 152 -15934
rect 106 -18322 112 -15946
rect 146 -18322 152 -15946
rect 106 -18334 152 -18322
rect -96 -18381 96 -18375
rect -96 -18415 -84 -18381
rect 84 -18415 96 -18381
rect -96 -18421 96 -18415
rect -96 -18489 96 -18483
rect -96 -18523 -84 -18489
rect 84 -18523 96 -18489
rect -96 -18529 96 -18523
rect -152 -18582 -106 -18570
rect -152 -20958 -146 -18582
rect -112 -20958 -106 -18582
rect -152 -20970 -106 -20958
rect 106 -18582 152 -18570
rect 106 -20958 112 -18582
rect 146 -20958 152 -18582
rect 106 -20970 152 -20958
rect -96 -21017 96 -21011
rect -96 -21051 -84 -21017
rect 84 -21051 96 -21017
rect -96 -21057 96 -21051
rect -96 -21125 96 -21119
rect -96 -21159 -84 -21125
rect 84 -21159 96 -21125
rect -96 -21165 96 -21159
rect -152 -21218 -106 -21206
rect -152 -23594 -146 -21218
rect -112 -23594 -106 -21218
rect -152 -23606 -106 -23594
rect 106 -21218 152 -21206
rect 106 -23594 112 -21218
rect 146 -23594 152 -21218
rect 106 -23606 152 -23594
rect -96 -23653 96 -23647
rect -96 -23687 -84 -23653
rect 84 -23687 96 -23653
rect -96 -23693 96 -23687
rect -96 -23761 96 -23755
rect -96 -23795 -84 -23761
rect 84 -23795 96 -23761
rect -96 -23801 96 -23795
rect -152 -23854 -106 -23842
rect -152 -26230 -146 -23854
rect -112 -26230 -106 -23854
rect -152 -26242 -106 -26230
rect 106 -23854 152 -23842
rect 106 -26230 112 -23854
rect 146 -26230 152 -23854
rect 106 -26242 152 -26230
rect -96 -26289 96 -26283
rect -96 -26323 -84 -26289
rect 84 -26323 96 -26289
rect -96 -26329 96 -26323
rect -96 -26397 96 -26391
rect -96 -26431 -84 -26397
rect 84 -26431 96 -26397
rect -96 -26437 96 -26431
rect -152 -26490 -106 -26478
rect -152 -28866 -146 -26490
rect -112 -28866 -106 -26490
rect -152 -28878 -106 -28866
rect 106 -26490 152 -26478
rect 106 -28866 112 -26490
rect 146 -28866 152 -26490
rect 106 -28878 152 -28866
rect -96 -28925 96 -28919
rect -96 -28959 -84 -28925
rect 84 -28959 96 -28925
rect -96 -28965 96 -28959
rect -96 -29033 96 -29027
rect -96 -29067 -84 -29033
rect 84 -29067 96 -29033
rect -96 -29073 96 -29067
rect -152 -29126 -106 -29114
rect -152 -31502 -146 -29126
rect -112 -31502 -106 -29126
rect -152 -31514 -106 -31502
rect 106 -29126 152 -29114
rect 106 -31502 112 -29126
rect 146 -31502 152 -29126
rect 106 -31514 152 -31502
rect -96 -31561 96 -31555
rect -96 -31595 -84 -31561
rect 84 -31595 96 -31561
rect -96 -31601 96 -31595
rect -96 -31669 96 -31663
rect -96 -31703 -84 -31669
rect 84 -31703 96 -31669
rect -96 -31709 96 -31703
rect -152 -31762 -106 -31750
rect -152 -34138 -146 -31762
rect -112 -34138 -106 -31762
rect -152 -34150 -106 -34138
rect 106 -31762 152 -31750
rect 106 -34138 112 -31762
rect 146 -34138 152 -31762
rect 106 -34150 152 -34138
rect -96 -34197 96 -34191
rect -96 -34231 -84 -34197
rect 84 -34231 96 -34197
rect -96 -34237 96 -34231
rect -96 -34305 96 -34299
rect -96 -34339 -84 -34305
rect 84 -34339 96 -34305
rect -96 -34345 96 -34339
rect -152 -34398 -106 -34386
rect -152 -36774 -146 -34398
rect -112 -36774 -106 -34398
rect -152 -36786 -106 -36774
rect 106 -34398 152 -34386
rect 106 -36774 112 -34398
rect 146 -36774 152 -34398
rect 106 -36786 152 -36774
rect -96 -36833 96 -36827
rect -96 -36867 -84 -36833
rect 84 -36867 96 -36833
rect -96 -36873 96 -36867
rect -96 -36941 96 -36935
rect -96 -36975 -84 -36941
rect 84 -36975 96 -36941
rect -96 -36981 96 -36975
rect -152 -37034 -106 -37022
rect -152 -39410 -146 -37034
rect -112 -39410 -106 -37034
rect -152 -39422 -106 -39410
rect 106 -37034 152 -37022
rect 106 -39410 112 -37034
rect 146 -39410 152 -37034
rect 106 -39422 152 -39410
rect -96 -39469 96 -39463
rect -96 -39503 -84 -39469
rect 84 -39503 96 -39469
rect -96 -39509 96 -39503
rect -96 -39577 96 -39571
rect -96 -39611 -84 -39577
rect 84 -39611 96 -39577
rect -96 -39617 96 -39611
rect -152 -39670 -106 -39658
rect -152 -42046 -146 -39670
rect -112 -42046 -106 -39670
rect -152 -42058 -106 -42046
rect 106 -39670 152 -39658
rect 106 -42046 112 -39670
rect 146 -42046 152 -39670
rect 106 -42058 152 -42046
rect -96 -42105 96 -42099
rect -96 -42139 -84 -42105
rect 84 -42139 96 -42105
rect -96 -42145 96 -42139
rect -96 -42213 96 -42207
rect -96 -42247 -84 -42213
rect 84 -42247 96 -42213
rect -96 -42253 96 -42247
rect -152 -42306 -106 -42294
rect -152 -44682 -146 -42306
rect -112 -44682 -106 -42306
rect -152 -44694 -106 -44682
rect 106 -42306 152 -42294
rect 106 -44682 112 -42306
rect 146 -44682 152 -42306
rect 106 -44694 152 -44682
rect -96 -44741 96 -44735
rect -96 -44775 -84 -44741
rect 84 -44775 96 -44741
rect -96 -44781 96 -44775
rect -96 -44849 96 -44843
rect -96 -44883 -84 -44849
rect 84 -44883 96 -44849
rect -96 -44889 96 -44883
rect -152 -44942 -106 -44930
rect -152 -47318 -146 -44942
rect -112 -47318 -106 -44942
rect -152 -47330 -106 -47318
rect 106 -44942 152 -44930
rect 106 -47318 112 -44942
rect 146 -47318 152 -44942
rect 106 -47330 152 -47318
rect -96 -47377 96 -47371
rect -96 -47411 -84 -47377
rect 84 -47411 96 -47377
rect -96 -47417 96 -47411
rect -96 -47485 96 -47479
rect -96 -47519 -84 -47485
rect 84 -47519 96 -47485
rect -96 -47525 96 -47519
rect -152 -47578 -106 -47566
rect -152 -49954 -146 -47578
rect -112 -49954 -106 -47578
rect -152 -49966 -106 -49954
rect 106 -47578 152 -47566
rect 106 -49954 112 -47578
rect 146 -49954 152 -47578
rect 106 -49966 152 -49954
rect -96 -50013 96 -50007
rect -96 -50047 -84 -50013
rect 84 -50047 96 -50013
rect -96 -50053 96 -50047
rect -96 -50121 96 -50115
rect -96 -50155 -84 -50121
rect 84 -50155 96 -50121
rect -96 -50161 96 -50155
rect -152 -50214 -106 -50202
rect -152 -52590 -146 -50214
rect -112 -52590 -106 -50214
rect -152 -52602 -106 -52590
rect 106 -50214 152 -50202
rect 106 -52590 112 -50214
rect 146 -52590 152 -50214
rect 106 -52602 152 -52590
rect -96 -52649 96 -52643
rect -96 -52683 -84 -52649
rect 84 -52683 96 -52649
rect -96 -52689 96 -52683
rect -96 -52757 96 -52751
rect -96 -52791 -84 -52757
rect 84 -52791 96 -52757
rect -96 -52797 96 -52791
rect -152 -52850 -106 -52838
rect -152 -55226 -146 -52850
rect -112 -55226 -106 -52850
rect -152 -55238 -106 -55226
rect 106 -52850 152 -52838
rect 106 -55226 112 -52850
rect 146 -55226 152 -52850
rect 106 -55238 152 -55226
rect -96 -55285 96 -55279
rect -96 -55319 -84 -55285
rect 84 -55319 96 -55285
rect -96 -55325 96 -55319
rect -96 -55393 96 -55387
rect -96 -55427 -84 -55393
rect 84 -55427 96 -55393
rect -96 -55433 96 -55427
rect -152 -55486 -106 -55474
rect -152 -57862 -146 -55486
rect -112 -57862 -106 -55486
rect -152 -57874 -106 -57862
rect 106 -55486 152 -55474
rect 106 -57862 112 -55486
rect 146 -57862 152 -55486
rect 106 -57874 152 -57862
rect -96 -57921 96 -57915
rect -96 -57955 -84 -57921
rect 84 -57955 96 -57921
rect -96 -57961 96 -57955
rect -96 -58029 96 -58023
rect -96 -58063 -84 -58029
rect 84 -58063 96 -58029
rect -96 -58069 96 -58063
rect -152 -58122 -106 -58110
rect -152 -60498 -146 -58122
rect -112 -60498 -106 -58122
rect -152 -60510 -106 -60498
rect 106 -58122 152 -58110
rect 106 -60498 112 -58122
rect 146 -60498 152 -58122
rect 106 -60510 152 -60498
rect -96 -60557 96 -60551
rect -96 -60591 -84 -60557
rect 84 -60591 96 -60557
rect -96 -60597 96 -60591
rect -96 -60665 96 -60659
rect -96 -60699 -84 -60665
rect 84 -60699 96 -60665
rect -96 -60705 96 -60699
rect -152 -60758 -106 -60746
rect -152 -63134 -146 -60758
rect -112 -63134 -106 -60758
rect -152 -63146 -106 -63134
rect 106 -60758 152 -60746
rect 106 -63134 112 -60758
rect 146 -63134 152 -60758
rect 106 -63146 152 -63134
rect -96 -63193 96 -63187
rect -96 -63227 -84 -63193
rect 84 -63227 96 -63193
rect -96 -63233 96 -63227
rect -96 -63301 96 -63295
rect -96 -63335 -84 -63301
rect 84 -63335 96 -63301
rect -96 -63341 96 -63335
rect -152 -63394 -106 -63382
rect -152 -65770 -146 -63394
rect -112 -65770 -106 -63394
rect -152 -65782 -106 -65770
rect 106 -63394 152 -63382
rect 106 -65770 112 -63394
rect 146 -65770 152 -63394
rect 106 -65782 152 -65770
rect -96 -65829 96 -65823
rect -96 -65863 -84 -65829
rect 84 -65863 96 -65829
rect -96 -65869 96 -65863
rect -96 -65937 96 -65931
rect -96 -65971 -84 -65937
rect 84 -65971 96 -65937
rect -96 -65977 96 -65971
rect -152 -66030 -106 -66018
rect -152 -68406 -146 -66030
rect -112 -68406 -106 -66030
rect -152 -68418 -106 -68406
rect 106 -66030 152 -66018
rect 106 -68406 112 -66030
rect 146 -68406 152 -66030
rect 106 -68418 152 -68406
rect -96 -68465 96 -68459
rect -96 -68499 -84 -68465
rect 84 -68499 96 -68465
rect -96 -68505 96 -68499
rect -96 -68573 96 -68567
rect -96 -68607 -84 -68573
rect 84 -68607 96 -68573
rect -96 -68613 96 -68607
rect -152 -68666 -106 -68654
rect -152 -71042 -146 -68666
rect -112 -71042 -106 -68666
rect -152 -71054 -106 -71042
rect 106 -68666 152 -68654
rect 106 -71042 112 -68666
rect 146 -71042 152 -68666
rect 106 -71054 152 -71042
rect -96 -71101 96 -71095
rect -96 -71135 -84 -71101
rect 84 -71135 96 -71101
rect -96 -71141 96 -71135
rect -96 -71209 96 -71203
rect -96 -71243 -84 -71209
rect 84 -71243 96 -71209
rect -96 -71249 96 -71243
rect -152 -71302 -106 -71290
rect -152 -73678 -146 -71302
rect -112 -73678 -106 -71302
rect -152 -73690 -106 -73678
rect 106 -71302 152 -71290
rect 106 -73678 112 -71302
rect 146 -73678 152 -71302
rect 106 -73690 152 -73678
rect -96 -73737 96 -73731
rect -96 -73771 -84 -73737
rect 84 -73771 96 -73737
rect -96 -73777 96 -73771
rect -96 -73845 96 -73839
rect -96 -73879 -84 -73845
rect 84 -73879 96 -73845
rect -96 -73885 96 -73879
rect -152 -73938 -106 -73926
rect -152 -76314 -146 -73938
rect -112 -76314 -106 -73938
rect -152 -76326 -106 -76314
rect 106 -73938 152 -73926
rect 106 -76314 112 -73938
rect 146 -76314 152 -73938
rect 106 -76326 152 -76314
rect -96 -76373 96 -76367
rect -96 -76407 -84 -76373
rect 84 -76407 96 -76373
rect -96 -76413 96 -76407
rect -96 -76481 96 -76475
rect -96 -76515 -84 -76481
rect 84 -76515 96 -76481
rect -96 -76521 96 -76515
rect -152 -76574 -106 -76562
rect -152 -78950 -146 -76574
rect -112 -78950 -106 -76574
rect -152 -78962 -106 -78950
rect 106 -76574 152 -76562
rect 106 -78950 112 -76574
rect 146 -78950 152 -76574
rect 106 -78962 152 -78950
rect -96 -79009 96 -79003
rect -96 -79043 -84 -79009
rect 84 -79043 96 -79009
rect -96 -79049 96 -79043
rect -96 -79117 96 -79111
rect -96 -79151 -84 -79117
rect 84 -79151 96 -79117
rect -96 -79157 96 -79151
rect -152 -79210 -106 -79198
rect -152 -81586 -146 -79210
rect -112 -81586 -106 -79210
rect -152 -81598 -106 -81586
rect 106 -79210 152 -79198
rect 106 -81586 112 -79210
rect 146 -81586 152 -79210
rect 106 -81598 152 -81586
rect -96 -81645 96 -81639
rect -96 -81679 -84 -81645
rect 84 -81679 96 -81645
rect -96 -81685 96 -81679
rect -96 -81753 96 -81747
rect -96 -81787 -84 -81753
rect 84 -81787 96 -81753
rect -96 -81793 96 -81787
rect -152 -81846 -106 -81834
rect -152 -84222 -146 -81846
rect -112 -84222 -106 -81846
rect -152 -84234 -106 -84222
rect 106 -81846 152 -81834
rect 106 -84222 112 -81846
rect 146 -84222 152 -81846
rect 106 -84234 152 -84222
rect -96 -84281 96 -84275
rect -96 -84315 -84 -84281
rect 84 -84315 96 -84281
rect -96 -84321 96 -84315
rect -96 -84389 96 -84383
rect -96 -84423 -84 -84389
rect 84 -84423 96 -84389
rect -96 -84429 96 -84423
rect -152 -84482 -106 -84470
rect -152 -86858 -146 -84482
rect -112 -86858 -106 -84482
rect -152 -86870 -106 -86858
rect 106 -84482 152 -84470
rect 106 -86858 112 -84482
rect 146 -86858 152 -84482
rect 106 -86870 152 -86858
rect -96 -86917 96 -86911
rect -96 -86951 -84 -86917
rect 84 -86951 96 -86917
rect -96 -86957 96 -86951
rect -96 -87025 96 -87019
rect -96 -87059 -84 -87025
rect 84 -87059 96 -87025
rect -96 -87065 96 -87059
rect -152 -87118 -106 -87106
rect -152 -89494 -146 -87118
rect -112 -89494 -106 -87118
rect -152 -89506 -106 -89494
rect 106 -87118 152 -87106
rect 106 -89494 112 -87118
rect 146 -89494 152 -87118
rect 106 -89506 152 -89494
rect -96 -89553 96 -89547
rect -96 -89587 -84 -89553
rect 84 -89587 96 -89553
rect -96 -89593 96 -89587
rect -96 -89661 96 -89655
rect -96 -89695 -84 -89661
rect 84 -89695 96 -89661
rect -96 -89701 96 -89695
rect -152 -89754 -106 -89742
rect -152 -92130 -146 -89754
rect -112 -92130 -106 -89754
rect -152 -92142 -106 -92130
rect 106 -89754 152 -89742
rect 106 -92130 112 -89754
rect 146 -92130 152 -89754
rect 106 -92142 152 -92130
rect -96 -92189 96 -92183
rect -96 -92223 -84 -92189
rect 84 -92223 96 -92189
rect -96 -92229 96 -92223
rect -96 -92297 96 -92291
rect -96 -92331 -84 -92297
rect 84 -92331 96 -92297
rect -96 -92337 96 -92331
rect -152 -92390 -106 -92378
rect -152 -94766 -146 -92390
rect -112 -94766 -106 -92390
rect -152 -94778 -106 -94766
rect 106 -92390 152 -92378
rect 106 -94766 112 -92390
rect 146 -94766 152 -92390
rect 106 -94778 152 -94766
rect -96 -94825 96 -94819
rect -96 -94859 -84 -94825
rect 84 -94859 96 -94825
rect -96 -94865 96 -94859
rect -96 -94933 96 -94927
rect -96 -94967 -84 -94933
rect 84 -94967 96 -94933
rect -96 -94973 96 -94967
rect -152 -95026 -106 -95014
rect -152 -97402 -146 -95026
rect -112 -97402 -106 -95026
rect -152 -97414 -106 -97402
rect 106 -95026 152 -95014
rect 106 -97402 112 -95026
rect 146 -97402 152 -95026
rect 106 -97414 152 -97402
rect -96 -97461 96 -97455
rect -96 -97495 -84 -97461
rect 84 -97495 96 -97461
rect -96 -97501 96 -97495
rect -96 -97569 96 -97563
rect -96 -97603 -84 -97569
rect 84 -97603 96 -97569
rect -96 -97609 96 -97603
rect -152 -97662 -106 -97650
rect -152 -100038 -146 -97662
rect -112 -100038 -106 -97662
rect -152 -100050 -106 -100038
rect 106 -97662 152 -97650
rect 106 -100038 112 -97662
rect 146 -100038 152 -97662
rect 106 -100050 152 -100038
rect -96 -100097 96 -100091
rect -96 -100131 -84 -100097
rect 84 -100131 96 -100097
rect -96 -100137 96 -100131
rect -96 -100205 96 -100199
rect -96 -100239 -84 -100205
rect 84 -100239 96 -100205
rect -96 -100245 96 -100239
rect -152 -100298 -106 -100286
rect -152 -102674 -146 -100298
rect -112 -102674 -106 -100298
rect -152 -102686 -106 -102674
rect 106 -100298 152 -100286
rect 106 -102674 112 -100298
rect 146 -102674 152 -100298
rect 106 -102686 152 -102674
rect -96 -102733 96 -102727
rect -96 -102767 -84 -102733
rect 84 -102767 96 -102733
rect -96 -102773 96 -102767
rect -96 -102841 96 -102835
rect -96 -102875 -84 -102841
rect 84 -102875 96 -102841
rect -96 -102881 96 -102875
rect -152 -102934 -106 -102922
rect -152 -105310 -146 -102934
rect -112 -105310 -106 -102934
rect -152 -105322 -106 -105310
rect 106 -102934 152 -102922
rect 106 -105310 112 -102934
rect 146 -105310 152 -102934
rect 106 -105322 152 -105310
rect -96 -105369 96 -105363
rect -96 -105403 -84 -105369
rect 84 -105403 96 -105369
rect -96 -105409 96 -105403
rect -96 -105477 96 -105471
rect -96 -105511 -84 -105477
rect 84 -105511 96 -105477
rect -96 -105517 96 -105511
rect -152 -105570 -106 -105558
rect -152 -107946 -146 -105570
rect -112 -107946 -106 -105570
rect -152 -107958 -106 -107946
rect 106 -105570 152 -105558
rect 106 -107946 112 -105570
rect 146 -107946 152 -105570
rect 106 -107958 152 -107946
rect -96 -108005 96 -107999
rect -96 -108039 -84 -108005
rect 84 -108039 96 -108005
rect -96 -108045 96 -108039
rect -96 -108113 96 -108107
rect -96 -108147 -84 -108113
rect 84 -108147 96 -108113
rect -96 -108153 96 -108147
rect -152 -108206 -106 -108194
rect -152 -110582 -146 -108206
rect -112 -110582 -106 -108206
rect -152 -110594 -106 -110582
rect 106 -108206 152 -108194
rect 106 -110582 112 -108206
rect 146 -110582 152 -108206
rect 106 -110594 152 -110582
rect -96 -110641 96 -110635
rect -96 -110675 -84 -110641
rect 84 -110675 96 -110641
rect -96 -110681 96 -110675
rect -96 -110749 96 -110743
rect -96 -110783 -84 -110749
rect 84 -110783 96 -110749
rect -96 -110789 96 -110783
rect -152 -110842 -106 -110830
rect -152 -113218 -146 -110842
rect -112 -113218 -106 -110842
rect -152 -113230 -106 -113218
rect 106 -110842 152 -110830
rect 106 -113218 112 -110842
rect 146 -113218 152 -110842
rect 106 -113230 152 -113218
rect -96 -113277 96 -113271
rect -96 -113311 -84 -113277
rect 84 -113311 96 -113277
rect -96 -113317 96 -113311
rect -96 -113385 96 -113379
rect -96 -113419 -84 -113385
rect 84 -113419 96 -113385
rect -96 -113425 96 -113419
rect -152 -113478 -106 -113466
rect -152 -115854 -146 -113478
rect -112 -115854 -106 -113478
rect -152 -115866 -106 -115854
rect 106 -113478 152 -113466
rect 106 -115854 112 -113478
rect 146 -115854 152 -113478
rect 106 -115866 152 -115854
rect -96 -115913 96 -115907
rect -96 -115947 -84 -115913
rect 84 -115947 96 -115913
rect -96 -115953 96 -115947
rect -96 -116021 96 -116015
rect -96 -116055 -84 -116021
rect 84 -116055 96 -116021
rect -96 -116061 96 -116055
rect -152 -116114 -106 -116102
rect -152 -118490 -146 -116114
rect -112 -118490 -106 -116114
rect -152 -118502 -106 -118490
rect 106 -116114 152 -116102
rect 106 -118490 112 -116114
rect 146 -118490 152 -116114
rect 106 -118502 152 -118490
rect -96 -118549 96 -118543
rect -96 -118583 -84 -118549
rect 84 -118583 96 -118549
rect -96 -118589 96 -118583
rect -96 -118657 96 -118651
rect -96 -118691 -84 -118657
rect 84 -118691 96 -118657
rect -96 -118697 96 -118691
rect -152 -118750 -106 -118738
rect -152 -121126 -146 -118750
rect -112 -121126 -106 -118750
rect -152 -121138 -106 -121126
rect 106 -118750 152 -118738
rect 106 -121126 112 -118750
rect 146 -121126 152 -118750
rect 106 -121138 152 -121126
rect -96 -121185 96 -121179
rect -96 -121219 -84 -121185
rect 84 -121219 96 -121185
rect -96 -121225 96 -121219
rect -96 -121293 96 -121287
rect -96 -121327 -84 -121293
rect 84 -121327 96 -121293
rect -96 -121333 96 -121327
rect -152 -121386 -106 -121374
rect -152 -123762 -146 -121386
rect -112 -123762 -106 -121386
rect -152 -123774 -106 -123762
rect 106 -121386 152 -121374
rect 106 -123762 112 -121386
rect 146 -123762 152 -121386
rect 106 -123774 152 -123762
rect -96 -123821 96 -123815
rect -96 -123855 -84 -123821
rect 84 -123855 96 -123821
rect -96 -123861 96 -123855
rect -96 -123929 96 -123923
rect -96 -123963 -84 -123929
rect 84 -123963 96 -123929
rect -96 -123969 96 -123963
rect -152 -124022 -106 -124010
rect -152 -126398 -146 -124022
rect -112 -126398 -106 -124022
rect -152 -126410 -106 -126398
rect 106 -124022 152 -124010
rect 106 -126398 112 -124022
rect 146 -126398 152 -124022
rect 106 -126410 152 -126398
rect -96 -126457 96 -126451
rect -96 -126491 -84 -126457
rect 84 -126491 96 -126457
rect -96 -126497 96 -126491
rect -96 -126565 96 -126559
rect -96 -126599 -84 -126565
rect 84 -126599 96 -126565
rect -96 -126605 96 -126599
rect -152 -126658 -106 -126646
rect -152 -129034 -146 -126658
rect -112 -129034 -106 -126658
rect -152 -129046 -106 -129034
rect 106 -126658 152 -126646
rect 106 -129034 112 -126658
rect 146 -129034 152 -126658
rect 106 -129046 152 -129034
rect -96 -129093 96 -129087
rect -96 -129127 -84 -129093
rect 84 -129127 96 -129093
rect -96 -129133 96 -129127
rect -96 -129201 96 -129195
rect -96 -129235 -84 -129201
rect 84 -129235 96 -129201
rect -96 -129241 96 -129235
rect -152 -129294 -106 -129282
rect -152 -131670 -146 -129294
rect -112 -131670 -106 -129294
rect -152 -131682 -106 -131670
rect 106 -129294 152 -129282
rect 106 -131670 112 -129294
rect 146 -131670 152 -129294
rect 106 -131682 152 -131670
rect -96 -131729 96 -131723
rect -96 -131763 -84 -131729
rect 84 -131763 96 -131729
rect -96 -131769 96 -131763
rect -96 -131837 96 -131831
rect -96 -131871 -84 -131837
rect 84 -131871 96 -131837
rect -96 -131877 96 -131871
rect -152 -131930 -106 -131918
rect -152 -134306 -146 -131930
rect -112 -134306 -106 -131930
rect -152 -134318 -106 -134306
rect 106 -131930 152 -131918
rect 106 -134306 112 -131930
rect 146 -134306 152 -131930
rect 106 -134318 152 -134306
rect -96 -134365 96 -134359
rect -96 -134399 -84 -134365
rect 84 -134399 96 -134365
rect -96 -134405 96 -134399
rect -96 -134473 96 -134467
rect -96 -134507 -84 -134473
rect 84 -134507 96 -134473
rect -96 -134513 96 -134507
rect -152 -134566 -106 -134554
rect -152 -136942 -146 -134566
rect -112 -136942 -106 -134566
rect -152 -136954 -106 -136942
rect 106 -134566 152 -134554
rect 106 -136942 112 -134566
rect 146 -136942 152 -134566
rect 106 -136954 152 -136942
rect -96 -137001 96 -136995
rect -96 -137035 -84 -137001
rect 84 -137035 96 -137001
rect -96 -137041 96 -137035
rect -96 -137109 96 -137103
rect -96 -137143 -84 -137109
rect 84 -137143 96 -137109
rect -96 -137149 96 -137143
rect -152 -137202 -106 -137190
rect -152 -139578 -146 -137202
rect -112 -139578 -106 -137202
rect -152 -139590 -106 -139578
rect 106 -137202 152 -137190
rect 106 -139578 112 -137202
rect 146 -139578 152 -137202
rect 106 -139590 152 -139578
rect -96 -139637 96 -139631
rect -96 -139671 -84 -139637
rect 84 -139671 96 -139637
rect -96 -139677 96 -139671
rect -96 -139745 96 -139739
rect -96 -139779 -84 -139745
rect 84 -139779 96 -139745
rect -96 -139785 96 -139779
rect -152 -139838 -106 -139826
rect -152 -142214 -146 -139838
rect -112 -142214 -106 -139838
rect -152 -142226 -106 -142214
rect 106 -139838 152 -139826
rect 106 -142214 112 -139838
rect 146 -142214 152 -139838
rect 106 -142226 152 -142214
rect -96 -142273 96 -142267
rect -96 -142307 -84 -142273
rect 84 -142307 96 -142273
rect -96 -142313 96 -142307
rect -96 -142381 96 -142375
rect -96 -142415 -84 -142381
rect 84 -142415 96 -142381
rect -96 -142421 96 -142415
rect -152 -142474 -106 -142462
rect -152 -144850 -146 -142474
rect -112 -144850 -106 -142474
rect -152 -144862 -106 -144850
rect 106 -142474 152 -142462
rect 106 -144850 112 -142474
rect 146 -144850 152 -142474
rect 106 -144862 152 -144850
rect -96 -144909 96 -144903
rect -96 -144943 -84 -144909
rect 84 -144943 96 -144909
rect -96 -144949 96 -144943
rect -96 -145017 96 -145011
rect -96 -145051 -84 -145017
rect 84 -145051 96 -145017
rect -96 -145057 96 -145051
rect -152 -145110 -106 -145098
rect -152 -147486 -146 -145110
rect -112 -147486 -106 -145110
rect -152 -147498 -106 -147486
rect 106 -145110 152 -145098
rect 106 -147486 112 -145110
rect 146 -147486 152 -145110
rect 106 -147498 152 -147486
rect -96 -147545 96 -147539
rect -96 -147579 -84 -147545
rect 84 -147579 96 -147545
rect -96 -147585 96 -147579
rect -96 -147653 96 -147647
rect -96 -147687 -84 -147653
rect 84 -147687 96 -147653
rect -96 -147693 96 -147687
rect -152 -147746 -106 -147734
rect -152 -150122 -146 -147746
rect -112 -150122 -106 -147746
rect -152 -150134 -106 -150122
rect 106 -147746 152 -147734
rect 106 -150122 112 -147746
rect 146 -150122 152 -147746
rect 106 -150134 152 -150122
rect -96 -150181 96 -150175
rect -96 -150215 -84 -150181
rect 84 -150215 96 -150181
rect -96 -150221 96 -150215
rect -96 -150289 96 -150283
rect -96 -150323 -84 -150289
rect 84 -150323 96 -150289
rect -96 -150329 96 -150323
rect -152 -150382 -106 -150370
rect -152 -152758 -146 -150382
rect -112 -152758 -106 -150382
rect -152 -152770 -106 -152758
rect 106 -150382 152 -150370
rect 106 -152758 112 -150382
rect 146 -152758 152 -150382
rect 106 -152770 152 -152758
rect -96 -152817 96 -152811
rect -96 -152851 -84 -152817
rect 84 -152851 96 -152817
rect -96 -152857 96 -152851
rect -96 -152925 96 -152919
rect -96 -152959 -84 -152925
rect 84 -152959 96 -152925
rect -96 -152965 96 -152959
rect -152 -153018 -106 -153006
rect -152 -155394 -146 -153018
rect -112 -155394 -106 -153018
rect -152 -155406 -106 -155394
rect 106 -153018 152 -153006
rect 106 -155394 112 -153018
rect 146 -155394 152 -153018
rect 106 -155406 152 -155394
rect -96 -155453 96 -155447
rect -96 -155487 -84 -155453
rect 84 -155487 96 -155453
rect -96 -155493 96 -155487
rect -96 -155561 96 -155555
rect -96 -155595 -84 -155561
rect 84 -155595 96 -155561
rect -96 -155601 96 -155595
rect -152 -155654 -106 -155642
rect -152 -158030 -146 -155654
rect -112 -158030 -106 -155654
rect -152 -158042 -106 -158030
rect 106 -155654 152 -155642
rect 106 -158030 112 -155654
rect 146 -158030 152 -155654
rect 106 -158042 152 -158030
rect -96 -158089 96 -158083
rect -96 -158123 -84 -158089
rect 84 -158123 96 -158089
rect -96 -158129 96 -158123
rect -96 -158197 96 -158191
rect -96 -158231 -84 -158197
rect 84 -158231 96 -158197
rect -96 -158237 96 -158231
rect -152 -158290 -106 -158278
rect -152 -160666 -146 -158290
rect -112 -160666 -106 -158290
rect -152 -160678 -106 -160666
rect 106 -158290 152 -158278
rect 106 -160666 112 -158290
rect 146 -160666 152 -158290
rect 106 -160678 152 -160666
rect -96 -160725 96 -160719
rect -96 -160759 -84 -160725
rect 84 -160759 96 -160725
rect -96 -160765 96 -160759
rect -96 -160833 96 -160827
rect -96 -160867 -84 -160833
rect 84 -160867 96 -160833
rect -96 -160873 96 -160867
rect -152 -160926 -106 -160914
rect -152 -163302 -146 -160926
rect -112 -163302 -106 -160926
rect -152 -163314 -106 -163302
rect 106 -160926 152 -160914
rect 106 -163302 112 -160926
rect 146 -163302 152 -160926
rect 106 -163314 152 -163302
rect -96 -163361 96 -163355
rect -96 -163395 -84 -163361
rect 84 -163395 96 -163361
rect -96 -163401 96 -163395
rect -96 -163469 96 -163463
rect -96 -163503 -84 -163469
rect 84 -163503 96 -163469
rect -96 -163509 96 -163503
rect -152 -163562 -106 -163550
rect -152 -165938 -146 -163562
rect -112 -165938 -106 -163562
rect -152 -165950 -106 -165938
rect 106 -163562 152 -163550
rect 106 -165938 112 -163562
rect 146 -165938 152 -163562
rect 106 -165950 152 -165938
rect -96 -165997 96 -165991
rect -96 -166031 -84 -165997
rect 84 -166031 96 -165997
rect -96 -166037 96 -166031
rect -96 -166105 96 -166099
rect -96 -166139 -84 -166105
rect 84 -166139 96 -166105
rect -96 -166145 96 -166139
rect -152 -166198 -106 -166186
rect -152 -168574 -146 -166198
rect -112 -168574 -106 -166198
rect -152 -168586 -106 -168574
rect 106 -166198 152 -166186
rect 106 -168574 112 -166198
rect 146 -168574 152 -166198
rect 106 -168586 152 -168574
rect -96 -168633 96 -168627
rect -96 -168667 -84 -168633
rect 84 -168667 96 -168633
rect -96 -168673 96 -168667
rect -96 -168741 96 -168735
rect -96 -168775 -84 -168741
rect 84 -168775 96 -168741
rect -96 -168781 96 -168775
rect -152 -168834 -106 -168822
rect -152 -171210 -146 -168834
rect -112 -171210 -106 -168834
rect -152 -171222 -106 -171210
rect 106 -168834 152 -168822
rect 106 -171210 112 -168834
rect 146 -171210 152 -168834
rect 106 -171222 152 -171210
rect -96 -171269 96 -171263
rect -96 -171303 -84 -171269
rect 84 -171303 96 -171269
rect -96 -171309 96 -171303
rect -96 -171377 96 -171371
rect -96 -171411 -84 -171377
rect 84 -171411 96 -171377
rect -96 -171417 96 -171411
rect -152 -171470 -106 -171458
rect -152 -173846 -146 -171470
rect -112 -173846 -106 -171470
rect -152 -173858 -106 -173846
rect 106 -171470 152 -171458
rect 106 -173846 112 -171470
rect 146 -173846 152 -171470
rect 106 -173858 152 -173846
rect -96 -173905 96 -173899
rect -96 -173939 -84 -173905
rect 84 -173939 96 -173905
rect -96 -173945 96 -173939
rect -96 -174013 96 -174007
rect -96 -174047 -84 -174013
rect 84 -174047 96 -174013
rect -96 -174053 96 -174047
rect -152 -174106 -106 -174094
rect -152 -176482 -146 -174106
rect -112 -176482 -106 -174106
rect -152 -176494 -106 -176482
rect 106 -174106 152 -174094
rect 106 -176482 112 -174106
rect 146 -176482 152 -174106
rect 106 -176494 152 -176482
rect -96 -176541 96 -176535
rect -96 -176575 -84 -176541
rect 84 -176575 96 -176541
rect -96 -176581 96 -176575
rect -96 -176649 96 -176643
rect -96 -176683 -84 -176649
rect 84 -176683 96 -176649
rect -96 -176689 96 -176683
rect -152 -176742 -106 -176730
rect -152 -179118 -146 -176742
rect -112 -179118 -106 -176742
rect -152 -179130 -106 -179118
rect 106 -176742 152 -176730
rect 106 -179118 112 -176742
rect 146 -179118 152 -176742
rect 106 -179130 152 -179118
rect -96 -179177 96 -179171
rect -96 -179211 -84 -179177
rect 84 -179211 96 -179177
rect -96 -179217 96 -179211
rect -96 -179285 96 -179279
rect -96 -179319 -84 -179285
rect 84 -179319 96 -179285
rect -96 -179325 96 -179319
rect -152 -179378 -106 -179366
rect -152 -181754 -146 -179378
rect -112 -181754 -106 -179378
rect -152 -181766 -106 -181754
rect 106 -179378 152 -179366
rect 106 -181754 112 -179378
rect 146 -181754 152 -179378
rect 106 -181766 152 -181754
rect -96 -181813 96 -181807
rect -96 -181847 -84 -181813
rect 84 -181847 96 -181813
rect -96 -181853 96 -181847
rect -96 -181921 96 -181915
rect -96 -181955 -84 -181921
rect 84 -181955 96 -181921
rect -96 -181961 96 -181955
rect -152 -182014 -106 -182002
rect -152 -184390 -146 -182014
rect -112 -184390 -106 -182014
rect -152 -184402 -106 -184390
rect 106 -182014 152 -182002
rect 106 -184390 112 -182014
rect 146 -184390 152 -182014
rect 106 -184402 152 -184390
rect -96 -184449 96 -184443
rect -96 -184483 -84 -184449
rect 84 -184483 96 -184449
rect -96 -184489 96 -184483
rect -96 -184557 96 -184551
rect -96 -184591 -84 -184557
rect 84 -184591 96 -184557
rect -96 -184597 96 -184591
rect -152 -184650 -106 -184638
rect -152 -187026 -146 -184650
rect -112 -187026 -106 -184650
rect -152 -187038 -106 -187026
rect 106 -184650 152 -184638
rect 106 -187026 112 -184650
rect 146 -187026 152 -184650
rect 106 -187038 152 -187026
rect -96 -187085 96 -187079
rect -96 -187119 -84 -187085
rect 84 -187119 96 -187085
rect -96 -187125 96 -187119
rect -96 -187193 96 -187187
rect -96 -187227 -84 -187193
rect 84 -187227 96 -187193
rect -96 -187233 96 -187227
rect -152 -187286 -106 -187274
rect -152 -189662 -146 -187286
rect -112 -189662 -106 -187286
rect -152 -189674 -106 -189662
rect 106 -187286 152 -187274
rect 106 -189662 112 -187286
rect 146 -189662 152 -187286
rect 106 -189674 152 -189662
rect -96 -189721 96 -189715
rect -96 -189755 -84 -189721
rect 84 -189755 96 -189721
rect -96 -189761 96 -189755
rect -96 -189829 96 -189823
rect -96 -189863 -84 -189829
rect 84 -189863 96 -189829
rect -96 -189869 96 -189863
rect -152 -189922 -106 -189910
rect -152 -192298 -146 -189922
rect -112 -192298 -106 -189922
rect -152 -192310 -106 -192298
rect 106 -189922 152 -189910
rect 106 -192298 112 -189922
rect 146 -192298 152 -189922
rect 106 -192310 152 -192298
rect -96 -192357 96 -192351
rect -96 -192391 -84 -192357
rect 84 -192391 96 -192357
rect -96 -192397 96 -192391
rect -96 -192465 96 -192459
rect -96 -192499 -84 -192465
rect 84 -192499 96 -192465
rect -96 -192505 96 -192499
rect -152 -192558 -106 -192546
rect -152 -194934 -146 -192558
rect -112 -194934 -106 -192558
rect -152 -194946 -106 -194934
rect 106 -192558 152 -192546
rect 106 -194934 112 -192558
rect 146 -194934 152 -192558
rect 106 -194946 152 -194934
rect -96 -194993 96 -194987
rect -96 -195027 -84 -194993
rect 84 -195027 96 -194993
rect -96 -195033 96 -195027
rect -96 -195101 96 -195095
rect -96 -195135 -84 -195101
rect 84 -195135 96 -195101
rect -96 -195141 96 -195135
rect -152 -195194 -106 -195182
rect -152 -197570 -146 -195194
rect -112 -197570 -106 -195194
rect -152 -197582 -106 -197570
rect 106 -195194 152 -195182
rect 106 -197570 112 -195194
rect 146 -197570 152 -195194
rect 106 -197582 152 -197570
rect -96 -197629 96 -197623
rect -96 -197663 -84 -197629
rect 84 -197663 96 -197629
rect -96 -197669 96 -197663
rect -96 -197737 96 -197731
rect -96 -197771 -84 -197737
rect 84 -197771 96 -197737
rect -96 -197777 96 -197771
rect -152 -197830 -106 -197818
rect -152 -200206 -146 -197830
rect -112 -200206 -106 -197830
rect -152 -200218 -106 -200206
rect 106 -197830 152 -197818
rect 106 -200206 112 -197830
rect 146 -200206 152 -197830
rect 106 -200218 152 -200206
rect -96 -200265 96 -200259
rect -96 -200299 -84 -200265
rect 84 -200299 96 -200265
rect -96 -200305 96 -200299
rect -96 -200373 96 -200367
rect -96 -200407 -84 -200373
rect 84 -200407 96 -200373
rect -96 -200413 96 -200407
rect -152 -200466 -106 -200454
rect -152 -202842 -146 -200466
rect -112 -202842 -106 -200466
rect -152 -202854 -106 -202842
rect 106 -200466 152 -200454
rect 106 -202842 112 -200466
rect 146 -202842 152 -200466
rect 106 -202854 152 -202842
rect -96 -202901 96 -202895
rect -96 -202935 -84 -202901
rect 84 -202935 96 -202901
rect -96 -202941 96 -202935
rect -96 -203009 96 -203003
rect -96 -203043 -84 -203009
rect 84 -203043 96 -203009
rect -96 -203049 96 -203043
rect -152 -203102 -106 -203090
rect -152 -205478 -146 -203102
rect -112 -205478 -106 -203102
rect -152 -205490 -106 -205478
rect 106 -203102 152 -203090
rect 106 -205478 112 -203102
rect 146 -205478 152 -203102
rect 106 -205490 152 -205478
rect -96 -205537 96 -205531
rect -96 -205571 -84 -205537
rect 84 -205571 96 -205537
rect -96 -205577 96 -205571
rect -96 -205645 96 -205639
rect -96 -205679 -84 -205645
rect 84 -205679 96 -205645
rect -96 -205685 96 -205679
rect -152 -205738 -106 -205726
rect -152 -208114 -146 -205738
rect -112 -208114 -106 -205738
rect -152 -208126 -106 -208114
rect 106 -205738 152 -205726
rect 106 -208114 112 -205738
rect 146 -208114 152 -205738
rect 106 -208126 152 -208114
rect -96 -208173 96 -208167
rect -96 -208207 -84 -208173
rect 84 -208207 96 -208173
rect -96 -208213 96 -208207
rect -96 -208281 96 -208275
rect -96 -208315 -84 -208281
rect 84 -208315 96 -208281
rect -96 -208321 96 -208315
rect -152 -208374 -106 -208362
rect -152 -210750 -146 -208374
rect -112 -210750 -106 -208374
rect -152 -210762 -106 -210750
rect 106 -208374 152 -208362
rect 106 -210750 112 -208374
rect 146 -210750 152 -208374
rect 106 -210762 152 -210750
rect -96 -210809 96 -210803
rect -96 -210843 -84 -210809
rect 84 -210843 96 -210809
rect -96 -210849 96 -210843
rect -96 -210917 96 -210911
rect -96 -210951 -84 -210917
rect 84 -210951 96 -210917
rect -96 -210957 96 -210951
rect -152 -211010 -106 -210998
rect -152 -213386 -146 -211010
rect -112 -213386 -106 -211010
rect -152 -213398 -106 -213386
rect 106 -211010 152 -210998
rect 106 -213386 112 -211010
rect 146 -213386 152 -211010
rect 106 -213398 152 -213386
rect -96 -213445 96 -213439
rect -96 -213479 -84 -213445
rect 84 -213479 96 -213445
rect -96 -213485 96 -213479
rect -96 -213553 96 -213547
rect -96 -213587 -84 -213553
rect 84 -213587 96 -213553
rect -96 -213593 96 -213587
rect -152 -213646 -106 -213634
rect -152 -216022 -146 -213646
rect -112 -216022 -106 -213646
rect -152 -216034 -106 -216022
rect 106 -213646 152 -213634
rect 106 -216022 112 -213646
rect 146 -216022 152 -213646
rect 106 -216034 152 -216022
rect -96 -216081 96 -216075
rect -96 -216115 -84 -216081
rect 84 -216115 96 -216081
rect -96 -216121 96 -216115
rect -96 -216189 96 -216183
rect -96 -216223 -84 -216189
rect 84 -216223 96 -216189
rect -96 -216229 96 -216223
rect -152 -216282 -106 -216270
rect -152 -218658 -146 -216282
rect -112 -218658 -106 -216282
rect -152 -218670 -106 -218658
rect 106 -216282 152 -216270
rect 106 -218658 112 -216282
rect 146 -218658 152 -216282
rect 106 -218670 152 -218658
rect -96 -218717 96 -218711
rect -96 -218751 -84 -218717
rect 84 -218751 96 -218717
rect -96 -218757 96 -218751
rect -96 -218825 96 -218819
rect -96 -218859 -84 -218825
rect 84 -218859 96 -218825
rect -96 -218865 96 -218859
rect -152 -218918 -106 -218906
rect -152 -221294 -146 -218918
rect -112 -221294 -106 -218918
rect -152 -221306 -106 -221294
rect 106 -218918 152 -218906
rect 106 -221294 112 -218918
rect 146 -221294 152 -218918
rect 106 -221306 152 -221294
rect -96 -221353 96 -221347
rect -96 -221387 -84 -221353
rect 84 -221387 96 -221353
rect -96 -221393 96 -221387
rect -96 -221461 96 -221455
rect -96 -221495 -84 -221461
rect 84 -221495 96 -221461
rect -96 -221501 96 -221495
rect -152 -221554 -106 -221542
rect -152 -223930 -146 -221554
rect -112 -223930 -106 -221554
rect -152 -223942 -106 -223930
rect 106 -221554 152 -221542
rect 106 -223930 112 -221554
rect 146 -223930 152 -221554
rect 106 -223942 152 -223930
rect -96 -223989 96 -223983
rect -96 -224023 -84 -223989
rect 84 -224023 96 -223989
rect -96 -224029 96 -224023
rect -96 -224097 96 -224091
rect -96 -224131 -84 -224097
rect 84 -224131 96 -224097
rect -96 -224137 96 -224131
rect -152 -224190 -106 -224178
rect -152 -226566 -146 -224190
rect -112 -226566 -106 -224190
rect -152 -226578 -106 -226566
rect 106 -224190 152 -224178
rect 106 -226566 112 -224190
rect 146 -226566 152 -224190
rect 106 -226578 152 -226566
rect -96 -226625 96 -226619
rect -96 -226659 -84 -226625
rect 84 -226659 96 -226625
rect -96 -226665 96 -226659
rect -96 -226733 96 -226727
rect -96 -226767 -84 -226733
rect 84 -226767 96 -226733
rect -96 -226773 96 -226767
rect -152 -226826 -106 -226814
rect -152 -229202 -146 -226826
rect -112 -229202 -106 -226826
rect -152 -229214 -106 -229202
rect 106 -226826 152 -226814
rect 106 -229202 112 -226826
rect 146 -229202 152 -226826
rect 106 -229214 152 -229202
rect -96 -229261 96 -229255
rect -96 -229295 -84 -229261
rect 84 -229295 96 -229261
rect -96 -229301 96 -229295
rect -96 -229369 96 -229363
rect -96 -229403 -84 -229369
rect 84 -229403 96 -229369
rect -96 -229409 96 -229403
rect -152 -229462 -106 -229450
rect -152 -231838 -146 -229462
rect -112 -231838 -106 -229462
rect -152 -231850 -106 -231838
rect 106 -229462 152 -229450
rect 106 -231838 112 -229462
rect 146 -231838 152 -229462
rect 106 -231850 152 -231838
rect -96 -231897 96 -231891
rect -96 -231931 -84 -231897
rect 84 -231931 96 -231897
rect -96 -231937 96 -231931
rect -96 -232005 96 -231999
rect -96 -232039 -84 -232005
rect 84 -232039 96 -232005
rect -96 -232045 96 -232039
rect -152 -232098 -106 -232086
rect -152 -234474 -146 -232098
rect -112 -234474 -106 -232098
rect -152 -234486 -106 -234474
rect 106 -232098 152 -232086
rect 106 -234474 112 -232098
rect 146 -234474 152 -232098
rect 106 -234486 152 -234474
rect -96 -234533 96 -234527
rect -96 -234567 -84 -234533
rect 84 -234567 96 -234533
rect -96 -234573 96 -234567
rect -96 -234641 96 -234635
rect -96 -234675 -84 -234641
rect 84 -234675 96 -234641
rect -96 -234681 96 -234675
rect -152 -234734 -106 -234722
rect -152 -237110 -146 -234734
rect -112 -237110 -106 -234734
rect -152 -237122 -106 -237110
rect 106 -234734 152 -234722
rect 106 -237110 112 -234734
rect 146 -237110 152 -234734
rect 106 -237122 152 -237110
rect -96 -237169 96 -237163
rect -96 -237203 -84 -237169
rect 84 -237203 96 -237169
rect -96 -237209 96 -237203
rect -96 -237277 96 -237271
rect -96 -237311 -84 -237277
rect 84 -237311 96 -237277
rect -96 -237317 96 -237311
rect -152 -237370 -106 -237358
rect -152 -239746 -146 -237370
rect -112 -239746 -106 -237370
rect -152 -239758 -106 -239746
rect 106 -237370 152 -237358
rect 106 -239746 112 -237370
rect 146 -239746 152 -237370
rect 106 -239758 152 -239746
rect -96 -239805 96 -239799
rect -96 -239839 -84 -239805
rect 84 -239839 96 -239805
rect -96 -239845 96 -239839
rect -96 -239913 96 -239907
rect -96 -239947 -84 -239913
rect 84 -239947 96 -239913
rect -96 -239953 96 -239947
rect -152 -240006 -106 -239994
rect -152 -242382 -146 -240006
rect -112 -242382 -106 -240006
rect -152 -242394 -106 -242382
rect 106 -240006 152 -239994
rect 106 -242382 112 -240006
rect 146 -242382 152 -240006
rect 106 -242394 152 -242382
rect -96 -242441 96 -242435
rect -96 -242475 -84 -242441
rect 84 -242475 96 -242441
rect -96 -242481 96 -242475
rect -96 -242549 96 -242543
rect -96 -242583 -84 -242549
rect 84 -242583 96 -242549
rect -96 -242589 96 -242583
rect -152 -242642 -106 -242630
rect -152 -245018 -146 -242642
rect -112 -245018 -106 -242642
rect -152 -245030 -106 -245018
rect 106 -242642 152 -242630
rect 106 -245018 112 -242642
rect 146 -245018 152 -242642
rect 106 -245030 152 -245018
rect -96 -245077 96 -245071
rect -96 -245111 -84 -245077
rect 84 -245111 96 -245077
rect -96 -245117 96 -245111
rect -96 -245185 96 -245179
rect -96 -245219 -84 -245185
rect 84 -245219 96 -245185
rect -96 -245225 96 -245219
rect -152 -245278 -106 -245266
rect -152 -247654 -146 -245278
rect -112 -247654 -106 -245278
rect -152 -247666 -106 -247654
rect 106 -245278 152 -245266
rect 106 -247654 112 -245278
rect 146 -247654 152 -245278
rect 106 -247666 152 -247654
rect -96 -247713 96 -247707
rect -96 -247747 -84 -247713
rect 84 -247747 96 -247713
rect -96 -247753 96 -247747
rect -96 -247821 96 -247815
rect -96 -247855 -84 -247821
rect 84 -247855 96 -247821
rect -96 -247861 96 -247855
rect -152 -247914 -106 -247902
rect -152 -250290 -146 -247914
rect -112 -250290 -106 -247914
rect -152 -250302 -106 -250290
rect 106 -247914 152 -247902
rect 106 -250290 112 -247914
rect 146 -250290 152 -247914
rect 106 -250302 152 -250290
rect -96 -250349 96 -250343
rect -96 -250383 -84 -250349
rect 84 -250383 96 -250349
rect -96 -250389 96 -250383
rect -96 -250457 96 -250451
rect -96 -250491 -84 -250457
rect 84 -250491 96 -250457
rect -96 -250497 96 -250491
rect -152 -250550 -106 -250538
rect -152 -252926 -146 -250550
rect -112 -252926 -106 -250550
rect -152 -252938 -106 -252926
rect 106 -250550 152 -250538
rect 106 -252926 112 -250550
rect 146 -252926 152 -250550
rect 106 -252938 152 -252926
rect -96 -252985 96 -252979
rect -96 -253019 -84 -252985
rect 84 -253019 96 -252985
rect -96 -253025 96 -253019
rect -96 -253093 96 -253087
rect -96 -253127 -84 -253093
rect 84 -253127 96 -253093
rect -96 -253133 96 -253127
rect -152 -253186 -106 -253174
rect -152 -255562 -146 -253186
rect -112 -255562 -106 -253186
rect -152 -255574 -106 -255562
rect 106 -253186 152 -253174
rect 106 -255562 112 -253186
rect 146 -255562 152 -253186
rect 106 -255574 152 -255562
rect -96 -255621 96 -255615
rect -96 -255655 -84 -255621
rect 84 -255655 96 -255621
rect -96 -255661 96 -255655
rect -96 -255729 96 -255723
rect -96 -255763 -84 -255729
rect 84 -255763 96 -255729
rect -96 -255769 96 -255763
rect -152 -255822 -106 -255810
rect -152 -258198 -146 -255822
rect -112 -258198 -106 -255822
rect -152 -258210 -106 -258198
rect 106 -255822 152 -255810
rect 106 -258198 112 -255822
rect 146 -258198 152 -255822
rect 106 -258210 152 -258198
rect -96 -258257 96 -258251
rect -96 -258291 -84 -258257
rect 84 -258291 96 -258257
rect -96 -258297 96 -258291
rect -96 -258365 96 -258359
rect -96 -258399 -84 -258365
rect 84 -258399 96 -258365
rect -96 -258405 96 -258399
rect -152 -258458 -106 -258446
rect -152 -260834 -146 -258458
rect -112 -260834 -106 -258458
rect -152 -260846 -106 -260834
rect 106 -258458 152 -258446
rect 106 -260834 112 -258458
rect 146 -260834 152 -258458
rect 106 -260846 152 -260834
rect -96 -260893 96 -260887
rect -96 -260927 -84 -260893
rect 84 -260927 96 -260893
rect -96 -260933 96 -260927
rect -96 -261001 96 -260995
rect -96 -261035 -84 -261001
rect 84 -261035 96 -261001
rect -96 -261041 96 -261035
rect -152 -261094 -106 -261082
rect -152 -263470 -146 -261094
rect -112 -263470 -106 -261094
rect -152 -263482 -106 -263470
rect 106 -261094 152 -261082
rect 106 -263470 112 -261094
rect 146 -263470 152 -261094
rect 106 -263482 152 -263470
rect -96 -263529 96 -263523
rect -96 -263563 -84 -263529
rect 84 -263563 96 -263529
rect -96 -263569 96 -263563
rect -96 -263637 96 -263631
rect -96 -263671 -84 -263637
rect 84 -263671 96 -263637
rect -96 -263677 96 -263671
rect -152 -263730 -106 -263718
rect -152 -266106 -146 -263730
rect -112 -266106 -106 -263730
rect -152 -266118 -106 -266106
rect 106 -263730 152 -263718
rect 106 -266106 112 -263730
rect 146 -266106 152 -263730
rect 106 -266118 152 -266106
rect -96 -266165 96 -266159
rect -96 -266199 -84 -266165
rect 84 -266199 96 -266165
rect -96 -266205 96 -266199
rect -96 -266273 96 -266267
rect -96 -266307 -84 -266273
rect 84 -266307 96 -266273
rect -96 -266313 96 -266307
rect -152 -266366 -106 -266354
rect -152 -268742 -146 -266366
rect -112 -268742 -106 -266366
rect -152 -268754 -106 -268742
rect 106 -266366 152 -266354
rect 106 -268742 112 -266366
rect 146 -268742 152 -266366
rect 106 -268754 152 -268742
rect -96 -268801 96 -268795
rect -96 -268835 -84 -268801
rect 84 -268835 96 -268801
rect -96 -268841 96 -268835
rect -96 -268909 96 -268903
rect -96 -268943 -84 -268909
rect 84 -268943 96 -268909
rect -96 -268949 96 -268943
rect -152 -269002 -106 -268990
rect -152 -271378 -146 -269002
rect -112 -271378 -106 -269002
rect -152 -271390 -106 -271378
rect 106 -269002 152 -268990
rect 106 -271378 112 -269002
rect 146 -271378 152 -269002
rect 106 -271390 152 -271378
rect -96 -271437 96 -271431
rect -96 -271471 -84 -271437
rect 84 -271471 96 -271437
rect -96 -271477 96 -271471
rect -96 -271545 96 -271539
rect -96 -271579 -84 -271545
rect 84 -271579 96 -271545
rect -96 -271585 96 -271579
rect -152 -271638 -106 -271626
rect -152 -274014 -146 -271638
rect -112 -274014 -106 -271638
rect -152 -274026 -106 -274014
rect 106 -271638 152 -271626
rect 106 -274014 112 -271638
rect 146 -274014 152 -271638
rect 106 -274026 152 -274014
rect -96 -274073 96 -274067
rect -96 -274107 -84 -274073
rect 84 -274107 96 -274073
rect -96 -274113 96 -274107
rect -96 -274181 96 -274175
rect -96 -274215 -84 -274181
rect 84 -274215 96 -274181
rect -96 -274221 96 -274215
rect -152 -274274 -106 -274262
rect -152 -276650 -146 -274274
rect -112 -276650 -106 -274274
rect -152 -276662 -106 -276650
rect 106 -274274 152 -274262
rect 106 -276650 112 -274274
rect 146 -276650 152 -274274
rect 106 -276662 152 -276650
rect -96 -276709 96 -276703
rect -96 -276743 -84 -276709
rect 84 -276743 96 -276709
rect -96 -276749 96 -276743
rect -96 -276817 96 -276811
rect -96 -276851 -84 -276817
rect 84 -276851 96 -276817
rect -96 -276857 96 -276851
rect -152 -276910 -106 -276898
rect -152 -279286 -146 -276910
rect -112 -279286 -106 -276910
rect -152 -279298 -106 -279286
rect 106 -276910 152 -276898
rect 106 -279286 112 -276910
rect 146 -279286 152 -276910
rect 106 -279298 152 -279286
rect -96 -279345 96 -279339
rect -96 -279379 -84 -279345
rect 84 -279379 96 -279345
rect -96 -279385 96 -279379
rect -96 -279453 96 -279447
rect -96 -279487 -84 -279453
rect 84 -279487 96 -279453
rect -96 -279493 96 -279487
rect -152 -279546 -106 -279534
rect -152 -281922 -146 -279546
rect -112 -281922 -106 -279546
rect -152 -281934 -106 -281922
rect 106 -279546 152 -279534
rect 106 -281922 112 -279546
rect 146 -281922 152 -279546
rect 106 -281934 152 -281922
rect -96 -281981 96 -281975
rect -96 -282015 -84 -281981
rect 84 -282015 96 -281981
rect -96 -282021 96 -282015
rect -96 -282089 96 -282083
rect -96 -282123 -84 -282089
rect 84 -282123 96 -282089
rect -96 -282129 96 -282123
rect -152 -282182 -106 -282170
rect -152 -284558 -146 -282182
rect -112 -284558 -106 -282182
rect -152 -284570 -106 -284558
rect 106 -282182 152 -282170
rect 106 -284558 112 -282182
rect 146 -284558 152 -282182
rect 106 -284570 152 -284558
rect -96 -284617 96 -284611
rect -96 -284651 -84 -284617
rect 84 -284651 96 -284617
rect -96 -284657 96 -284651
rect -96 -284725 96 -284719
rect -96 -284759 -84 -284725
rect 84 -284759 96 -284725
rect -96 -284765 96 -284759
rect -152 -284818 -106 -284806
rect -152 -287194 -146 -284818
rect -112 -287194 -106 -284818
rect -152 -287206 -106 -287194
rect 106 -284818 152 -284806
rect 106 -287194 112 -284818
rect 146 -287194 152 -284818
rect 106 -287206 152 -287194
rect -96 -287253 96 -287247
rect -96 -287287 -84 -287253
rect 84 -287287 96 -287253
rect -96 -287293 96 -287287
rect -96 -287361 96 -287355
rect -96 -287395 -84 -287361
rect 84 -287395 96 -287361
rect -96 -287401 96 -287395
rect -152 -287454 -106 -287442
rect -152 -289830 -146 -287454
rect -112 -289830 -106 -287454
rect -152 -289842 -106 -289830
rect 106 -287454 152 -287442
rect 106 -289830 112 -287454
rect 146 -289830 152 -287454
rect 106 -289842 152 -289830
rect -96 -289889 96 -289883
rect -96 -289923 -84 -289889
rect 84 -289923 96 -289889
rect -96 -289929 96 -289923
rect -96 -289997 96 -289991
rect -96 -290031 -84 -289997
rect 84 -290031 96 -289997
rect -96 -290037 96 -290031
rect -152 -290090 -106 -290078
rect -152 -292466 -146 -290090
rect -112 -292466 -106 -290090
rect -152 -292478 -106 -292466
rect 106 -290090 152 -290078
rect 106 -292466 112 -290090
rect 146 -292466 152 -290090
rect 106 -292478 152 -292466
rect -96 -292525 96 -292519
rect -96 -292559 -84 -292525
rect 84 -292559 96 -292525
rect -96 -292565 96 -292559
rect -96 -292633 96 -292627
rect -96 -292667 -84 -292633
rect 84 -292667 96 -292633
rect -96 -292673 96 -292667
rect -152 -292726 -106 -292714
rect -152 -295102 -146 -292726
rect -112 -295102 -106 -292726
rect -152 -295114 -106 -295102
rect 106 -292726 152 -292714
rect 106 -295102 112 -292726
rect 146 -295102 152 -292726
rect 106 -295114 152 -295102
rect -96 -295161 96 -295155
rect -96 -295195 -84 -295161
rect 84 -295195 96 -295161
rect -96 -295201 96 -295195
rect -96 -295269 96 -295263
rect -96 -295303 -84 -295269
rect 84 -295303 96 -295269
rect -96 -295309 96 -295303
rect -152 -295362 -106 -295350
rect -152 -297738 -146 -295362
rect -112 -297738 -106 -295362
rect -152 -297750 -106 -297738
rect 106 -295362 152 -295350
rect 106 -297738 112 -295362
rect 146 -297738 152 -295362
rect 106 -297750 152 -297738
rect -96 -297797 96 -297791
rect -96 -297831 -84 -297797
rect 84 -297831 96 -297797
rect -96 -297837 96 -297831
rect -96 -297905 96 -297899
rect -96 -297939 -84 -297905
rect 84 -297939 96 -297905
rect -96 -297945 96 -297939
rect -152 -297998 -106 -297986
rect -152 -300374 -146 -297998
rect -112 -300374 -106 -297998
rect -152 -300386 -106 -300374
rect 106 -297998 152 -297986
rect 106 -300374 112 -297998
rect 146 -300374 152 -297998
rect 106 -300386 152 -300374
rect -96 -300433 96 -300427
rect -96 -300467 -84 -300433
rect 84 -300467 96 -300433
rect -96 -300473 96 -300467
rect -96 -300541 96 -300535
rect -96 -300575 -84 -300541
rect 84 -300575 96 -300541
rect -96 -300581 96 -300575
rect -152 -300634 -106 -300622
rect -152 -303010 -146 -300634
rect -112 -303010 -106 -300634
rect -152 -303022 -106 -303010
rect 106 -300634 152 -300622
rect 106 -303010 112 -300634
rect 146 -303010 152 -300634
rect 106 -303022 152 -303010
rect -96 -303069 96 -303063
rect -96 -303103 -84 -303069
rect 84 -303103 96 -303069
rect -96 -303109 96 -303103
rect -96 -303177 96 -303171
rect -96 -303211 -84 -303177
rect 84 -303211 96 -303177
rect -96 -303217 96 -303211
rect -152 -303270 -106 -303258
rect -152 -305646 -146 -303270
rect -112 -305646 -106 -303270
rect -152 -305658 -106 -305646
rect 106 -303270 152 -303258
rect 106 -305646 112 -303270
rect 146 -305646 152 -303270
rect 106 -305658 152 -305646
rect -96 -305705 96 -305699
rect -96 -305739 -84 -305705
rect 84 -305739 96 -305705
rect -96 -305745 96 -305739
rect -96 -305813 96 -305807
rect -96 -305847 -84 -305813
rect 84 -305847 96 -305813
rect -96 -305853 96 -305847
rect -152 -305906 -106 -305894
rect -152 -308282 -146 -305906
rect -112 -308282 -106 -305906
rect -152 -308294 -106 -308282
rect 106 -305906 152 -305894
rect 106 -308282 112 -305906
rect 146 -308282 152 -305906
rect 106 -308294 152 -308282
rect -96 -308341 96 -308335
rect -96 -308375 -84 -308341
rect 84 -308375 96 -308341
rect -96 -308381 96 -308375
rect -96 -308449 96 -308443
rect -96 -308483 -84 -308449
rect 84 -308483 96 -308449
rect -96 -308489 96 -308483
rect -152 -308542 -106 -308530
rect -152 -310918 -146 -308542
rect -112 -310918 -106 -308542
rect -152 -310930 -106 -310918
rect 106 -308542 152 -308530
rect 106 -310918 112 -308542
rect 146 -310918 152 -308542
rect 106 -310930 152 -310918
rect -96 -310977 96 -310971
rect -96 -311011 -84 -310977
rect 84 -311011 96 -310977
rect -96 -311017 96 -311011
rect -96 -311085 96 -311079
rect -96 -311119 -84 -311085
rect 84 -311119 96 -311085
rect -96 -311125 96 -311119
rect -152 -311178 -106 -311166
rect -152 -313554 -146 -311178
rect -112 -313554 -106 -311178
rect -152 -313566 -106 -313554
rect 106 -311178 152 -311166
rect 106 -313554 112 -311178
rect 146 -313554 152 -311178
rect 106 -313566 152 -313554
rect -96 -313613 96 -313607
rect -96 -313647 -84 -313613
rect 84 -313647 96 -313613
rect -96 -313653 96 -313647
rect -96 -313721 96 -313715
rect -96 -313755 -84 -313721
rect 84 -313755 96 -313721
rect -96 -313761 96 -313755
rect -152 -313814 -106 -313802
rect -152 -316190 -146 -313814
rect -112 -316190 -106 -313814
rect -152 -316202 -106 -316190
rect 106 -313814 152 -313802
rect 106 -316190 112 -313814
rect 146 -316190 152 -313814
rect 106 -316202 152 -316190
rect -96 -316249 96 -316243
rect -96 -316283 -84 -316249
rect 84 -316283 96 -316249
rect -96 -316289 96 -316283
rect -96 -316357 96 -316351
rect -96 -316391 -84 -316357
rect 84 -316391 96 -316357
rect -96 -316397 96 -316391
rect -152 -316450 -106 -316438
rect -152 -318826 -146 -316450
rect -112 -318826 -106 -316450
rect -152 -318838 -106 -318826
rect 106 -316450 152 -316438
rect 106 -318826 112 -316450
rect 146 -318826 152 -316450
rect 106 -318838 152 -318826
rect -96 -318885 96 -318879
rect -96 -318919 -84 -318885
rect 84 -318919 96 -318885
rect -96 -318925 96 -318919
rect -96 -318993 96 -318987
rect -96 -319027 -84 -318993
rect 84 -319027 96 -318993
rect -96 -319033 96 -319027
rect -152 -319086 -106 -319074
rect -152 -321462 -146 -319086
rect -112 -321462 -106 -319086
rect -152 -321474 -106 -321462
rect 106 -319086 152 -319074
rect 106 -321462 112 -319086
rect 146 -321462 152 -319086
rect 106 -321474 152 -321462
rect -96 -321521 96 -321515
rect -96 -321555 -84 -321521
rect 84 -321555 96 -321521
rect -96 -321561 96 -321555
rect -96 -321629 96 -321623
rect -96 -321663 -84 -321629
rect 84 -321663 96 -321629
rect -96 -321669 96 -321663
rect -152 -321722 -106 -321710
rect -152 -324098 -146 -321722
rect -112 -324098 -106 -321722
rect -152 -324110 -106 -324098
rect 106 -321722 152 -321710
rect 106 -324098 112 -321722
rect 146 -324098 152 -321722
rect 106 -324110 152 -324098
rect -96 -324157 96 -324151
rect -96 -324191 -84 -324157
rect 84 -324191 96 -324157
rect -96 -324197 96 -324191
rect -96 -324265 96 -324259
rect -96 -324299 -84 -324265
rect 84 -324299 96 -324265
rect -96 -324305 96 -324299
rect -152 -324358 -106 -324346
rect -152 -326734 -146 -324358
rect -112 -326734 -106 -324358
rect -152 -326746 -106 -326734
rect 106 -324358 152 -324346
rect 106 -326734 112 -324358
rect 146 -326734 152 -324358
rect 106 -326746 152 -326734
rect -96 -326793 96 -326787
rect -96 -326827 -84 -326793
rect 84 -326827 96 -326793
rect -96 -326833 96 -326827
rect -96 -326901 96 -326895
rect -96 -326935 -84 -326901
rect 84 -326935 96 -326901
rect -96 -326941 96 -326935
rect -152 -326994 -106 -326982
rect -152 -329370 -146 -326994
rect -112 -329370 -106 -326994
rect -152 -329382 -106 -329370
rect 106 -326994 152 -326982
rect 106 -329370 112 -326994
rect 146 -329370 152 -326994
rect 106 -329382 152 -329370
rect -96 -329429 96 -329423
rect -96 -329463 -84 -329429
rect 84 -329463 96 -329429
rect -96 -329469 96 -329463
rect -96 -329537 96 -329531
rect -96 -329571 -84 -329537
rect 84 -329571 96 -329537
rect -96 -329577 96 -329571
rect -152 -329630 -106 -329618
rect -152 -332006 -146 -329630
rect -112 -332006 -106 -329630
rect -152 -332018 -106 -332006
rect 106 -329630 152 -329618
rect 106 -332006 112 -329630
rect 146 -332006 152 -329630
rect 106 -332018 152 -332006
rect -96 -332065 96 -332059
rect -96 -332099 -84 -332065
rect 84 -332099 96 -332065
rect -96 -332105 96 -332099
rect -96 -332173 96 -332167
rect -96 -332207 -84 -332173
rect 84 -332207 96 -332173
rect -96 -332213 96 -332207
rect -152 -332266 -106 -332254
rect -152 -334642 -146 -332266
rect -112 -334642 -106 -332266
rect -152 -334654 -106 -334642
rect 106 -332266 152 -332254
rect 106 -334642 112 -332266
rect 146 -334642 152 -332266
rect 106 -334654 152 -334642
rect -96 -334701 96 -334695
rect -96 -334735 -84 -334701
rect 84 -334735 96 -334701
rect -96 -334741 96 -334735
rect -96 -334809 96 -334803
rect -96 -334843 -84 -334809
rect 84 -334843 96 -334809
rect -96 -334849 96 -334843
rect -152 -334902 -106 -334890
rect -152 -337278 -146 -334902
rect -112 -337278 -106 -334902
rect -152 -337290 -106 -337278
rect 106 -334902 152 -334890
rect 106 -337278 112 -334902
rect 146 -337278 152 -334902
rect 106 -337290 152 -337278
rect -96 -337337 96 -337331
rect -96 -337371 -84 -337337
rect 84 -337371 96 -337337
rect -96 -337377 96 -337371
<< properties >>
string FIXED_BBOX -263 -337492 263 337492
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 12.0 l 1.0 m 256 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
