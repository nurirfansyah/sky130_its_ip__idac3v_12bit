magic
tech sky130A
magscale 1 2
timestamp 1717438951
<< metal1 >>
rect 4864 2590 5064 2790
rect 4864 2362 5064 2562
rect 4864 -630 5064 -430
rect 4864 -858 5064 -658
rect 4864 -1086 5064 -886
rect 5218 -1314 5418 -1114
rect 33354 -1314 34457 -1114
rect 4864 -2462 5064 -2262
rect 4864 -2690 5064 -2490
rect 4864 -2918 5064 -2718
rect 4864 -3146 5064 -2946
use icell8scs  x1
timestamp 1717438951
transform 1 0 0 0 1 0
box 4862 -5160 33945 2790
use icell8scs  x2
timestamp 1717438951
transform 1 0 29039 0 1 0
box 4862 -5160 33945 2790
<< labels >>
flabel metal1 4864 2362 5064 2562 0 FreeSans 256 0 0 0 iout
port 0 nsew
flabel metal1 4864 -630 5064 -430 0 FreeSans 256 0 0 0 avdd
port 1 nsew
flabel metal1 4864 -858 5064 -658 0 FreeSans 256 0 0 0 pbias
port 2 nsew
flabel metal1 4864 2590 5064 2790 0 FreeSans 256 0 0 0 ioutn
port 3 nsew
flabel metal1 5218 -1314 5418 -1114 0 FreeSans 256 0 0 0 sw
port 4 nsew
flabel metal1 4864 -1086 5064 -886 0 FreeSans 256 0 0 0 pcbias
port 5 nsew
flabel metal1 4864 -2462 5064 -2262 0 FreeSans 256 0 0 0 idir_sel
port 6 nsew
flabel metal1 4864 -2690 5064 -2490 0 FreeSans 256 0 0 0 ncbias
port 7 nsew
flabel metal1 4864 -2918 5064 -2718 0 FreeSans 256 0 0 0 nbias
port 8 nsew
flabel metal1 4864 -3146 5064 -2946 0 FreeSans 256 0 0 0 avss
port 9 nsew
<< end >>
