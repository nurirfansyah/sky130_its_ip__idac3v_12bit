magic
tech sky130A
magscale 1 2
timestamp 1717439242
<< nwell >>
rect -1458 -1097 1458 1097
<< mvpmos >>
rect -1200 -800 1200 800
<< mvpdiff >>
rect -1258 788 -1200 800
rect -1258 -788 -1246 788
rect -1212 -788 -1200 788
rect -1258 -800 -1200 -788
rect 1200 788 1258 800
rect 1200 -788 1212 788
rect 1246 -788 1258 788
rect 1200 -800 1258 -788
<< mvpdiffc >>
rect -1246 -788 -1212 788
rect 1212 -788 1246 788
<< mvnsubdiff >>
rect -1392 1019 1392 1031
rect -1392 985 -1284 1019
rect 1284 985 1392 1019
rect -1392 973 1392 985
rect -1392 923 -1334 973
rect -1392 -923 -1380 923
rect -1346 -923 -1334 923
rect 1334 923 1392 973
rect -1392 -973 -1334 -923
rect 1334 -923 1346 923
rect 1380 -923 1392 923
rect 1334 -973 1392 -923
rect -1392 -985 1392 -973
rect -1392 -1019 -1284 -985
rect 1284 -1019 1392 -985
rect -1392 -1031 1392 -1019
<< mvnsubdiffcont >>
rect -1284 985 1284 1019
rect -1380 -923 -1346 923
rect 1346 -923 1380 923
rect -1284 -1019 1284 -985
<< poly >>
rect -1200 881 1200 897
rect -1200 847 -1184 881
rect 1184 847 1200 881
rect -1200 800 1200 847
rect -1200 -847 1200 -800
rect -1200 -881 -1184 -847
rect 1184 -881 1200 -847
rect -1200 -897 1200 -881
<< polycont >>
rect -1184 847 1184 881
rect -1184 -881 1184 -847
<< locali >>
rect -1380 985 -1284 1019
rect 1284 985 1380 1019
rect -1380 923 -1346 985
rect 1346 923 1380 985
rect -1200 847 -1184 881
rect 1184 847 1200 881
rect -1246 788 -1212 804
rect -1246 -804 -1212 -788
rect 1212 788 1246 804
rect 1212 -804 1246 -788
rect -1200 -881 -1184 -847
rect 1184 -881 1200 -847
rect -1380 -985 -1346 -923
rect 1346 -985 1380 -923
rect -1380 -1019 -1284 -985
rect 1284 -1019 1380 -985
<< viali >>
rect -1184 847 1184 881
rect -1246 -788 -1212 788
rect 1212 -788 1246 788
rect -1184 -881 1184 -847
<< metal1 >>
rect -1196 881 1196 887
rect -1196 847 -1184 881
rect 1184 847 1196 881
rect -1196 841 1196 847
rect -1252 788 -1206 800
rect -1252 -788 -1246 788
rect -1212 -788 -1206 788
rect -1252 -800 -1206 -788
rect 1206 788 1252 800
rect 1206 -788 1212 788
rect 1246 -788 1252 788
rect 1206 -800 1252 -788
rect -1196 -847 1196 -841
rect -1196 -881 -1184 -847
rect 1184 -881 1196 -847
rect -1196 -887 1196 -881
<< properties >>
string FIXED_BBOX -1363 -1002 1363 1002
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 8.0 l 12.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
