magic
tech sky130A
magscale 1 2
timestamp 1717438951
<< metal1 >>
rect 19010 -1314 19937 -1114
use icell4scs  x1
timestamp 1717438951
transform 1 0 0 0 1 0
box 4862 -5160 19426 2790
use icell4scs  x2
timestamp 1717438951
transform 1 0 14519 0 1 0
box 4862 -5160 19426 2790
<< end >>
